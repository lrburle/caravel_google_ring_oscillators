VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO scs130hd_mpr2aa_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130hd_mpr2aa_8 0 0 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT 8.41 0.35 8.74 1.08 ;
      RECT 8.37 0.235 8.55 0.885 ;
      RECT 4.87 2.035 5.2 2.365 ;
      RECT 3.665 2.05 5.2 2.35 ;
      RECT 3.665 0.93 3.965 2.35 ;
      RECT 3.41 0.915 3.74 1.245 ;
      RECT 8.89 1.475 9.22 2.205 ;
      RECT 6.81 1.075 7.14 1.805 ;
      RECT 5.25 0.515 5.58 1.245 ;
      RECT 4.37 0.515 4.7 1.245 ;
      RECT 2.69 0.915 3.02 1.645 ;
      RECT 1.69 0.355 2.02 1.085 ;
      RECT 0.25 1.075 0.58 1.805 ;
    LAYER via2 ;
      RECT 8.955 1.54 9.155 1.74 ;
      RECT 8.475 0.815 8.675 1.015 ;
      RECT 6.875 1.54 7.075 1.74 ;
      RECT 5.315 0.98 5.515 1.18 ;
      RECT 4.935 2.1 5.135 2.3 ;
      RECT 4.435 0.98 4.635 1.18 ;
      RECT 3.475 0.98 3.675 1.18 ;
      RECT 2.755 0.98 2.955 1.18 ;
      RECT 1.755 0.42 1.955 0.62 ;
      RECT 0.315 1.54 0.515 1.74 ;
    LAYER met2 ;
      RECT 5.985 0.955 6.22 1.215 ;
      RECT 9.13 0.735 9.295 0.995 ;
      RECT 9.035 0.725 9.05 0.995 ;
      RECT 7.635 0.295 7.675 0.435 ;
      RECT 9.05 0.73 9.13 0.995 ;
      RECT 8.995 0.725 9.035 0.961 ;
      RECT 8.981 0.725 8.995 0.961 ;
      RECT 8.895 0.73 8.981 0.963 ;
      RECT 8.85 0.737 8.895 0.965 ;
      RECT 8.82 0.737 8.85 0.967 ;
      RECT 8.795 0.732 8.82 0.969 ;
      RECT 8.765 0.728 8.795 0.978 ;
      RECT 8.755 0.725 8.765 0.99 ;
      RECT 8.75 0.725 8.755 0.998 ;
      RECT 8.745 0.725 8.75 1.003 ;
      RECT 8.735 0.724 8.745 1.013 ;
      RECT 8.73 0.723 8.735 1.023 ;
      RECT 8.715 0.722 8.73 1.028 ;
      RECT 8.687 0.719 8.715 1.055 ;
      RECT 8.601 0.711 8.687 1.055 ;
      RECT 8.515 0.7 8.601 1.055 ;
      RECT 8.475 0.685 8.515 1.055 ;
      RECT 8.435 0.659 8.475 1.055 ;
      RECT 8.43 0.641 8.435 0.867 ;
      RECT 8.42 0.637 8.43 0.857 ;
      RECT 8.405 0.627 8.42 0.844 ;
      RECT 8.385 0.611 8.405 0.829 ;
      RECT 8.37 0.596 8.385 0.814 ;
      RECT 8.36 0.585 8.37 0.804 ;
      RECT 8.335 0.569 8.36 0.793 ;
      RECT 8.33 0.556 8.335 0.783 ;
      RECT 8.325 0.552 8.33 0.778 ;
      RECT 8.27 0.538 8.325 0.756 ;
      RECT 8.231 0.519 8.27 0.72 ;
      RECT 8.145 0.493 8.231 0.673 ;
      RECT 8.141 0.475 8.145 0.639 ;
      RECT 8.055 0.456 8.141 0.617 ;
      RECT 8.05 0.438 8.055 0.595 ;
      RECT 8.045 0.436 8.05 0.593 ;
      RECT 8.035 0.435 8.045 0.588 ;
      RECT 7.975 0.422 8.035 0.574 ;
      RECT 7.93 0.4 7.975 0.553 ;
      RECT 7.87 0.377 7.93 0.532 ;
      RECT 7.806 0.352 7.87 0.507 ;
      RECT 7.72 0.322 7.806 0.476 ;
      RECT 7.705 0.302 7.72 0.455 ;
      RECT 7.675 0.297 7.705 0.446 ;
      RECT 7.622 0.295 7.635 0.435 ;
      RECT 7.536 0.295 7.622 0.437 ;
      RECT 7.45 0.295 7.536 0.439 ;
      RECT 7.43 0.295 7.45 0.443 ;
      RECT 7.385 0.297 7.43 0.454 ;
      RECT 7.345 0.307 7.385 0.47 ;
      RECT 7.341 0.316 7.345 0.478 ;
      RECT 7.255 0.336 7.341 0.494 ;
      RECT 7.245 0.355 7.255 0.512 ;
      RECT 7.24 0.357 7.245 0.515 ;
      RECT 7.23 0.361 7.24 0.518 ;
      RECT 7.21 0.366 7.23 0.528 ;
      RECT 7.18 0.376 7.21 0.548 ;
      RECT 7.175 0.383 7.18 0.562 ;
      RECT 7.165 0.387 7.175 0.569 ;
      RECT 7.15 0.395 7.165 0.58 ;
      RECT 7.14 0.405 7.15 0.591 ;
      RECT 7.13 0.412 7.14 0.599 ;
      RECT 7.105 0.425 7.13 0.614 ;
      RECT 7.041 0.461 7.105 0.653 ;
      RECT 6.955 0.524 7.041 0.717 ;
      RECT 6.92 0.575 6.955 0.77 ;
      RECT 6.915 0.592 6.92 0.787 ;
      RECT 6.9 0.601 6.915 0.794 ;
      RECT 6.88 0.616 6.9 0.808 ;
      RECT 6.875 0.627 6.88 0.818 ;
      RECT 6.855 0.64 6.875 0.828 ;
      RECT 6.85 0.65 6.855 0.838 ;
      RECT 6.835 0.655 6.85 0.847 ;
      RECT 6.825 0.665 6.835 0.858 ;
      RECT 6.795 0.682 6.825 0.875 ;
      RECT 6.785 0.7 6.795 0.893 ;
      RECT 6.77 0.711 6.785 0.904 ;
      RECT 6.73 0.735 6.77 0.92 ;
      RECT 6.695 0.769 6.73 0.937 ;
      RECT 6.665 0.792 6.695 0.949 ;
      RECT 6.65 0.802 6.665 0.958 ;
      RECT 6.61 0.812 6.65 0.969 ;
      RECT 6.59 0.823 6.61 0.981 ;
      RECT 6.585 0.827 6.59 0.988 ;
      RECT 6.57 0.831 6.585 0.993 ;
      RECT 6.56 0.836 6.57 0.998 ;
      RECT 6.555 0.839 6.56 1.001 ;
      RECT 6.525 0.845 6.555 1.008 ;
      RECT 6.49 0.855 6.525 1.022 ;
      RECT 6.43 0.87 6.49 1.042 ;
      RECT 6.375 0.89 6.43 1.066 ;
      RECT 6.346 0.905 6.375 1.084 ;
      RECT 6.26 0.925 6.346 1.109 ;
      RECT 6.255 0.94 6.26 1.129 ;
      RECT 6.245 0.943 6.255 1.13 ;
      RECT 6.22 0.95 6.245 1.215 ;
      RECT 8.915 1.443 9.195 1.78 ;
      RECT 8.915 1.453 9.2 1.738 ;
      RECT 8.915 1.462 9.205 1.635 ;
      RECT 8.915 1.477 9.21 1.503 ;
      RECT 8.915 1.305 9.175 1.78 ;
      RECT 6.635 2.185 6.645 2.375 ;
      RECT 4.895 2.06 5.175 2.34 ;
      RECT 7.94 1 7.945 1.485 ;
      RECT 7.835 1 7.895 1.26 ;
      RECT 8.16 1.97 8.165 2.045 ;
      RECT 8.15 1.837 8.16 2.08 ;
      RECT 8.14 1.672 8.15 2.101 ;
      RECT 8.135 1.542 8.14 2.117 ;
      RECT 8.125 1.432 8.135 2.133 ;
      RECT 8.12 1.331 8.125 2.15 ;
      RECT 8.115 1.313 8.12 2.16 ;
      RECT 8.11 1.295 8.115 2.17 ;
      RECT 8.1 1.27 8.11 2.185 ;
      RECT 8.095 1.25 8.1 2.2 ;
      RECT 8.075 1 8.095 2.225 ;
      RECT 8.06 1 8.075 2.258 ;
      RECT 8.03 1 8.06 2.28 ;
      RECT 8.01 1 8.03 2.294 ;
      RECT 7.99 1 8.01 1.81 ;
      RECT 8.005 1.877 8.01 2.299 ;
      RECT 8 1.907 8.005 2.301 ;
      RECT 7.995 1.92 8 2.304 ;
      RECT 7.99 1.93 7.995 2.308 ;
      RECT 7.985 1 7.99 1.728 ;
      RECT 7.985 1.94 7.99 2.31 ;
      RECT 7.98 1 7.985 1.705 ;
      RECT 7.97 1.962 7.985 2.31 ;
      RECT 7.965 1 7.98 1.65 ;
      RECT 7.96 1.987 7.97 2.31 ;
      RECT 7.96 1 7.965 1.595 ;
      RECT 7.95 1 7.96 1.543 ;
      RECT 7.955 2 7.96 2.311 ;
      RECT 7.95 2.012 7.955 2.312 ;
      RECT 7.945 1 7.95 1.503 ;
      RECT 7.945 2.025 7.95 2.313 ;
      RECT 7.93 2.04 7.945 2.314 ;
      RECT 7.935 1 7.94 1.465 ;
      RECT 7.93 1 7.935 1.43 ;
      RECT 7.925 1 7.93 1.405 ;
      RECT 7.92 2.067 7.93 2.316 ;
      RECT 7.915 1 7.925 1.363 ;
      RECT 7.915 2.085 7.92 2.317 ;
      RECT 7.91 1 7.915 1.323 ;
      RECT 7.91 2.092 7.915 2.318 ;
      RECT 7.905 1 7.91 1.295 ;
      RECT 7.9 2.11 7.91 2.319 ;
      RECT 7.895 1 7.905 1.275 ;
      RECT 7.89 2.13 7.9 2.321 ;
      RECT 7.88 2.147 7.89 2.322 ;
      RECT 7.845 2.17 7.88 2.325 ;
      RECT 7.79 2.188 7.845 2.331 ;
      RECT 7.704 2.196 7.79 2.34 ;
      RECT 7.618 2.207 7.704 2.351 ;
      RECT 7.532 2.217 7.618 2.362 ;
      RECT 7.446 2.227 7.532 2.374 ;
      RECT 7.36 2.237 7.446 2.385 ;
      RECT 7.34 2.243 7.36 2.391 ;
      RECT 7.26 2.245 7.34 2.395 ;
      RECT 7.255 2.244 7.26 2.4 ;
      RECT 7.247 2.243 7.255 2.4 ;
      RECT 7.161 2.239 7.247 2.398 ;
      RECT 7.075 2.231 7.161 2.395 ;
      RECT 6.989 2.222 7.075 2.391 ;
      RECT 6.903 2.214 6.989 2.388 ;
      RECT 6.817 2.206 6.903 2.384 ;
      RECT 6.731 2.197 6.817 2.381 ;
      RECT 6.645 2.189 6.731 2.377 ;
      RECT 6.59 2.182 6.635 2.375 ;
      RECT 6.505 2.175 6.59 2.373 ;
      RECT 6.431 2.167 6.505 2.369 ;
      RECT 6.345 2.159 6.431 2.366 ;
      RECT 6.342 2.155 6.345 2.364 ;
      RECT 6.256 2.151 6.342 2.363 ;
      RECT 6.17 2.143 6.256 2.36 ;
      RECT 6.085 2.138 6.17 2.357 ;
      RECT 5.999 2.135 6.085 2.354 ;
      RECT 5.913 2.133 5.999 2.351 ;
      RECT 5.827 2.13 5.913 2.348 ;
      RECT 5.741 2.127 5.827 2.345 ;
      RECT 5.655 2.124 5.741 2.342 ;
      RECT 5.579 2.122 5.655 2.339 ;
      RECT 5.493 2.119 5.579 2.336 ;
      RECT 5.407 2.116 5.493 2.334 ;
      RECT 5.321 2.114 5.407 2.331 ;
      RECT 5.235 2.111 5.321 2.328 ;
      RECT 5.175 2.102 5.235 2.326 ;
      RECT 7.685 1.72 7.76 1.98 ;
      RECT 7.665 1.7 7.67 1.98 ;
      RECT 6.985 1.485 7.09 1.78 ;
      RECT 1.43 1.46 1.5 1.72 ;
      RECT 7.325 1.335 7.33 1.706 ;
      RECT 7.315 1.39 7.32 1.706 ;
      RECT 7.62 0.56 7.68 0.82 ;
      RECT 7.675 1.715 7.685 1.98 ;
      RECT 7.67 1.705 7.675 1.98 ;
      RECT 7.59 1.652 7.665 1.98 ;
      RECT 7.615 0.56 7.62 0.84 ;
      RECT 7.605 0.56 7.615 0.86 ;
      RECT 7.59 0.56 7.605 0.89 ;
      RECT 7.575 0.56 7.59 0.933 ;
      RECT 7.57 1.595 7.59 1.98 ;
      RECT 7.56 0.56 7.575 0.97 ;
      RECT 7.555 1.575 7.57 1.98 ;
      RECT 7.555 0.56 7.56 0.993 ;
      RECT 7.545 0.56 7.555 1.018 ;
      RECT 7.515 1.542 7.555 1.98 ;
      RECT 7.52 0.56 7.545 1.068 ;
      RECT 7.515 0.56 7.52 1.123 ;
      RECT 7.51 0.56 7.515 1.165 ;
      RECT 7.5 1.505 7.515 1.98 ;
      RECT 7.505 0.56 7.51 1.208 ;
      RECT 7.5 0.56 7.505 1.273 ;
      RECT 7.495 0.56 7.5 1.295 ;
      RECT 7.495 1.493 7.5 1.845 ;
      RECT 7.49 0.56 7.495 1.363 ;
      RECT 7.49 1.485 7.495 1.828 ;
      RECT 7.485 0.56 7.49 1.408 ;
      RECT 7.48 1.467 7.49 1.805 ;
      RECT 7.48 0.56 7.485 1.445 ;
      RECT 7.47 0.56 7.48 1.785 ;
      RECT 7.465 0.56 7.47 1.768 ;
      RECT 7.46 0.56 7.465 1.753 ;
      RECT 7.455 0.56 7.46 1.738 ;
      RECT 7.435 0.56 7.455 1.728 ;
      RECT 7.43 0.56 7.435 1.718 ;
      RECT 7.42 0.56 7.43 1.714 ;
      RECT 7.415 0.837 7.42 1.713 ;
      RECT 7.41 0.86 7.415 1.712 ;
      RECT 7.405 0.89 7.41 1.711 ;
      RECT 7.4 0.917 7.405 1.71 ;
      RECT 7.395 0.945 7.4 1.71 ;
      RECT 7.39 0.972 7.395 1.71 ;
      RECT 7.385 0.992 7.39 1.71 ;
      RECT 7.38 1.02 7.385 1.71 ;
      RECT 7.37 1.062 7.38 1.71 ;
      RECT 7.36 1.107 7.37 1.709 ;
      RECT 7.355 1.16 7.36 1.708 ;
      RECT 7.35 1.192 7.355 1.707 ;
      RECT 7.345 1.212 7.35 1.706 ;
      RECT 7.34 1.25 7.345 1.706 ;
      RECT 7.335 1.272 7.34 1.706 ;
      RECT 7.33 1.297 7.335 1.706 ;
      RECT 7.32 1.362 7.325 1.706 ;
      RECT 7.305 1.422 7.315 1.706 ;
      RECT 7.29 1.432 7.305 1.706 ;
      RECT 7.27 1.442 7.29 1.706 ;
      RECT 7.24 1.447 7.27 1.703 ;
      RECT 7.18 1.457 7.24 1.7 ;
      RECT 7.16 1.466 7.18 1.705 ;
      RECT 7.135 1.472 7.16 1.718 ;
      RECT 7.115 1.477 7.135 1.733 ;
      RECT 7.09 1.482 7.115 1.78 ;
      RECT 6.961 1.484 6.985 1.78 ;
      RECT 6.875 1.479 6.961 1.78 ;
      RECT 6.835 1.476 6.875 1.78 ;
      RECT 6.785 1.478 6.835 1.76 ;
      RECT 6.755 1.482 6.785 1.76 ;
      RECT 6.676 1.492 6.755 1.76 ;
      RECT 6.59 1.507 6.676 1.761 ;
      RECT 6.54 1.517 6.59 1.762 ;
      RECT 6.532 1.52 6.54 1.762 ;
      RECT 6.446 1.522 6.532 1.763 ;
      RECT 6.36 1.526 6.446 1.763 ;
      RECT 6.274 1.53 6.36 1.764 ;
      RECT 6.188 1.533 6.274 1.765 ;
      RECT 6.102 1.537 6.188 1.765 ;
      RECT 6.016 1.541 6.102 1.766 ;
      RECT 5.93 1.544 6.016 1.767 ;
      RECT 5.844 1.548 5.93 1.767 ;
      RECT 5.758 1.552 5.844 1.768 ;
      RECT 5.672 1.556 5.758 1.769 ;
      RECT 5.586 1.559 5.672 1.769 ;
      RECT 5.5 1.563 5.586 1.77 ;
      RECT 5.47 1.565 5.5 1.77 ;
      RECT 5.384 1.568 5.47 1.771 ;
      RECT 5.298 1.572 5.384 1.772 ;
      RECT 5.212 1.576 5.298 1.773 ;
      RECT 5.126 1.579 5.212 1.773 ;
      RECT 5.04 1.583 5.126 1.774 ;
      RECT 5.005 1.588 5.04 1.775 ;
      RECT 4.95 1.598 5.005 1.782 ;
      RECT 4.925 1.61 4.95 1.792 ;
      RECT 4.89 1.623 4.925 1.8 ;
      RECT 4.85 1.64 4.89 1.823 ;
      RECT 4.83 1.653 4.85 1.85 ;
      RECT 4.8 1.665 4.83 1.878 ;
      RECT 4.795 1.673 4.8 1.898 ;
      RECT 4.79 1.676 4.795 1.908 ;
      RECT 4.74 1.688 4.79 1.942 ;
      RECT 4.73 1.703 4.74 1.975 ;
      RECT 4.72 1.709 4.73 1.988 ;
      RECT 4.71 1.716 4.72 2 ;
      RECT 4.685 1.729 4.71 2.018 ;
      RECT 4.67 1.744 4.685 2.04 ;
      RECT 4.66 1.752 4.67 2.056 ;
      RECT 4.645 1.761 4.66 2.071 ;
      RECT 4.635 1.771 4.645 2.085 ;
      RECT 4.616 1.784 4.635 2.102 ;
      RECT 4.53 1.829 4.616 2.167 ;
      RECT 4.515 1.874 4.53 2.225 ;
      RECT 4.51 1.883 4.515 2.238 ;
      RECT 4.5 1.89 4.51 2.243 ;
      RECT 4.495 1.895 4.5 2.247 ;
      RECT 4.475 1.905 4.495 2.254 ;
      RECT 4.45 1.925 4.475 2.268 ;
      RECT 4.415 1.95 4.45 2.288 ;
      RECT 4.4 1.973 4.415 2.303 ;
      RECT 4.39 1.983 4.4 2.308 ;
      RECT 4.38 1.991 4.39 2.315 ;
      RECT 4.37 2 4.38 2.321 ;
      RECT 4.35 2.012 4.37 2.323 ;
      RECT 4.34 2.025 4.35 2.325 ;
      RECT 4.315 2.04 4.34 2.328 ;
      RECT 4.295 2.057 4.315 2.332 ;
      RECT 4.255 2.085 4.295 2.338 ;
      RECT 4.19 2.132 4.255 2.347 ;
      RECT 4.175 2.165 4.19 2.355 ;
      RECT 4.17 2.172 4.175 2.357 ;
      RECT 4.12 2.197 4.17 2.362 ;
      RECT 4.105 2.221 4.12 2.369 ;
      RECT 4.055 2.226 4.105 2.37 ;
      RECT 3.969 2.23 4.055 2.37 ;
      RECT 3.883 2.23 3.969 2.37 ;
      RECT 3.797 2.23 3.883 2.371 ;
      RECT 3.711 2.23 3.797 2.371 ;
      RECT 3.625 2.23 3.711 2.371 ;
      RECT 3.559 2.23 3.625 2.371 ;
      RECT 3.473 2.23 3.559 2.372 ;
      RECT 3.387 2.23 3.473 2.372 ;
      RECT 3.301 2.231 3.387 2.373 ;
      RECT 3.215 2.231 3.301 2.373 ;
      RECT 3.129 2.231 3.215 2.373 ;
      RECT 3.043 2.231 3.129 2.374 ;
      RECT 2.957 2.231 3.043 2.374 ;
      RECT 2.871 2.232 2.957 2.375 ;
      RECT 2.785 2.232 2.871 2.375 ;
      RECT 2.765 2.232 2.785 2.375 ;
      RECT 2.679 2.232 2.765 2.375 ;
      RECT 2.593 2.232 2.679 2.375 ;
      RECT 2.507 2.233 2.593 2.375 ;
      RECT 2.421 2.233 2.507 2.375 ;
      RECT 2.335 2.233 2.421 2.375 ;
      RECT 2.249 2.234 2.335 2.375 ;
      RECT 2.163 2.234 2.249 2.375 ;
      RECT 2.077 2.234 2.163 2.375 ;
      RECT 1.991 2.234 2.077 2.375 ;
      RECT 1.905 2.235 1.991 2.375 ;
      RECT 1.855 2.232 1.905 2.375 ;
      RECT 1.845 2.23 1.855 2.374 ;
      RECT 1.841 2.23 1.845 2.373 ;
      RECT 1.755 2.225 1.841 2.368 ;
      RECT 1.733 2.218 1.755 2.362 ;
      RECT 1.647 2.209 1.733 2.356 ;
      RECT 1.561 2.196 1.647 2.347 ;
      RECT 1.475 2.182 1.561 2.337 ;
      RECT 1.43 2.172 1.475 2.33 ;
      RECT 1.41 1.46 1.43 1.738 ;
      RECT 1.41 2.165 1.43 2.326 ;
      RECT 1.38 1.46 1.41 1.76 ;
      RECT 1.37 2.132 1.41 2.323 ;
      RECT 1.365 1.46 1.38 1.78 ;
      RECT 1.365 2.097 1.37 2.321 ;
      RECT 1.36 1.46 1.365 1.905 ;
      RECT 1.36 2.057 1.365 2.321 ;
      RECT 1.35 1.46 1.36 2.321 ;
      RECT 1.275 1.46 1.35 2.315 ;
      RECT 1.245 1.46 1.275 2.305 ;
      RECT 1.24 1.46 1.245 2.297 ;
      RECT 1.235 1.502 1.24 2.29 ;
      RECT 1.225 1.571 1.235 2.281 ;
      RECT 1.22 1.641 1.225 2.233 ;
      RECT 1.215 1.705 1.22 2.13 ;
      RECT 1.21 1.74 1.215 2.085 ;
      RECT 1.208 1.777 1.21 1.977 ;
      RECT 1.205 1.785 1.208 1.97 ;
      RECT 1.2 1.85 1.205 1.913 ;
      RECT 5.275 0.94 5.555 1.22 ;
      RECT 5.265 0.94 5.555 1.083 ;
      RECT 5.22 0.805 5.48 1.065 ;
      RECT 5.22 0.92 5.535 1.065 ;
      RECT 5.22 0.89 5.53 1.065 ;
      RECT 5.22 0.877 5.52 1.065 ;
      RECT 5.22 0.867 5.515 1.065 ;
      RECT 1.195 0.85 1.455 1.11 ;
      RECT 4.965 0.4 5.225 0.66 ;
      RECT 4.955 0.425 5.225 0.62 ;
      RECT 4.95 0.425 4.955 0.619 ;
      RECT 4.88 0.42 4.95 0.611 ;
      RECT 4.795 0.407 4.88 0.594 ;
      RECT 4.791 0.399 4.795 0.584 ;
      RECT 4.705 0.392 4.791 0.574 ;
      RECT 4.696 0.384 4.705 0.564 ;
      RECT 4.61 0.377 4.696 0.552 ;
      RECT 4.59 0.368 4.61 0.538 ;
      RECT 4.535 0.363 4.59 0.53 ;
      RECT 4.525 0.357 4.535 0.524 ;
      RECT 4.505 0.355 4.525 0.52 ;
      RECT 4.497 0.354 4.505 0.516 ;
      RECT 4.411 0.346 4.497 0.505 ;
      RECT 4.325 0.332 4.411 0.485 ;
      RECT 4.265 0.32 4.325 0.47 ;
      RECT 4.255 0.315 4.265 0.465 ;
      RECT 4.205 0.315 4.255 0.467 ;
      RECT 4.158 0.317 4.205 0.471 ;
      RECT 4.072 0.324 4.158 0.476 ;
      RECT 3.986 0.332 4.072 0.482 ;
      RECT 3.9 0.341 3.986 0.488 ;
      RECT 3.841 0.347 3.9 0.493 ;
      RECT 3.755 0.352 3.841 0.499 ;
      RECT 3.68 0.357 3.755 0.505 ;
      RECT 3.641 0.359 3.68 0.51 ;
      RECT 3.555 0.356 3.641 0.515 ;
      RECT 3.47 0.354 3.555 0.522 ;
      RECT 3.438 0.353 3.47 0.525 ;
      RECT 3.352 0.352 3.438 0.526 ;
      RECT 3.266 0.351 3.352 0.527 ;
      RECT 3.18 0.35 3.266 0.527 ;
      RECT 3.094 0.349 3.18 0.528 ;
      RECT 3.008 0.348 3.094 0.529 ;
      RECT 2.922 0.347 3.008 0.53 ;
      RECT 2.836 0.346 2.922 0.53 ;
      RECT 2.75 0.345 2.836 0.531 ;
      RECT 2.7 0.345 2.75 0.532 ;
      RECT 2.686 0.346 2.7 0.532 ;
      RECT 2.6 0.353 2.686 0.533 ;
      RECT 2.526 0.364 2.6 0.534 ;
      RECT 2.44 0.373 2.526 0.535 ;
      RECT 2.405 0.38 2.44 0.55 ;
      RECT 2.38 0.383 2.405 0.58 ;
      RECT 2.355 0.392 2.38 0.609 ;
      RECT 2.345 0.403 2.355 0.629 ;
      RECT 2.335 0.411 2.345 0.643 ;
      RECT 2.33 0.417 2.335 0.653 ;
      RECT 2.305 0.434 2.33 0.67 ;
      RECT 2.29 0.456 2.305 0.698 ;
      RECT 2.26 0.482 2.29 0.728 ;
      RECT 2.24 0.511 2.26 0.758 ;
      RECT 2.235 0.526 2.24 0.775 ;
      RECT 2.215 0.541 2.235 0.79 ;
      RECT 2.205 0.559 2.215 0.808 ;
      RECT 2.195 0.57 2.205 0.823 ;
      RECT 2.145 0.602 2.195 0.849 ;
      RECT 2.14 0.632 2.145 0.869 ;
      RECT 2.13 0.645 2.14 0.875 ;
      RECT 2.121 0.655 2.13 0.883 ;
      RECT 2.11 0.666 2.121 0.891 ;
      RECT 2.105 0.676 2.11 0.897 ;
      RECT 2.09 0.697 2.105 0.904 ;
      RECT 2.075 0.727 2.09 0.912 ;
      RECT 2.04 0.757 2.075 0.918 ;
      RECT 2.015 0.775 2.04 0.925 ;
      RECT 1.965 0.783 2.015 0.934 ;
      RECT 1.94 0.788 1.965 0.943 ;
      RECT 1.885 0.794 1.94 0.953 ;
      RECT 1.88 0.799 1.885 0.961 ;
      RECT 1.866 0.802 1.88 0.963 ;
      RECT 1.78 0.814 1.866 0.975 ;
      RECT 1.77 0.826 1.78 0.988 ;
      RECT 1.685 0.839 1.77 1 ;
      RECT 1.641 0.856 1.685 1.014 ;
      RECT 1.555 0.873 1.641 1.03 ;
      RECT 1.525 0.887 1.555 1.044 ;
      RECT 1.515 0.892 1.525 1.049 ;
      RECT 1.455 0.895 1.515 1.058 ;
      RECT 4.345 1.165 4.605 1.425 ;
      RECT 4.345 1.165 4.625 1.278 ;
      RECT 4.345 1.165 4.65 1.245 ;
      RECT 4.345 1.165 4.655 1.225 ;
      RECT 4.395 0.94 4.675 1.22 ;
      RECT 3.95 1.675 4.21 1.935 ;
      RECT 3.94 1.532 4.135 1.873 ;
      RECT 3.935 1.64 4.15 1.865 ;
      RECT 3.93 1.69 4.21 1.855 ;
      RECT 3.92 1.767 4.21 1.84 ;
      RECT 3.94 1.615 4.15 1.873 ;
      RECT 3.95 1.49 4.135 1.935 ;
      RECT 3.95 1.385 4.115 1.935 ;
      RECT 3.96 1.372 4.115 1.935 ;
      RECT 3.96 1.33 4.105 1.935 ;
      RECT 3.965 1.255 4.105 1.935 ;
      RECT 3.995 0.905 4.105 1.935 ;
      RECT 4 0.635 4.125 1.258 ;
      RECT 3.97 1.21 4.125 1.258 ;
      RECT 3.985 1.012 4.105 1.935 ;
      RECT 3.975 1.122 4.125 1.258 ;
      RECT 4 0.635 4.14 1.115 ;
      RECT 4 0.635 4.16 0.99 ;
      RECT 3.965 0.635 4.225 0.895 ;
      RECT 3.435 0.94 3.715 1.22 ;
      RECT 3.42 0.94 3.715 1.2 ;
      RECT 1.475 1.805 1.735 2.065 ;
      RECT 3.26 1.66 3.52 1.92 ;
      RECT 3.24 1.68 3.52 1.895 ;
      RECT 3.197 1.68 3.24 1.894 ;
      RECT 3.111 1.681 3.197 1.891 ;
      RECT 3.025 1.682 3.111 1.887 ;
      RECT 2.95 1.684 3.025 1.884 ;
      RECT 2.927 1.685 2.95 1.882 ;
      RECT 2.841 1.686 2.927 1.88 ;
      RECT 2.755 1.687 2.841 1.877 ;
      RECT 2.731 1.688 2.755 1.875 ;
      RECT 2.645 1.69 2.731 1.872 ;
      RECT 2.56 1.692 2.645 1.873 ;
      RECT 2.503 1.693 2.56 1.879 ;
      RECT 2.417 1.695 2.503 1.889 ;
      RECT 2.331 1.698 2.417 1.902 ;
      RECT 2.245 1.7 2.331 1.914 ;
      RECT 2.231 1.701 2.245 1.921 ;
      RECT 2.145 1.702 2.231 1.929 ;
      RECT 2.105 1.704 2.145 1.938 ;
      RECT 2.096 1.705 2.105 1.941 ;
      RECT 2.01 1.713 2.096 1.947 ;
      RECT 1.99 1.722 2.01 1.955 ;
      RECT 1.905 1.737 1.99 1.963 ;
      RECT 1.845 1.76 1.905 1.974 ;
      RECT 1.835 1.772 1.845 1.979 ;
      RECT 1.795 1.782 1.835 1.983 ;
      RECT 1.74 1.799 1.795 1.991 ;
      RECT 1.735 1.809 1.74 1.995 ;
      RECT 2.801 0.94 2.86 1.337 ;
      RECT 2.715 0.94 2.92 1.328 ;
      RECT 2.71 0.97 2.92 1.323 ;
      RECT 2.676 0.97 2.92 1.321 ;
      RECT 2.59 0.97 2.92 1.315 ;
      RECT 2.545 0.97 2.94 1.293 ;
      RECT 2.545 0.97 2.96 1.248 ;
      RECT 2.505 0.97 2.96 1.238 ;
      RECT 2.715 0.94 2.995 1.22 ;
      RECT 2.45 0.94 2.71 1.2 ;
      RECT 1.635 0.42 1.895 0.68 ;
      RECT 1.715 0.38 1.995 0.66 ;
      RECT 0.275 1.5 0.555 1.78 ;
      RECT 0.245 1.462 0.5 1.765 ;
      RECT 0.24 1.463 0.5 1.763 ;
      RECT 0.235 1.464 0.5 1.757 ;
      RECT 0.23 1.467 0.5 1.75 ;
      RECT 0.225 1.5 0.555 1.743 ;
      RECT 0.195 1.47 0.5 1.73 ;
      RECT 0.195 1.497 0.52 1.73 ;
      RECT 0.195 1.487 0.515 1.73 ;
      RECT 0.195 1.472 0.51 1.73 ;
      RECT 0.275 1.459 0.49 1.78 ;
      RECT 0.361 1.457 0.49 1.78 ;
      RECT 0.447 1.455 0.475 1.78 ;
    LAYER via1 ;
      RECT 9.09 0.79 9.24 0.94 ;
      RECT 8.97 1.36 9.12 1.51 ;
      RECT 7.89 1.055 8.04 1.205 ;
      RECT 7.555 1.775 7.705 1.925 ;
      RECT 7.475 0.615 7.625 0.765 ;
      RECT 6.04 1.01 6.19 1.16 ;
      RECT 5.275 0.86 5.425 1.01 ;
      RECT 5.02 0.455 5.17 0.605 ;
      RECT 4.4 1.22 4.55 1.37 ;
      RECT 4.02 0.69 4.17 0.84 ;
      RECT 4.005 1.73 4.155 1.88 ;
      RECT 3.475 0.995 3.625 1.145 ;
      RECT 3.315 1.715 3.465 1.865 ;
      RECT 2.505 0.995 2.655 1.145 ;
      RECT 1.69 0.475 1.84 0.625 ;
      RECT 1.53 1.86 1.68 2.01 ;
      RECT 1.295 1.515 1.445 1.665 ;
      RECT 1.25 0.905 1.4 1.055 ;
      RECT 0.25 1.525 0.4 1.675 ;
    LAYER met1 ;
      RECT 8.5 0.965 8.685 1.175 ;
      RECT 8.49 0.97 8.7 1.168 ;
      RECT 8.49 0.97 8.786 1.145 ;
      RECT 8.49 0.97 8.845 1.12 ;
      RECT 8.49 0.97 8.9 1.1 ;
      RECT 8.49 0.97 8.91 1.088 ;
      RECT 8.49 0.97 9.105 1.027 ;
      RECT 8.49 0.97 9.135 1.01 ;
      RECT 8.49 0.97 9.155 1 ;
      RECT 9.035 0.735 9.295 0.995 ;
      RECT 9.02 0.825 9.035 1.042 ;
      RECT 8.555 0.957 9.295 0.995 ;
      RECT 9.006 0.836 9.02 1.048 ;
      RECT 8.595 0.95 9.295 0.995 ;
      RECT 8.92 0.876 9.006 1.067 ;
      RECT 8.845 0.937 9.295 0.995 ;
      RECT 8.915 0.912 8.92 1.084 ;
      RECT 8.9 0.922 9.295 0.995 ;
      RECT 8.91 0.917 8.915 1.086 ;
      RECT 9.205 1.422 9.21 1.514 ;
      RECT 9.2 1.4 9.205 1.531 ;
      RECT 9.195 1.39 9.2 1.543 ;
      RECT 9.185 1.381 9.195 1.553 ;
      RECT 9.18 1.376 9.185 1.561 ;
      RECT 9.175 1.372 9.18 1.564 ;
      RECT 9.141 1.305 9.175 1.575 ;
      RECT 9.055 1.305 9.141 1.61 ;
      RECT 8.975 1.305 9.055 1.658 ;
      RECT 8.915 1.305 8.975 1.683 ;
      RECT 8.855 1.405 8.915 1.69 ;
      RECT 8.82 1.43 8.855 1.696 ;
      RECT 8.795 1.445 8.82 1.7 ;
      RECT 8.781 1.454 8.795 1.702 ;
      RECT 8.695 1.481 8.781 1.708 ;
      RECT 8.63 1.522 8.695 1.717 ;
      RECT 8.615 1.542 8.63 1.722 ;
      RECT 8.585 1.552 8.615 1.725 ;
      RECT 8.58 1.562 8.585 1.728 ;
      RECT 8.55 1.567 8.58 1.73 ;
      RECT 8.53 1.572 8.55 1.734 ;
      RECT 8.445 1.575 8.53 1.741 ;
      RECT 8.43 1.572 8.445 1.747 ;
      RECT 8.42 1.569 8.43 1.749 ;
      RECT 8.4 1.566 8.42 1.751 ;
      RECT 8.38 1.562 8.4 1.752 ;
      RECT 8.365 1.558 8.38 1.754 ;
      RECT 8.355 1.555 8.365 1.755 ;
      RECT 8.315 1.549 8.355 1.753 ;
      RECT 8.305 1.544 8.315 1.751 ;
      RECT 8.29 1.541 8.305 1.747 ;
      RECT 8.265 1.536 8.29 1.74 ;
      RECT 8.215 1.527 8.265 1.728 ;
      RECT 8.145 1.513 8.215 1.71 ;
      RECT 8.087 1.498 8.145 1.692 ;
      RECT 8.001 1.481 8.087 1.672 ;
      RECT 7.915 1.46 8.001 1.647 ;
      RECT 7.865 1.445 7.915 1.628 ;
      RECT 7.861 1.439 7.865 1.62 ;
      RECT 7.775 1.429 7.861 1.607 ;
      RECT 7.74 1.414 7.775 1.59 ;
      RECT 7.725 1.407 7.74 1.583 ;
      RECT 7.665 1.395 7.725 1.571 ;
      RECT 7.645 1.382 7.665 1.559 ;
      RECT 7.605 1.373 7.645 1.551 ;
      RECT 7.6 1.365 7.605 1.544 ;
      RECT 7.52 1.355 7.6 1.53 ;
      RECT 7.505 1.342 7.52 1.515 ;
      RECT 7.5 1.34 7.505 1.513 ;
      RECT 7.421 1.328 7.5 1.5 ;
      RECT 7.335 1.303 7.421 1.475 ;
      RECT 7.32 1.272 7.335 1.46 ;
      RECT 7.305 1.247 7.32 1.456 ;
      RECT 7.29 1.24 7.305 1.452 ;
      RECT 7.115 1.245 7.12 1.448 ;
      RECT 7.11 1.25 7.115 1.443 ;
      RECT 7.12 1.24 7.29 1.45 ;
      RECT 7.835 1 7.94 1.26 ;
      RECT 8.65 0.525 8.655 0.75 ;
      RECT 8.78 0.525 8.835 0.735 ;
      RECT 8.835 0.53 8.845 0.728 ;
      RECT 8.741 0.525 8.78 0.738 ;
      RECT 8.655 0.525 8.741 0.745 ;
      RECT 8.635 0.53 8.65 0.751 ;
      RECT 8.625 0.57 8.635 0.753 ;
      RECT 8.595 0.58 8.625 0.755 ;
      RECT 8.59 0.585 8.595 0.757 ;
      RECT 8.565 0.59 8.59 0.759 ;
      RECT 8.55 0.595 8.565 0.761 ;
      RECT 8.535 0.597 8.55 0.763 ;
      RECT 8.53 0.602 8.535 0.765 ;
      RECT 8.48 0.61 8.53 0.768 ;
      RECT 8.455 0.619 8.48 0.773 ;
      RECT 8.445 0.626 8.455 0.778 ;
      RECT 8.44 0.629 8.445 0.782 ;
      RECT 8.42 0.632 8.44 0.791 ;
      RECT 8.39 0.64 8.42 0.811 ;
      RECT 8.361 0.653 8.39 0.833 ;
      RECT 8.275 0.687 8.361 0.877 ;
      RECT 8.27 0.713 8.275 0.915 ;
      RECT 8.265 0.717 8.27 0.924 ;
      RECT 8.23 0.73 8.265 0.957 ;
      RECT 8.22 0.744 8.23 0.995 ;
      RECT 8.215 0.748 8.22 1.008 ;
      RECT 8.21 0.752 8.215 1.013 ;
      RECT 8.2 0.76 8.21 1.025 ;
      RECT 8.195 0.767 8.2 1.04 ;
      RECT 8.17 0.78 8.195 1.065 ;
      RECT 8.13 0.809 8.17 1.12 ;
      RECT 8.115 0.834 8.13 1.175 ;
      RECT 8.105 0.845 8.115 1.198 ;
      RECT 8.1 0.852 8.105 1.21 ;
      RECT 8.095 0.856 8.1 1.218 ;
      RECT 8.04 0.884 8.095 1.26 ;
      RECT 8.02 0.92 8.04 1.26 ;
      RECT 8.005 0.935 8.02 1.26 ;
      RECT 7.95 0.967 8.005 1.26 ;
      RECT 7.94 0.997 7.95 1.26 ;
      RECT 7.55 0.612 7.735 0.85 ;
      RECT 7.535 0.614 7.745 0.845 ;
      RECT 7.42 0.56 7.68 0.82 ;
      RECT 7.415 0.597 7.68 0.774 ;
      RECT 7.41 0.607 7.68 0.771 ;
      RECT 7.405 0.647 7.745 0.765 ;
      RECT 7.4 0.68 7.745 0.755 ;
      RECT 7.41 0.622 7.76 0.693 ;
      RECT 7.707 1.72 7.72 2.25 ;
      RECT 7.621 1.72 7.72 2.249 ;
      RECT 7.621 1.72 7.725 2.248 ;
      RECT 7.535 1.72 7.725 2.246 ;
      RECT 7.53 1.72 7.725 2.243 ;
      RECT 7.53 1.72 7.735 2.241 ;
      RECT 7.525 2.012 7.735 2.238 ;
      RECT 7.525 2.022 7.74 2.235 ;
      RECT 7.525 2.09 7.745 2.231 ;
      RECT 7.515 2.095 7.745 2.23 ;
      RECT 7.515 2.187 7.75 2.227 ;
      RECT 7.5 1.72 7.76 1.98 ;
      RECT 6.73 0.71 6.775 2.245 ;
      RECT 6.93 0.71 6.96 0.925 ;
      RECT 5.305 0.45 5.425 0.66 ;
      RECT 4.965 0.4 5.225 0.66 ;
      RECT 4.965 0.445 5.26 0.65 ;
      RECT 6.97 0.726 6.975 0.78 ;
      RECT 6.965 0.719 6.97 0.913 ;
      RECT 6.96 0.713 6.965 0.92 ;
      RECT 6.915 0.71 6.93 0.933 ;
      RECT 6.91 0.71 6.915 0.955 ;
      RECT 6.905 0.71 6.91 1.003 ;
      RECT 6.9 0.71 6.905 1.023 ;
      RECT 6.89 0.71 6.9 1.13 ;
      RECT 6.885 0.71 6.89 1.193 ;
      RECT 6.88 0.71 6.885 1.25 ;
      RECT 6.875 0.71 6.88 1.258 ;
      RECT 6.86 0.71 6.875 1.365 ;
      RECT 6.85 0.71 6.86 1.5 ;
      RECT 6.84 0.71 6.85 1.61 ;
      RECT 6.83 0.71 6.84 1.667 ;
      RECT 6.825 0.71 6.83 1.707 ;
      RECT 6.82 0.71 6.825 1.743 ;
      RECT 6.81 0.71 6.82 1.783 ;
      RECT 6.805 0.71 6.81 1.825 ;
      RECT 6.785 0.71 6.805 1.89 ;
      RECT 6.79 2.035 6.795 2.215 ;
      RECT 6.785 2.017 6.79 2.223 ;
      RECT 6.78 0.71 6.785 1.953 ;
      RECT 6.78 1.997 6.785 2.23 ;
      RECT 6.775 0.71 6.78 2.24 ;
      RECT 6.72 0.71 6.73 1.01 ;
      RECT 6.725 1.257 6.73 2.245 ;
      RECT 6.72 1.322 6.725 2.245 ;
      RECT 6.715 0.711 6.72 1 ;
      RECT 6.71 1.387 6.72 2.245 ;
      RECT 6.705 0.712 6.715 0.99 ;
      RECT 6.695 1.5 6.71 2.245 ;
      RECT 6.7 0.713 6.705 0.98 ;
      RECT 6.68 0.714 6.7 0.958 ;
      RECT 6.685 1.597 6.695 2.245 ;
      RECT 6.68 1.672 6.685 2.245 ;
      RECT 6.67 0.713 6.68 0.935 ;
      RECT 6.675 1.715 6.68 2.245 ;
      RECT 6.67 1.742 6.675 2.245 ;
      RECT 6.66 0.711 6.67 0.923 ;
      RECT 6.665 1.785 6.67 2.245 ;
      RECT 6.66 1.812 6.665 2.245 ;
      RECT 6.65 0.71 6.66 0.91 ;
      RECT 6.655 1.827 6.66 2.245 ;
      RECT 6.615 1.885 6.655 2.245 ;
      RECT 6.645 0.709 6.65 0.895 ;
      RECT 6.64 0.707 6.645 0.888 ;
      RECT 6.63 0.704 6.64 0.878 ;
      RECT 6.625 0.701 6.63 0.863 ;
      RECT 6.61 0.697 6.625 0.856 ;
      RECT 6.605 1.94 6.615 2.245 ;
      RECT 6.605 0.694 6.61 0.851 ;
      RECT 6.59 0.69 6.605 0.845 ;
      RECT 6.6 1.957 6.605 2.245 ;
      RECT 6.59 2.02 6.6 2.245 ;
      RECT 6.51 0.675 6.59 0.825 ;
      RECT 6.585 2.027 6.59 2.24 ;
      RECT 6.58 2.035 6.585 2.23 ;
      RECT 6.5 0.661 6.51 0.809 ;
      RECT 6.485 0.657 6.5 0.807 ;
      RECT 6.475 0.652 6.485 0.803 ;
      RECT 6.45 0.645 6.475 0.795 ;
      RECT 6.445 0.64 6.45 0.79 ;
      RECT 6.435 0.64 6.445 0.788 ;
      RECT 6.425 0.638 6.435 0.786 ;
      RECT 6.395 0.63 6.425 0.78 ;
      RECT 6.38 0.622 6.395 0.773 ;
      RECT 6.36 0.617 6.38 0.766 ;
      RECT 6.355 0.613 6.36 0.761 ;
      RECT 6.325 0.606 6.355 0.755 ;
      RECT 6.3 0.597 6.325 0.745 ;
      RECT 6.27 0.59 6.3 0.737 ;
      RECT 6.245 0.58 6.27 0.728 ;
      RECT 6.23 0.572 6.245 0.722 ;
      RECT 6.205 0.567 6.23 0.717 ;
      RECT 6.195 0.563 6.205 0.712 ;
      RECT 6.175 0.558 6.195 0.707 ;
      RECT 6.14 0.553 6.175 0.7 ;
      RECT 6.08 0.548 6.14 0.693 ;
      RECT 6.067 0.544 6.08 0.691 ;
      RECT 5.981 0.539 6.067 0.688 ;
      RECT 5.895 0.529 5.981 0.684 ;
      RECT 5.854 0.522 5.895 0.681 ;
      RECT 5.768 0.515 5.854 0.678 ;
      RECT 5.682 0.505 5.768 0.674 ;
      RECT 5.596 0.495 5.682 0.669 ;
      RECT 5.51 0.485 5.596 0.665 ;
      RECT 5.5 0.47 5.51 0.663 ;
      RECT 5.49 0.455 5.5 0.663 ;
      RECT 5.425 0.45 5.49 0.662 ;
      RECT 5.26 0.447 5.305 0.655 ;
      RECT 6.505 1.352 6.51 1.543 ;
      RECT 6.5 1.347 6.505 1.55 ;
      RECT 6.486 1.345 6.5 1.556 ;
      RECT 6.4 1.345 6.486 1.558 ;
      RECT 6.396 1.345 6.4 1.561 ;
      RECT 6.31 1.345 6.396 1.579 ;
      RECT 6.3 1.35 6.31 1.598 ;
      RECT 6.29 1.405 6.3 1.602 ;
      RECT 6.265 1.42 6.29 1.609 ;
      RECT 6.225 1.44 6.265 1.622 ;
      RECT 6.22 1.452 6.225 1.632 ;
      RECT 6.205 1.458 6.22 1.637 ;
      RECT 6.2 1.463 6.205 1.641 ;
      RECT 6.18 1.47 6.2 1.646 ;
      RECT 6.11 1.495 6.18 1.663 ;
      RECT 6.07 1.523 6.11 1.683 ;
      RECT 6.065 1.533 6.07 1.691 ;
      RECT 6.045 1.54 6.065 1.693 ;
      RECT 6.04 1.547 6.045 1.696 ;
      RECT 6.01 1.555 6.04 1.699 ;
      RECT 6.005 1.56 6.01 1.703 ;
      RECT 5.931 1.564 6.005 1.711 ;
      RECT 5.845 1.573 5.931 1.727 ;
      RECT 5.841 1.578 5.845 1.736 ;
      RECT 5.755 1.583 5.841 1.746 ;
      RECT 5.715 1.591 5.755 1.758 ;
      RECT 5.665 1.597 5.715 1.765 ;
      RECT 5.58 1.606 5.665 1.78 ;
      RECT 5.505 1.617 5.58 1.798 ;
      RECT 5.47 1.624 5.505 1.808 ;
      RECT 5.395 1.632 5.47 1.813 ;
      RECT 5.34 1.641 5.395 1.813 ;
      RECT 5.315 1.646 5.34 1.811 ;
      RECT 5.305 1.649 5.315 1.809 ;
      RECT 5.27 1.651 5.305 1.807 ;
      RECT 5.24 1.653 5.27 1.803 ;
      RECT 5.195 1.652 5.24 1.799 ;
      RECT 5.175 1.647 5.195 1.796 ;
      RECT 5.125 1.632 5.175 1.793 ;
      RECT 5.115 1.617 5.125 1.788 ;
      RECT 5.065 1.602 5.115 1.778 ;
      RECT 5.015 1.577 5.065 1.758 ;
      RECT 5.005 1.562 5.015 1.74 ;
      RECT 5 1.56 5.005 1.734 ;
      RECT 4.98 1.555 5 1.729 ;
      RECT 4.975 1.547 4.98 1.723 ;
      RECT 4.96 1.541 4.975 1.716 ;
      RECT 4.955 1.536 4.96 1.708 ;
      RECT 4.935 1.531 4.955 1.7 ;
      RECT 4.92 1.524 4.935 1.693 ;
      RECT 4.905 1.518 4.92 1.684 ;
      RECT 4.9 1.512 4.905 1.677 ;
      RECT 4.855 1.487 4.9 1.663 ;
      RECT 4.84 1.457 4.855 1.645 ;
      RECT 4.825 1.44 4.84 1.636 ;
      RECT 4.8 1.42 4.825 1.624 ;
      RECT 4.76 1.39 4.8 1.604 ;
      RECT 4.75 1.36 4.76 1.589 ;
      RECT 4.735 1.35 4.75 1.582 ;
      RECT 4.68 1.315 4.735 1.561 ;
      RECT 4.665 1.278 4.68 1.54 ;
      RECT 4.655 1.265 4.665 1.532 ;
      RECT 4.605 1.235 4.655 1.514 ;
      RECT 4.59 1.165 4.605 1.495 ;
      RECT 4.545 1.165 4.59 1.478 ;
      RECT 4.52 1.165 4.545 1.46 ;
      RECT 4.51 1.165 4.52 1.453 ;
      RECT 4.431 1.165 4.51 1.446 ;
      RECT 4.345 1.165 4.431 1.438 ;
      RECT 4.33 1.197 4.345 1.433 ;
      RECT 4.255 1.207 4.33 1.429 ;
      RECT 4.235 1.217 4.255 1.424 ;
      RECT 4.21 1.217 4.235 1.421 ;
      RECT 4.2 1.207 4.21 1.42 ;
      RECT 4.19 1.18 4.2 1.419 ;
      RECT 4.15 1.175 4.19 1.417 ;
      RECT 4.105 1.175 4.15 1.413 ;
      RECT 4.08 1.175 4.105 1.408 ;
      RECT 4.03 1.175 4.08 1.395 ;
      RECT 3.99 1.18 4 1.38 ;
      RECT 4 1.175 4.03 1.385 ;
      RECT 5.985 0.955 6.245 1.215 ;
      RECT 5.98 0.977 6.245 1.173 ;
      RECT 5.22 0.805 5.44 1.17 ;
      RECT 5.202 0.892 5.44 1.169 ;
      RECT 5.185 0.897 5.44 1.166 ;
      RECT 5.185 0.897 5.46 1.165 ;
      RECT 5.155 0.907 5.46 1.163 ;
      RECT 5.15 0.922 5.46 1.159 ;
      RECT 5.15 0.922 5.465 1.158 ;
      RECT 5.145 0.98 5.465 1.156 ;
      RECT 5.145 0.98 5.475 1.153 ;
      RECT 5.14 1.045 5.475 1.148 ;
      RECT 5.22 0.805 5.48 1.065 ;
      RECT 3.965 0.635 4.225 0.895 ;
      RECT 3.965 0.678 4.311 0.869 ;
      RECT 3.965 0.678 4.355 0.868 ;
      RECT 3.965 0.678 4.375 0.866 ;
      RECT 3.965 0.678 4.475 0.865 ;
      RECT 3.965 0.678 4.495 0.863 ;
      RECT 3.965 0.678 4.505 0.858 ;
      RECT 4.375 0.645 4.565 0.855 ;
      RECT 4.375 0.647 4.57 0.853 ;
      RECT 4.365 0.652 4.575 0.845 ;
      RECT 4.311 0.676 4.575 0.845 ;
      RECT 4.355 0.67 4.365 0.867 ;
      RECT 4.365 0.65 4.57 0.853 ;
      RECT 3.32 1.71 3.525 1.94 ;
      RECT 3.26 1.66 3.315 1.92 ;
      RECT 3.32 1.66 3.52 1.94 ;
      RECT 4.29 1.975 4.295 2.002 ;
      RECT 4.28 1.885 4.29 2.007 ;
      RECT 4.275 1.807 4.28 2.013 ;
      RECT 4.265 1.797 4.275 2.02 ;
      RECT 4.26 1.787 4.265 2.026 ;
      RECT 4.25 1.782 4.26 2.028 ;
      RECT 4.235 1.774 4.25 2.036 ;
      RECT 4.22 1.765 4.235 2.048 ;
      RECT 4.21 1.757 4.22 2.058 ;
      RECT 4.175 1.675 4.21 2.076 ;
      RECT 4.14 1.675 4.175 2.095 ;
      RECT 4.125 1.675 4.14 2.103 ;
      RECT 4.07 1.675 4.125 2.103 ;
      RECT 4.036 1.675 4.07 2.094 ;
      RECT 3.95 1.675 4.036 2.07 ;
      RECT 3.94 1.735 3.95 2.052 ;
      RECT 3.9 1.737 3.94 2.043 ;
      RECT 3.895 1.739 3.9 2.033 ;
      RECT 3.875 1.741 3.895 2.028 ;
      RECT 3.865 1.744 3.875 2.023 ;
      RECT 3.855 1.745 3.865 2.018 ;
      RECT 3.831 1.746 3.855 2.01 ;
      RECT 3.745 1.751 3.831 1.988 ;
      RECT 3.69 1.75 3.745 1.961 ;
      RECT 3.675 1.743 3.69 1.948 ;
      RECT 3.64 1.738 3.675 1.944 ;
      RECT 3.585 1.73 3.64 1.943 ;
      RECT 3.525 1.717 3.585 1.941 ;
      RECT 3.315 1.66 3.32 1.928 ;
      RECT 3.39 1.03 3.575 1.24 ;
      RECT 3.38 1.035 3.59 1.233 ;
      RECT 3.42 0.94 3.68 1.2 ;
      RECT 3.375 1.097 3.68 1.123 ;
      RECT 2.72 0.89 2.725 1.69 ;
      RECT 2.665 0.94 2.695 1.69 ;
      RECT 2.655 0.94 2.66 1.25 ;
      RECT 2.64 0.94 2.645 1.245 ;
      RECT 2.185 0.985 2.2 1.2 ;
      RECT 2.115 0.985 2.2 1.195 ;
      RECT 3.38 0.565 3.45 0.775 ;
      RECT 3.45 0.572 3.46 0.77 ;
      RECT 3.346 0.565 3.38 0.782 ;
      RECT 3.26 0.565 3.346 0.806 ;
      RECT 3.25 0.57 3.26 0.825 ;
      RECT 3.245 0.582 3.25 0.828 ;
      RECT 3.23 0.597 3.245 0.832 ;
      RECT 3.225 0.615 3.23 0.836 ;
      RECT 3.185 0.625 3.225 0.845 ;
      RECT 3.17 0.632 3.185 0.857 ;
      RECT 3.155 0.637 3.17 0.862 ;
      RECT 3.14 0.64 3.155 0.867 ;
      RECT 3.13 0.642 3.14 0.871 ;
      RECT 3.095 0.649 3.13 0.879 ;
      RECT 3.06 0.657 3.095 0.893 ;
      RECT 3.05 0.663 3.06 0.902 ;
      RECT 3.045 0.665 3.05 0.904 ;
      RECT 3.025 0.668 3.045 0.91 ;
      RECT 2.995 0.675 3.025 0.921 ;
      RECT 2.985 0.681 2.995 0.928 ;
      RECT 2.96 0.684 2.985 0.935 ;
      RECT 2.95 0.688 2.96 0.943 ;
      RECT 2.945 0.689 2.95 0.965 ;
      RECT 2.94 0.69 2.945 0.98 ;
      RECT 2.935 0.691 2.94 0.995 ;
      RECT 2.93 0.692 2.935 1.01 ;
      RECT 2.925 0.693 2.93 1.04 ;
      RECT 2.915 0.695 2.925 1.073 ;
      RECT 2.9 0.699 2.915 1.12 ;
      RECT 2.89 0.702 2.9 1.165 ;
      RECT 2.885 0.705 2.89 1.193 ;
      RECT 2.875 0.707 2.885 1.22 ;
      RECT 2.87 0.71 2.875 1.255 ;
      RECT 2.84 0.715 2.87 1.313 ;
      RECT 2.835 0.72 2.84 1.398 ;
      RECT 2.83 0.722 2.835 1.433 ;
      RECT 2.825 0.724 2.83 1.515 ;
      RECT 2.82 0.726 2.825 1.603 ;
      RECT 2.81 0.728 2.82 1.685 ;
      RECT 2.795 0.742 2.81 1.69 ;
      RECT 2.76 0.787 2.795 1.69 ;
      RECT 2.75 0.827 2.76 1.69 ;
      RECT 2.735 0.855 2.75 1.69 ;
      RECT 2.73 0.872 2.735 1.69 ;
      RECT 2.725 0.88 2.73 1.69 ;
      RECT 2.715 0.895 2.72 1.69 ;
      RECT 2.71 0.902 2.715 1.69 ;
      RECT 2.7 0.922 2.71 1.69 ;
      RECT 2.695 0.935 2.7 1.69 ;
      RECT 2.66 0.94 2.665 1.275 ;
      RECT 2.645 1.33 2.665 1.69 ;
      RECT 2.645 0.94 2.655 1.248 ;
      RECT 2.64 1.37 2.645 1.69 ;
      RECT 2.59 0.94 2.64 1.243 ;
      RECT 2.635 1.407 2.64 1.69 ;
      RECT 2.625 1.43 2.635 1.69 ;
      RECT 2.62 1.475 2.625 1.69 ;
      RECT 2.61 1.485 2.62 1.683 ;
      RECT 2.536 0.94 2.59 1.237 ;
      RECT 2.45 0.94 2.536 1.23 ;
      RECT 2.401 0.987 2.45 1.223 ;
      RECT 2.315 0.995 2.401 1.216 ;
      RECT 2.3 0.992 2.315 1.211 ;
      RECT 2.286 0.985 2.3 1.21 ;
      RECT 2.2 0.985 2.286 1.205 ;
      RECT 2.105 0.99 2.115 1.19 ;
      RECT 1.695 0.42 1.71 0.82 ;
      RECT 1.89 0.42 1.895 0.68 ;
      RECT 1.635 0.42 1.68 0.68 ;
      RECT 2.09 1.725 2.095 1.93 ;
      RECT 2.085 1.715 2.09 1.935 ;
      RECT 2.08 1.702 2.085 1.94 ;
      RECT 2.075 1.682 2.08 1.94 ;
      RECT 2.05 1.635 2.075 1.94 ;
      RECT 2.015 1.55 2.05 1.94 ;
      RECT 2.01 1.487 2.015 1.94 ;
      RECT 2.005 1.472 2.01 1.94 ;
      RECT 1.99 1.432 2.005 1.94 ;
      RECT 1.985 1.407 1.99 1.94 ;
      RECT 1.975 1.39 1.985 1.94 ;
      RECT 1.94 1.312 1.975 1.94 ;
      RECT 1.935 1.255 1.94 1.94 ;
      RECT 1.93 1.242 1.935 1.94 ;
      RECT 1.92 1.22 1.93 1.94 ;
      RECT 1.91 1.185 1.92 1.94 ;
      RECT 1.9 1.155 1.91 1.94 ;
      RECT 1.89 1.07 1.9 1.583 ;
      RECT 1.897 1.715 1.9 1.94 ;
      RECT 1.895 1.725 1.897 1.94 ;
      RECT 1.885 1.735 1.895 1.935 ;
      RECT 1.88 0.42 1.89 0.815 ;
      RECT 1.885 0.947 1.89 1.558 ;
      RECT 1.88 0.845 1.885 1.541 ;
      RECT 1.87 0.42 1.88 1.517 ;
      RECT 1.865 0.42 1.87 1.488 ;
      RECT 1.86 0.42 1.865 1.478 ;
      RECT 1.84 0.42 1.86 1.44 ;
      RECT 1.835 0.42 1.84 1.398 ;
      RECT 1.83 0.42 1.835 1.378 ;
      RECT 1.8 0.42 1.83 1.328 ;
      RECT 1.79 0.42 1.8 1.275 ;
      RECT 1.785 0.42 1.79 1.248 ;
      RECT 1.78 0.42 1.785 1.233 ;
      RECT 1.77 0.42 1.78 1.21 ;
      RECT 1.76 0.42 1.77 1.185 ;
      RECT 1.755 0.42 1.76 1.125 ;
      RECT 1.745 0.42 1.755 1.063 ;
      RECT 1.74 0.42 1.745 0.983 ;
      RECT 1.735 0.42 1.74 0.948 ;
      RECT 1.73 0.42 1.735 0.923 ;
      RECT 1.725 0.42 1.73 0.908 ;
      RECT 1.72 0.42 1.725 0.878 ;
      RECT 1.715 0.42 1.72 0.855 ;
      RECT 1.71 0.42 1.715 0.828 ;
      RECT 1.68 0.42 1.695 0.815 ;
      RECT 0.835 1.955 1.02 2.165 ;
      RECT 0.825 1.96 1.035 2.158 ;
      RECT 0.825 1.96 1.055 2.13 ;
      RECT 0.825 1.96 1.07 2.109 ;
      RECT 0.825 1.96 1.085 2.107 ;
      RECT 0.825 1.96 1.095 2.106 ;
      RECT 0.825 1.96 1.125 2.103 ;
      RECT 1.475 1.805 1.735 2.065 ;
      RECT 1.435 1.852 1.735 2.048 ;
      RECT 1.426 1.86 1.435 2.051 ;
      RECT 1.02 1.953 1.735 2.048 ;
      RECT 1.34 1.878 1.426 2.058 ;
      RECT 1.035 1.95 1.735 2.048 ;
      RECT 1.281 1.9 1.34 2.07 ;
      RECT 1.055 1.946 1.735 2.048 ;
      RECT 1.195 1.912 1.281 2.081 ;
      RECT 1.07 1.942 1.735 2.048 ;
      RECT 1.14 1.925 1.195 2.093 ;
      RECT 1.085 1.94 1.735 2.048 ;
      RECT 1.125 1.931 1.14 2.099 ;
      RECT 1.095 1.936 1.735 2.048 ;
      RECT 1.24 1.46 1.5 1.72 ;
      RECT 1.24 1.48 1.61 1.69 ;
      RECT 1.24 1.485 1.62 1.685 ;
      RECT 1.431 0.899 1.51 1.13 ;
      RECT 1.345 0.902 1.56 1.125 ;
      RECT 1.34 0.902 1.56 1.12 ;
      RECT 1.34 0.907 1.57 1.118 ;
      RECT 1.315 0.907 1.57 1.115 ;
      RECT 1.315 0.915 1.58 1.113 ;
      RECT 1.195 0.85 1.455 1.11 ;
      RECT 1.195 0.897 1.505 1.11 ;
      RECT 0.45 1.47 0.455 1.73 ;
      RECT 0.28 1.24 0.285 1.73 ;
      RECT 0.165 1.48 0.17 1.705 ;
      RECT 0.875 0.575 0.88 0.785 ;
      RECT 0.88 0.58 0.895 0.78 ;
      RECT 0.815 0.575 0.875 0.793 ;
      RECT 0.8 0.575 0.815 0.803 ;
      RECT 0.75 0.575 0.8 0.82 ;
      RECT 0.73 0.575 0.75 0.843 ;
      RECT 0.715 0.575 0.73 0.855 ;
      RECT 0.695 0.575 0.715 0.865 ;
      RECT 0.685 0.58 0.695 0.874 ;
      RECT 0.68 0.59 0.685 0.879 ;
      RECT 0.675 0.602 0.68 0.883 ;
      RECT 0.665 0.625 0.675 0.888 ;
      RECT 0.66 0.64 0.665 0.892 ;
      RECT 0.655 0.657 0.66 0.895 ;
      RECT 0.65 0.665 0.655 0.898 ;
      RECT 0.64 0.67 0.65 0.902 ;
      RECT 0.635 0.677 0.64 0.907 ;
      RECT 0.625 0.682 0.635 0.911 ;
      RECT 0.6 0.694 0.625 0.922 ;
      RECT 0.58 0.711 0.6 0.938 ;
      RECT 0.555 0.728 0.58 0.96 ;
      RECT 0.52 0.751 0.555 1.018 ;
      RECT 0.5 0.773 0.52 1.08 ;
      RECT 0.495 0.783 0.5 1.115 ;
      RECT 0.485 0.79 0.495 1.153 ;
      RECT 0.48 0.797 0.485 1.173 ;
      RECT 0.475 0.808 0.48 1.21 ;
      RECT 0.47 0.816 0.475 1.275 ;
      RECT 0.46 0.827 0.47 1.328 ;
      RECT 0.455 0.845 0.46 1.398 ;
      RECT 0.45 0.855 0.455 1.435 ;
      RECT 0.445 0.865 0.45 1.73 ;
      RECT 0.44 0.877 0.445 1.73 ;
      RECT 0.435 0.887 0.44 1.73 ;
      RECT 0.425 0.897 0.435 1.73 ;
      RECT 0.415 0.92 0.425 1.73 ;
      RECT 0.4 0.955 0.415 1.73 ;
      RECT 0.36 1.017 0.4 1.73 ;
      RECT 0.355 1.07 0.36 1.73 ;
      RECT 0.33 1.105 0.355 1.73 ;
      RECT 0.315 1.15 0.33 1.73 ;
      RECT 0.31 1.172 0.315 1.73 ;
      RECT 0.3 1.185 0.31 1.73 ;
      RECT 0.29 1.21 0.3 1.73 ;
      RECT 0.285 1.232 0.29 1.73 ;
      RECT 0.26 1.27 0.28 1.73 ;
      RECT 0.22 1.327 0.26 1.73 ;
      RECT 0.215 1.377 0.22 1.73 ;
      RECT 0.21 1.395 0.215 1.73 ;
      RECT 0.205 1.407 0.21 1.73 ;
      RECT 0.195 1.425 0.205 1.73 ;
      RECT 0.185 1.445 0.195 1.705 ;
      RECT 0.18 1.462 0.185 1.705 ;
      RECT 0.17 1.475 0.18 1.705 ;
      RECT 0.14 1.485 0.165 1.705 ;
      RECT 0.13 1.492 0.14 1.705 ;
      RECT 0.115 1.502 0.13 1.7 ;
      RECT 0 -0.24 9.66 0.24 ;
      RECT 0 2.48 9.66 2.96 ;
    LAYER mcon ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 8.975 1.375 9.145 1.545 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 8.655 0.545 8.825 0.715 ;
      RECT 8.51 0.985 8.68 1.155 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 7.9 1.025 8.07 1.195 ;
      RECT 7.555 0.66 7.725 0.83 ;
      RECT 7.545 2.02 7.715 2.19 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.13 1.26 7.3 1.43 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 6.78 0.735 6.95 0.905 ;
      RECT 6.6 2.05 6.77 2.22 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.32 1.365 6.49 1.535 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6 0.99 6.17 1.16 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.31 0.47 5.48 0.64 ;
      RECT 5.235 0.94 5.405 1.11 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.385 0.665 4.555 0.835 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.045 1.86 4.215 2.03 ;
      RECT 4.01 1.195 4.18 1.365 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 3.4 1.05 3.57 1.22 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.33 1.75 3.5 1.92 ;
      RECT 3.27 0.585 3.44 0.755 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.63 1.5 2.8 1.67 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.125 1.005 2.295 1.175 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 1.905 1.75 2.075 1.92 ;
      RECT 1.7 0.63 1.87 0.8 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.43 1.5 1.6 1.67 ;
      RECT 1.39 0.93 1.56 1.1 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 0.845 1.975 1.015 2.145 ;
      RECT 0.705 0.595 0.875 0.765 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.135 1.515 0.305 1.685 ;
    LAYER li ;
      RECT 8.13 -0.085 8.3 0.585 ;
      RECT 6.17 -0.085 6.34 0.585 ;
      RECT 3.73 -0.085 3.9 0.585 ;
      RECT 2.77 -0.085 2.94 0.585 ;
      RECT 2.25 -0.085 2.42 0.585 ;
      RECT 1.29 -0.085 1.46 0.585 ;
      RECT 0.33 -0.085 0.5 0.585 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 9.09 2.135 9.26 2.805 ;
      RECT 8.13 2.135 8.3 2.805 ;
      RECT 5.69 2.135 5.86 2.805 ;
      RECT 4.69 2.135 4.86 2.805 ;
      RECT 3.73 2.135 3.9 2.805 ;
      RECT 1.29 2.135 1.46 2.805 ;
      RECT 8.655 0.475 9.385 0.715 ;
      RECT 9.197 0.27 9.385 0.715 ;
      RECT 9.025 0.282 9.4 0.709 ;
      RECT 8.94 0.297 9.42 0.694 ;
      RECT 8.94 0.312 9.425 0.684 ;
      RECT 8.895 0.332 9.44 0.676 ;
      RECT 8.872 0.367 9.455 0.63 ;
      RECT 8.786 0.39 9.46 0.59 ;
      RECT 8.786 0.408 9.47 0.56 ;
      RECT 8.655 0.477 9.475 0.523 ;
      RECT 8.7 0.42 9.47 0.56 ;
      RECT 8.786 0.372 9.455 0.63 ;
      RECT 8.872 0.341 9.44 0.676 ;
      RECT 8.895 0.322 9.425 0.684 ;
      RECT 8.94 0.295 9.4 0.709 ;
      RECT 9.025 0.277 9.385 0.715 ;
      RECT 9.111 0.271 9.385 0.715 ;
      RECT 9.197 0.266 9.33 0.715 ;
      RECT 9.283 0.261 9.33 0.715 ;
      RECT 8.975 1.159 9.145 1.545 ;
      RECT 8.97 1.159 9.145 1.54 ;
      RECT 8.945 1.159 9.145 1.505 ;
      RECT 8.945 1.187 9.155 1.495 ;
      RECT 8.925 1.187 9.155 1.455 ;
      RECT 8.92 1.187 9.155 1.428 ;
      RECT 8.92 1.205 9.16 1.42 ;
      RECT 8.865 1.205 9.16 1.355 ;
      RECT 8.865 1.222 9.17 1.338 ;
      RECT 8.855 1.222 9.17 1.278 ;
      RECT 8.855 1.239 9.175 1.275 ;
      RECT 8.85 1.075 9.02 1.253 ;
      RECT 8.85 1.109 9.106 1.253 ;
      RECT 8.845 1.875 8.85 1.888 ;
      RECT 8.84 1.77 8.845 1.893 ;
      RECT 8.815 1.63 8.84 1.908 ;
      RECT 8.78 1.581 8.815 1.94 ;
      RECT 8.775 1.549 8.78 1.96 ;
      RECT 8.77 1.54 8.775 1.96 ;
      RECT 8.69 1.505 8.77 1.96 ;
      RECT 8.627 1.475 8.69 1.96 ;
      RECT 8.541 1.463 8.627 1.96 ;
      RECT 8.455 1.449 8.541 1.96 ;
      RECT 8.375 1.436 8.455 1.946 ;
      RECT 8.34 1.428 8.375 1.926 ;
      RECT 8.33 1.425 8.34 1.917 ;
      RECT 8.3 1.42 8.33 1.904 ;
      RECT 8.25 1.395 8.3 1.88 ;
      RECT 8.236 1.369 8.25 1.862 ;
      RECT 8.15 1.329 8.236 1.838 ;
      RECT 8.105 1.277 8.15 1.807 ;
      RECT 8.095 1.252 8.105 1.794 ;
      RECT 8.09 1.033 8.095 1.055 ;
      RECT 8.085 1.235 8.095 1.79 ;
      RECT 8.085 1.031 8.09 1.145 ;
      RECT 8.075 1.027 8.085 1.786 ;
      RECT 8.031 1.025 8.075 1.774 ;
      RECT 7.945 1.025 8.031 1.745 ;
      RECT 7.915 1.025 7.945 1.718 ;
      RECT 7.9 1.025 7.915 1.706 ;
      RECT 7.86 1.037 7.9 1.691 ;
      RECT 7.84 1.056 7.86 1.67 ;
      RECT 7.83 1.066 7.84 1.654 ;
      RECT 7.82 1.072 7.83 1.643 ;
      RECT 7.8 1.082 7.82 1.626 ;
      RECT 7.795 1.091 7.8 1.613 ;
      RECT 7.79 1.095 7.795 1.563 ;
      RECT 7.78 1.101 7.79 1.48 ;
      RECT 7.775 1.105 7.78 1.394 ;
      RECT 7.77 1.125 7.775 1.331 ;
      RECT 7.765 1.148 7.77 1.278 ;
      RECT 7.76 1.166 7.765 1.223 ;
      RECT 8.37 0.985 8.54 1.245 ;
      RECT 8.54 0.95 8.585 1.231 ;
      RECT 8.501 0.952 8.59 1.214 ;
      RECT 8.39 0.969 8.676 1.185 ;
      RECT 8.39 0.984 8.68 1.157 ;
      RECT 8.39 0.965 8.59 1.214 ;
      RECT 8.415 0.953 8.54 1.245 ;
      RECT 8.501 0.951 8.585 1.231 ;
      RECT 7.555 0.34 7.725 0.83 ;
      RECT 7.555 0.34 7.76 0.81 ;
      RECT 7.69 0.26 7.8 0.77 ;
      RECT 7.671 0.264 7.82 0.74 ;
      RECT 7.585 0.272 7.84 0.723 ;
      RECT 7.585 0.278 7.845 0.713 ;
      RECT 7.585 0.287 7.865 0.701 ;
      RECT 7.56 0.312 7.895 0.679 ;
      RECT 7.56 0.332 7.9 0.659 ;
      RECT 7.555 0.345 7.91 0.639 ;
      RECT 7.555 0.412 7.915 0.62 ;
      RECT 7.555 0.545 7.92 0.607 ;
      RECT 7.55 0.35 7.91 0.44 ;
      RECT 7.56 0.307 7.865 0.701 ;
      RECT 7.671 0.262 7.8 0.77 ;
      RECT 7.545 2.015 7.845 2.27 ;
      RECT 7.63 1.981 7.845 2.27 ;
      RECT 7.63 1.984 7.85 2.13 ;
      RECT 7.565 2.005 7.85 2.13 ;
      RECT 7.6 1.995 7.845 2.27 ;
      RECT 7.595 2 7.85 2.13 ;
      RECT 7.63 1.979 7.831 2.27 ;
      RECT 7.716 1.97 7.831 2.27 ;
      RECT 7.716 1.964 7.745 2.27 ;
      RECT 7.205 1.605 7.215 2.095 ;
      RECT 6.865 1.54 6.875 1.84 ;
      RECT 7.38 1.712 7.385 1.931 ;
      RECT 7.37 1.692 7.38 1.948 ;
      RECT 7.36 1.672 7.37 1.978 ;
      RECT 7.355 1.662 7.36 1.993 ;
      RECT 7.35 1.658 7.355 1.998 ;
      RECT 7.335 1.65 7.35 2.005 ;
      RECT 7.295 1.63 7.335 2.03 ;
      RECT 7.27 1.612 7.295 2.063 ;
      RECT 7.265 1.61 7.27 2.076 ;
      RECT 7.245 1.607 7.265 2.08 ;
      RECT 7.215 1.605 7.245 2.09 ;
      RECT 7.145 1.607 7.205 2.091 ;
      RECT 7.125 1.607 7.145 2.085 ;
      RECT 7.1 1.605 7.125 2.082 ;
      RECT 7.065 1.6 7.1 2.078 ;
      RECT 7.045 1.594 7.065 2.065 ;
      RECT 7.035 1.591 7.045 2.053 ;
      RECT 7.015 1.588 7.035 2.038 ;
      RECT 6.995 1.584 7.015 2.02 ;
      RECT 6.99 1.581 6.995 2.01 ;
      RECT 6.985 1.58 6.99 2.008 ;
      RECT 6.975 1.577 6.985 2 ;
      RECT 6.965 1.571 6.975 1.983 ;
      RECT 6.955 1.565 6.965 1.965 ;
      RECT 6.945 1.559 6.955 1.953 ;
      RECT 6.935 1.553 6.945 1.933 ;
      RECT 6.93 1.549 6.935 1.918 ;
      RECT 6.925 1.547 6.93 1.91 ;
      RECT 6.92 1.545 6.925 1.903 ;
      RECT 6.915 1.543 6.92 1.893 ;
      RECT 6.91 1.541 6.915 1.887 ;
      RECT 6.9 1.54 6.91 1.877 ;
      RECT 6.89 1.54 6.9 1.868 ;
      RECT 6.875 1.54 6.89 1.853 ;
      RECT 6.835 1.54 6.865 1.837 ;
      RECT 6.815 1.542 6.835 1.832 ;
      RECT 6.81 1.547 6.815 1.83 ;
      RECT 6.78 1.555 6.81 1.828 ;
      RECT 6.75 1.57 6.78 1.827 ;
      RECT 6.705 1.592 6.75 1.832 ;
      RECT 6.7 1.607 6.705 1.836 ;
      RECT 6.685 1.612 6.7 1.838 ;
      RECT 6.68 1.616 6.685 1.84 ;
      RECT 6.62 1.639 6.68 1.849 ;
      RECT 6.6 1.665 6.62 1.862 ;
      RECT 6.59 1.672 6.6 1.866 ;
      RECT 6.575 1.679 6.59 1.869 ;
      RECT 6.555 1.689 6.575 1.872 ;
      RECT 6.55 1.697 6.555 1.875 ;
      RECT 6.505 1.702 6.55 1.882 ;
      RECT 6.495 1.705 6.505 1.889 ;
      RECT 6.485 1.705 6.495 1.893 ;
      RECT 6.45 1.707 6.485 1.905 ;
      RECT 6.43 1.71 6.45 1.918 ;
      RECT 6.39 1.713 6.43 1.929 ;
      RECT 6.375 1.715 6.39 1.942 ;
      RECT 6.365 1.715 6.375 1.947 ;
      RECT 6.34 1.716 6.365 1.955 ;
      RECT 6.33 1.718 6.34 1.96 ;
      RECT 6.325 1.719 6.33 1.963 ;
      RECT 6.3 1.717 6.325 1.966 ;
      RECT 6.285 1.715 6.3 1.967 ;
      RECT 6.265 1.712 6.285 1.969 ;
      RECT 6.245 1.707 6.265 1.969 ;
      RECT 6.185 1.702 6.245 1.966 ;
      RECT 6.15 1.677 6.185 1.962 ;
      RECT 6.14 1.654 6.15 1.96 ;
      RECT 6.11 1.631 6.14 1.96 ;
      RECT 6.1 1.61 6.11 1.96 ;
      RECT 6.075 1.592 6.1 1.958 ;
      RECT 6.06 1.57 6.075 1.955 ;
      RECT 6.045 1.552 6.06 1.953 ;
      RECT 6.025 1.542 6.045 1.951 ;
      RECT 6.01 1.537 6.025 1.95 ;
      RECT 5.995 1.535 6.01 1.949 ;
      RECT 5.965 1.536 5.995 1.947 ;
      RECT 5.945 1.539 5.965 1.945 ;
      RECT 5.888 1.543 5.945 1.945 ;
      RECT 5.802 1.552 5.888 1.945 ;
      RECT 5.716 1.563 5.802 1.945 ;
      RECT 5.63 1.574 5.716 1.945 ;
      RECT 5.61 1.581 5.63 1.953 ;
      RECT 5.6 1.584 5.61 1.96 ;
      RECT 5.535 1.589 5.6 1.978 ;
      RECT 5.505 1.596 5.535 2.003 ;
      RECT 5.495 1.599 5.505 2.01 ;
      RECT 5.45 1.603 5.495 2.015 ;
      RECT 5.42 1.608 5.45 2.02 ;
      RECT 5.419 1.61 5.42 2.02 ;
      RECT 5.333 1.616 5.419 2.02 ;
      RECT 5.247 1.627 5.333 2.02 ;
      RECT 5.161 1.639 5.247 2.02 ;
      RECT 5.075 1.65 5.161 2.02 ;
      RECT 5.06 1.657 5.075 2.015 ;
      RECT 5.055 1.659 5.06 2.009 ;
      RECT 5.035 1.67 5.055 2.004 ;
      RECT 5.025 1.688 5.035 1.998 ;
      RECT 5.02 1.7 5.025 1.798 ;
      RECT 7.315 0.453 7.335 0.54 ;
      RECT 7.31 0.388 7.315 0.572 ;
      RECT 7.3 0.355 7.31 0.577 ;
      RECT 7.295 0.335 7.3 0.583 ;
      RECT 7.265 0.335 7.295 0.6 ;
      RECT 7.216 0.335 7.265 0.636 ;
      RECT 7.13 0.335 7.216 0.694 ;
      RECT 7.101 0.345 7.13 0.743 ;
      RECT 7.015 0.387 7.101 0.796 ;
      RECT 6.995 0.425 7.015 0.843 ;
      RECT 6.97 0.442 6.995 0.863 ;
      RECT 6.96 0.456 6.97 0.883 ;
      RECT 6.955 0.462 6.96 0.893 ;
      RECT 6.95 0.466 6.955 0.9 ;
      RECT 6.9 0.486 6.95 0.905 ;
      RECT 6.835 0.53 6.9 0.905 ;
      RECT 6.81 0.58 6.835 0.905 ;
      RECT 6.8 0.61 6.81 0.905 ;
      RECT 6.795 0.637 6.8 0.905 ;
      RECT 6.79 0.655 6.795 0.905 ;
      RECT 6.78 0.697 6.79 0.905 ;
      RECT 7.13 1.255 7.3 1.43 ;
      RECT 7.07 1.083 7.13 1.418 ;
      RECT 7.06 1.076 7.07 1.401 ;
      RECT 7.015 1.255 7.3 1.381 ;
      RECT 6.996 1.255 7.3 1.359 ;
      RECT 6.91 1.255 7.3 1.324 ;
      RECT 6.89 1.075 7.06 1.28 ;
      RECT 6.89 1.222 7.295 1.28 ;
      RECT 6.89 1.17 7.27 1.28 ;
      RECT 6.89 1.125 7.235 1.28 ;
      RECT 6.89 1.107 7.2 1.28 ;
      RECT 6.89 1.097 7.195 1.28 ;
      RECT 6.61 2.055 6.8 2.28 ;
      RECT 6.6 2.056 6.805 2.275 ;
      RECT 6.6 2.058 6.815 2.255 ;
      RECT 6.6 2.062 6.82 2.24 ;
      RECT 6.6 2.049 6.77 2.275 ;
      RECT 6.6 2.052 6.795 2.275 ;
      RECT 6.61 2.048 6.77 2.28 ;
      RECT 6.696 2.046 6.77 2.28 ;
      RECT 6.32 1.297 6.49 1.535 ;
      RECT 6.32 1.297 6.576 1.449 ;
      RECT 6.32 1.297 6.58 1.359 ;
      RECT 6.37 1.07 6.59 1.338 ;
      RECT 6.365 1.087 6.595 1.311 ;
      RECT 6.33 1.245 6.595 1.311 ;
      RECT 6.35 1.095 6.49 1.535 ;
      RECT 6.34 1.177 6.6 1.294 ;
      RECT 6.335 1.225 6.6 1.294 ;
      RECT 6.34 1.135 6.595 1.311 ;
      RECT 6.365 1.072 6.59 1.338 ;
      RECT 5.93 1.047 6.1 1.245 ;
      RECT 5.93 1.047 6.145 1.22 ;
      RECT 6 0.99 6.17 1.178 ;
      RECT 5.975 1.005 6.17 1.178 ;
      RECT 5.59 1.051 5.62 1.245 ;
      RECT 5.585 1.023 5.59 1.245 ;
      RECT 5.555 0.997 5.585 1.247 ;
      RECT 5.53 0.955 5.555 1.25 ;
      RECT 5.52 0.927 5.53 1.252 ;
      RECT 5.485 0.907 5.52 1.254 ;
      RECT 5.42 0.892 5.485 1.26 ;
      RECT 5.37 0.89 5.42 1.266 ;
      RECT 5.347 0.892 5.37 1.271 ;
      RECT 5.261 0.903 5.347 1.277 ;
      RECT 5.175 0.921 5.261 1.287 ;
      RECT 5.16 0.932 5.175 1.293 ;
      RECT 5.09 0.955 5.16 1.299 ;
      RECT 5.035 0.987 5.09 1.307 ;
      RECT 4.995 1.01 5.035 1.313 ;
      RECT 4.981 1.023 4.995 1.316 ;
      RECT 4.895 1.045 4.981 1.322 ;
      RECT 4.88 1.07 4.895 1.328 ;
      RECT 4.84 1.085 4.88 1.332 ;
      RECT 4.79 1.1 4.84 1.337 ;
      RECT 4.765 1.107 4.79 1.341 ;
      RECT 4.705 1.102 4.765 1.345 ;
      RECT 4.69 1.093 4.705 1.349 ;
      RECT 4.62 1.083 4.69 1.345 ;
      RECT 4.595 1.075 4.615 1.335 ;
      RECT 4.536 1.075 4.595 1.313 ;
      RECT 4.45 1.075 4.536 1.27 ;
      RECT 4.615 1.075 4.62 1.34 ;
      RECT 5.31 0.306 5.48 0.64 ;
      RECT 5.28 0.306 5.48 0.635 ;
      RECT 5.22 0.273 5.28 0.623 ;
      RECT 5.22 0.329 5.49 0.618 ;
      RECT 5.195 0.329 5.49 0.612 ;
      RECT 5.19 0.27 5.22 0.609 ;
      RECT 5.175 0.276 5.31 0.607 ;
      RECT 5.17 0.284 5.395 0.595 ;
      RECT 5.17 0.336 5.505 0.548 ;
      RECT 5.155 0.292 5.395 0.543 ;
      RECT 5.155 0.362 5.515 0.484 ;
      RECT 5.125 0.312 5.48 0.445 ;
      RECT 5.125 0.402 5.525 0.441 ;
      RECT 5.175 0.281 5.395 0.607 ;
      RECT 4.515 0.611 4.57 0.875 ;
      RECT 4.515 0.611 4.635 0.874 ;
      RECT 4.515 0.611 4.66 0.873 ;
      RECT 4.515 0.611 4.725 0.872 ;
      RECT 4.66 0.577 4.74 0.871 ;
      RECT 4.475 0.621 4.885 0.87 ;
      RECT 4.515 0.618 4.885 0.87 ;
      RECT 4.475 0.626 4.89 0.863 ;
      RECT 4.46 0.628 4.89 0.862 ;
      RECT 4.46 0.635 4.895 0.858 ;
      RECT 4.44 0.634 4.89 0.854 ;
      RECT 4.44 0.642 4.9 0.853 ;
      RECT 4.435 0.639 4.895 0.849 ;
      RECT 4.435 0.652 4.91 0.848 ;
      RECT 4.42 0.642 4.9 0.847 ;
      RECT 4.385 0.655 4.91 0.84 ;
      RECT 4.57 0.61 4.88 0.87 ;
      RECT 4.57 0.595 4.83 0.87 ;
      RECT 4.635 0.582 4.765 0.87 ;
      RECT 4.18 1.671 4.195 2.064 ;
      RECT 4.145 1.676 4.195 2.063 ;
      RECT 4.18 1.675 4.24 2.062 ;
      RECT 4.125 1.686 4.24 2.061 ;
      RECT 4.14 1.682 4.24 2.061 ;
      RECT 4.105 1.692 4.315 2.058 ;
      RECT 4.105 1.711 4.36 2.056 ;
      RECT 4.105 1.718 4.365 2.053 ;
      RECT 4.09 1.695 4.315 2.05 ;
      RECT 4.07 1.7 4.315 2.043 ;
      RECT 4.065 1.704 4.315 2.039 ;
      RECT 4.065 1.721 4.375 2.038 ;
      RECT 4.045 1.715 4.36 2.034 ;
      RECT 4.045 1.724 4.38 2.028 ;
      RECT 4.04 1.73 4.38 1.8 ;
      RECT 4.105 1.69 4.24 2.058 ;
      RECT 3.98 1.053 4.18 1.365 ;
      RECT 4.055 1.031 4.18 1.365 ;
      RECT 3.995 1.05 4.185 1.35 ;
      RECT 3.965 1.061 4.185 1.348 ;
      RECT 3.98 1.056 4.19 1.314 ;
      RECT 3.965 1.16 4.195 1.281 ;
      RECT 3.995 1.032 4.18 1.365 ;
      RECT 4.055 1.01 4.155 1.365 ;
      RECT 4.08 1.007 4.155 1.365 ;
      RECT 4.08 1.002 4.1 1.365 ;
      RECT 3.485 1.07 3.66 1.245 ;
      RECT 3.48 1.07 3.66 1.243 ;
      RECT 3.455 1.07 3.66 1.238 ;
      RECT 3.4 1.05 3.57 1.228 ;
      RECT 3.4 1.057 3.635 1.228 ;
      RECT 3.485 1.737 3.5 1.92 ;
      RECT 3.475 1.715 3.485 1.92 ;
      RECT 3.46 1.695 3.475 1.92 ;
      RECT 3.45 1.67 3.46 1.92 ;
      RECT 3.42 1.635 3.45 1.92 ;
      RECT 3.385 1.575 3.42 1.92 ;
      RECT 3.38 1.537 3.385 1.92 ;
      RECT 3.33 1.488 3.38 1.92 ;
      RECT 3.32 1.438 3.33 1.908 ;
      RECT 3.305 1.417 3.32 1.868 ;
      RECT 3.285 1.385 3.305 1.818 ;
      RECT 3.26 1.341 3.285 1.758 ;
      RECT 3.255 1.313 3.26 1.713 ;
      RECT 3.25 1.304 3.255 1.699 ;
      RECT 3.245 1.297 3.25 1.686 ;
      RECT 3.24 1.292 3.245 1.675 ;
      RECT 3.235 1.277 3.24 1.665 ;
      RECT 3.23 1.255 3.235 1.652 ;
      RECT 3.22 1.215 3.23 1.627 ;
      RECT 3.195 1.145 3.22 1.583 ;
      RECT 3.19 1.085 3.195 1.548 ;
      RECT 3.175 1.065 3.19 1.515 ;
      RECT 3.17 1.065 3.175 1.49 ;
      RECT 3.14 1.065 3.17 1.445 ;
      RECT 3.095 1.065 3.14 1.385 ;
      RECT 3.02 1.065 3.095 1.333 ;
      RECT 3.015 1.065 3.02 1.298 ;
      RECT 3.01 1.065 3.015 1.288 ;
      RECT 3.005 1.065 3.01 1.268 ;
      RECT 3.27 0.285 3.44 0.755 ;
      RECT 3.215 0.278 3.41 0.739 ;
      RECT 3.215 0.292 3.445 0.738 ;
      RECT 3.2 0.293 3.445 0.719 ;
      RECT 3.195 0.311 3.445 0.705 ;
      RECT 3.2 0.294 3.45 0.703 ;
      RECT 3.185 0.325 3.45 0.688 ;
      RECT 3.2 0.3 3.455 0.673 ;
      RECT 3.18 0.34 3.455 0.67 ;
      RECT 3.195 0.312 3.46 0.655 ;
      RECT 3.195 0.324 3.465 0.635 ;
      RECT 3.18 0.34 3.47 0.618 ;
      RECT 3.18 0.35 3.475 0.473 ;
      RECT 3.175 0.35 3.475 0.43 ;
      RECT 3.175 0.365 3.48 0.408 ;
      RECT 3.27 0.275 3.41 0.755 ;
      RECT 3.27 0.273 3.38 0.755 ;
      RECT 3.356 0.27 3.38 0.755 ;
      RECT 3.015 1.937 3.02 1.983 ;
      RECT 3.005 1.785 3.015 2.007 ;
      RECT 3 1.63 3.005 2.032 ;
      RECT 2.985 1.592 3 2.043 ;
      RECT 2.98 1.575 2.985 2.05 ;
      RECT 2.97 1.563 2.98 2.057 ;
      RECT 2.965 1.554 2.97 2.059 ;
      RECT 2.96 1.552 2.965 2.063 ;
      RECT 2.915 1.543 2.96 2.078 ;
      RECT 2.91 1.535 2.915 2.092 ;
      RECT 2.905 1.532 2.91 2.096 ;
      RECT 2.89 1.527 2.905 2.104 ;
      RECT 2.835 1.517 2.89 2.115 ;
      RECT 2.8 1.505 2.835 2.116 ;
      RECT 2.791 1.5 2.8 2.11 ;
      RECT 2.705 1.5 2.791 2.1 ;
      RECT 2.675 1.5 2.705 2.078 ;
      RECT 2.665 1.5 2.67 2.058 ;
      RECT 2.66 1.5 2.665 2.02 ;
      RECT 2.655 1.5 2.66 1.978 ;
      RECT 2.65 1.5 2.655 1.938 ;
      RECT 2.645 1.5 2.65 1.868 ;
      RECT 2.635 1.5 2.645 1.79 ;
      RECT 2.63 1.5 2.635 1.69 ;
      RECT 2.67 1.5 2.675 2.06 ;
      RECT 2.165 1.582 2.255 2.06 ;
      RECT 2.15 1.585 2.27 2.058 ;
      RECT 2.165 1.584 2.27 2.058 ;
      RECT 2.13 1.591 2.295 2.048 ;
      RECT 2.15 1.585 2.295 2.048 ;
      RECT 2.115 1.597 2.295 2.036 ;
      RECT 2.15 1.588 2.345 2.029 ;
      RECT 2.101 1.605 2.345 2.027 ;
      RECT 2.13 1.595 2.355 2.015 ;
      RECT 2.101 1.616 2.385 2.006 ;
      RECT 2.015 1.64 2.385 2 ;
      RECT 2.015 1.653 2.425 1.983 ;
      RECT 2.01 1.675 2.425 1.976 ;
      RECT 1.98 1.69 2.425 1.966 ;
      RECT 1.975 1.701 2.425 1.956 ;
      RECT 1.945 1.714 2.425 1.947 ;
      RECT 1.93 1.732 2.425 1.936 ;
      RECT 1.905 1.745 2.425 1.926 ;
      RECT 2.165 1.581 2.175 2.06 ;
      RECT 2.211 1.005 2.25 1.25 ;
      RECT 2.125 1.005 2.26 1.248 ;
      RECT 2.01 1.03 2.26 1.245 ;
      RECT 2.01 1.03 2.265 1.243 ;
      RECT 2.01 1.03 2.28 1.238 ;
      RECT 2.116 1.005 2.295 1.218 ;
      RECT 2.03 1.013 2.295 1.218 ;
      RECT 1.7 0.365 1.87 0.8 ;
      RECT 1.69 0.399 1.87 0.783 ;
      RECT 1.77 0.335 1.94 0.77 ;
      RECT 1.675 0.41 1.94 0.748 ;
      RECT 1.77 0.345 1.945 0.738 ;
      RECT 1.7 0.397 1.975 0.723 ;
      RECT 1.66 0.423 1.975 0.708 ;
      RECT 1.66 0.465 1.985 0.688 ;
      RECT 1.655 0.49 1.99 0.67 ;
      RECT 1.655 0.5 1.995 0.655 ;
      RECT 1.65 0.437 1.975 0.653 ;
      RECT 1.65 0.51 2 0.638 ;
      RECT 1.645 0.447 1.975 0.635 ;
      RECT 1.64 0.531 2.005 0.618 ;
      RECT 1.64 0.563 2.01 0.598 ;
      RECT 1.635 0.477 1.985 0.59 ;
      RECT 1.64 0.462 1.975 0.618 ;
      RECT 1.655 0.432 1.975 0.67 ;
      RECT 1.5 1.019 1.725 1.275 ;
      RECT 1.5 1.052 1.745 1.265 ;
      RECT 1.465 1.052 1.745 1.263 ;
      RECT 1.465 1.065 1.75 1.253 ;
      RECT 1.465 1.085 1.76 1.245 ;
      RECT 1.465 1.182 1.765 1.238 ;
      RECT 1.445 0.93 1.575 1.228 ;
      RECT 1.4 1.085 1.76 1.17 ;
      RECT 1.39 0.93 1.575 1.115 ;
      RECT 1.39 0.962 1.661 1.115 ;
      RECT 1.355 1.492 1.375 1.67 ;
      RECT 1.32 1.445 1.355 1.67 ;
      RECT 1.305 1.385 1.32 1.67 ;
      RECT 1.28 1.332 1.305 1.67 ;
      RECT 1.265 1.285 1.28 1.67 ;
      RECT 1.245 1.262 1.265 1.67 ;
      RECT 1.22 1.227 1.245 1.67 ;
      RECT 1.21 1.073 1.22 1.67 ;
      RECT 1.18 1.068 1.21 1.661 ;
      RECT 1.175 1.065 1.18 1.651 ;
      RECT 1.16 1.065 1.175 1.625 ;
      RECT 1.155 1.065 1.16 1.588 ;
      RECT 1.13 1.065 1.155 1.54 ;
      RECT 1.11 1.065 1.13 1.465 ;
      RECT 1.1 1.065 1.11 1.425 ;
      RECT 1.095 1.065 1.1 1.4 ;
      RECT 1.09 1.065 1.095 1.383 ;
      RECT 1.085 1.065 1.09 1.365 ;
      RECT 1.08 1.066 1.085 1.355 ;
      RECT 1.07 1.068 1.08 1.323 ;
      RECT 1.06 1.07 1.07 1.29 ;
      RECT 1.05 1.073 1.06 1.263 ;
      RECT 1.375 1.5 1.6 1.67 ;
      RECT 0.705 0.312 0.875 0.765 ;
      RECT 0.705 0.312 0.965 0.731 ;
      RECT 0.705 0.312 0.995 0.715 ;
      RECT 0.705 0.312 1.025 0.688 ;
      RECT 0.961 0.29 1.04 0.67 ;
      RECT 0.74 0.297 1.045 0.655 ;
      RECT 0.74 0.305 1.055 0.618 ;
      RECT 0.7 0.332 1.055 0.59 ;
      RECT 0.685 0.345 1.055 0.555 ;
      RECT 0.705 0.32 1.075 0.545 ;
      RECT 0.68 0.385 1.075 0.515 ;
      RECT 0.68 0.415 1.08 0.498 ;
      RECT 0.675 0.445 1.08 0.485 ;
      RECT 0.74 0.294 1.04 0.67 ;
      RECT 0.875 0.291 0.961 0.749 ;
      RECT 0.826 0.292 1.04 0.67 ;
      RECT 0.97 1.952 1.015 2.145 ;
      RECT 0.96 1.922 0.97 2.145 ;
      RECT 0.955 1.907 0.96 2.145 ;
      RECT 0.915 1.817 0.955 2.145 ;
      RECT 0.91 1.73 0.915 2.145 ;
      RECT 0.9 1.7 0.91 2.145 ;
      RECT 0.895 1.66 0.9 2.145 ;
      RECT 0.885 1.622 0.895 2.145 ;
      RECT 0.88 1.587 0.885 2.145 ;
      RECT 0.86 1.54 0.88 2.145 ;
      RECT 0.845 1.465 0.86 2.145 ;
      RECT 0.84 1.42 0.845 2.14 ;
      RECT 0.835 1.4 0.84 2.113 ;
      RECT 0.83 1.38 0.835 2.098 ;
      RECT 0.825 1.355 0.83 2.078 ;
      RECT 0.82 1.333 0.825 2.063 ;
      RECT 0.815 1.311 0.82 2.045 ;
      RECT 0.81 1.29 0.815 2.035 ;
      RECT 0.8 1.262 0.81 2.005 ;
      RECT 0.79 1.225 0.8 1.973 ;
      RECT 0.78 1.185 0.79 1.94 ;
      RECT 0.77 1.163 0.78 1.91 ;
      RECT 0.74 1.115 0.77 1.842 ;
      RECT 0.725 1.075 0.74 1.769 ;
      RECT 0.715 1.075 0.725 1.735 ;
      RECT 0.71 1.075 0.715 1.71 ;
      RECT 0.705 1.075 0.71 1.695 ;
      RECT 0.7 1.075 0.705 1.673 ;
      RECT 0.695 1.075 0.7 1.66 ;
      RECT 0.68 1.075 0.695 1.625 ;
      RECT 0.66 1.075 0.68 1.565 ;
      RECT 0.65 1.075 0.66 1.515 ;
      RECT 0.63 1.075 0.65 1.463 ;
      RECT 0.61 1.075 0.63 1.42 ;
      RECT 0.6 1.075 0.61 1.408 ;
      RECT 0.57 1.075 0.6 1.395 ;
      RECT 0.54 1.096 0.57 1.375 ;
      RECT 0.53 1.124 0.54 1.355 ;
      RECT 0.515 1.141 0.53 1.323 ;
      RECT 0.51 1.155 0.515 1.29 ;
      RECT 0.505 1.163 0.51 1.263 ;
      RECT 0.5 1.171 0.505 1.225 ;
      RECT 0.505 1.695 0.51 2.03 ;
      RECT 0.47 1.682 0.505 2.029 ;
      RECT 0.4 1.622 0.47 2.028 ;
      RECT 0.32 1.565 0.4 2.027 ;
      RECT 0.185 1.525 0.32 2.026 ;
      RECT 0.185 1.712 0.52 2.015 ;
      RECT 0.145 1.712 0.52 2.005 ;
      RECT 0.145 1.73 0.525 2 ;
      RECT 0.145 1.82 0.53 1.99 ;
      RECT 0.14 1.515 0.305 1.97 ;
      RECT 0.135 1.515 0.305 1.713 ;
      RECT 0.135 1.672 0.5 1.713 ;
      RECT 0.135 1.66 0.495 1.713 ;
  END
END scs130hd_mpr2aa_8

MACRO scs130hd_mpr2at_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130hd_mpr2at_8 0 0 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT 9.305 2.04 9.86 2.37 ;
      RECT 9.305 0.375 9.605 2.37 ;
      RECT 5.37 1.48 5.925 1.81 ;
      RECT 5.625 0.375 5.925 1.81 ;
      RECT 6.42 0.24 6.57 0.89 ;
      RECT 5.625 0.375 9.605 0.675 ;
      RECT 10.49 0.36 11.22 0.69 ;
      RECT 8.27 2.04 9 2.37 ;
      RECT 6.57 2.04 7.3 2.37 ;
      RECT 4.13 0.92 4.86 1.25 ;
      RECT 2.69 1.48 3.42 1.81 ;
      RECT 1.615 0.92 2.345 1.25 ;
      RECT 0.58 0.92 1.31 1.25 ;
      RECT 0.25 2.04 0.98 2.37 ;
    LAYER via2 ;
      RECT 10.555 0.425 10.755 0.625 ;
      RECT 9.595 2.105 9.795 2.305 ;
      RECT 8.595 2.105 8.795 2.305 ;
      RECT 6.635 2.105 6.835 2.305 ;
      RECT 5.435 1.545 5.635 1.745 ;
      RECT 4.195 0.985 4.395 1.185 ;
      RECT 2.755 1.545 2.955 1.745 ;
      RECT 2.015 0.985 2.215 1.185 ;
      RECT 0.795 0.985 0.995 1.185 ;
      RECT 0.315 2.105 0.515 2.305 ;
    LAYER met2 ;
      RECT 10.55 0.515 10.81 0.775 ;
      RECT 10.545 0.515 10.81 0.723 ;
      RECT 10.54 0.515 10.81 0.693 ;
      RECT 10.515 0.385 10.795 0.665 ;
      RECT 9.555 2.065 9.835 2.345 ;
      RECT 9.595 2.02 9.86 2.28 ;
      RECT 9.585 2.055 9.86 2.28 ;
      RECT 9.59 2.04 9.835 2.345 ;
      RECT 9.595 2.017 9.805 2.345 ;
      RECT 9.595 2.015 9.79 2.345 ;
      RECT 9.635 2.005 9.79 2.345 ;
      RECT 9.605 2.01 9.79 2.345 ;
      RECT 9.635 2.002 9.735 2.345 ;
      RECT 9.66 1.995 9.735 2.345 ;
      RECT 9.64 1.997 9.735 2.345 ;
      RECT 8.97 1.51 9.23 1.77 ;
      RECT 9.02 1.502 9.21 1.77 ;
      RECT 9.025 1.422 9.21 1.77 ;
      RECT 9.145 0.81 9.21 1.77 ;
      RECT 9.05 1.207 9.21 1.77 ;
      RECT 9.125 0.895 9.21 1.77 ;
      RECT 9.16 0.52 9.296 1.248 ;
      RECT 9.105 1.017 9.296 1.248 ;
      RECT 9.12 0.957 9.21 1.77 ;
      RECT 9.16 0.52 9.32 0.913 ;
      RECT 9.16 0.52 9.33 0.81 ;
      RECT 9.15 0.52 9.41 0.78 ;
      RECT 8.555 2.065 8.835 2.345 ;
      RECT 8.575 2.025 8.835 2.345 ;
      RECT 8.215 1.98 8.32 2.24 ;
      RECT 8.07 0.47 8.16 0.73 ;
      RECT 8.61 1.535 8.615 1.575 ;
      RECT 8.605 1.525 8.61 1.66 ;
      RECT 8.6 1.515 8.605 1.753 ;
      RECT 8.59 1.495 8.6 1.809 ;
      RECT 8.51 1.423 8.59 1.889 ;
      RECT 8.545 2.067 8.555 2.292 ;
      RECT 8.54 2.064 8.545 2.287 ;
      RECT 8.525 2.061 8.54 2.28 ;
      RECT 8.49 2.055 8.525 2.262 ;
      RECT 8.505 1.358 8.51 1.963 ;
      RECT 8.485 1.309 8.505 1.978 ;
      RECT 8.475 2.042 8.49 2.245 ;
      RECT 8.48 1.251 8.485 1.993 ;
      RECT 8.475 1.229 8.48 2.003 ;
      RECT 8.44 1.139 8.475 2.24 ;
      RECT 8.425 1.017 8.44 2.24 ;
      RECT 8.42 0.97 8.425 2.24 ;
      RECT 8.395 0.895 8.42 2.24 ;
      RECT 8.38 0.81 8.395 2.24 ;
      RECT 8.375 0.757 8.38 2.24 ;
      RECT 8.37 0.737 8.375 2.24 ;
      RECT 8.365 0.712 8.37 1.474 ;
      RECT 8.35 1.672 8.37 2.24 ;
      RECT 8.36 0.69 8.365 1.451 ;
      RECT 8.35 0.642 8.36 1.416 ;
      RECT 8.345 0.605 8.35 1.382 ;
      RECT 8.345 1.752 8.35 2.24 ;
      RECT 8.33 0.582 8.345 1.337 ;
      RECT 8.325 1.85 8.345 2.24 ;
      RECT 8.275 0.47 8.33 1.179 ;
      RECT 8.32 1.972 8.325 2.24 ;
      RECT 8.26 0.47 8.275 1.018 ;
      RECT 8.255 0.47 8.26 0.97 ;
      RECT 8.25 0.47 8.255 0.958 ;
      RECT 8.205 0.47 8.25 0.895 ;
      RECT 8.18 0.47 8.205 0.813 ;
      RECT 8.165 0.47 8.18 0.765 ;
      RECT 8.16 0.47 8.165 0.735 ;
      RECT 7.485 1.92 7.53 2.18 ;
      RECT 7.39 0.455 7.535 0.715 ;
      RECT 7.895 1.077 7.905 1.168 ;
      RECT 7.88 1.015 7.895 1.224 ;
      RECT 7.875 0.962 7.88 1.27 ;
      RECT 7.825 0.909 7.875 1.396 ;
      RECT 7.82 0.864 7.825 1.543 ;
      RECT 7.81 0.852 7.82 1.585 ;
      RECT 7.775 0.816 7.81 1.69 ;
      RECT 7.77 0.784 7.775 1.796 ;
      RECT 7.755 0.766 7.77 1.841 ;
      RECT 7.75 0.749 7.755 1.075 ;
      RECT 7.745 1.13 7.755 1.898 ;
      RECT 7.74 0.735 7.75 1.048 ;
      RECT 7.735 1.185 7.745 2.18 ;
      RECT 7.73 0.721 7.74 1.033 ;
      RECT 7.73 1.235 7.735 2.18 ;
      RECT 7.715 0.698 7.73 1.013 ;
      RECT 7.695 1.357 7.73 2.18 ;
      RECT 7.71 0.68 7.715 0.995 ;
      RECT 7.705 0.672 7.71 0.985 ;
      RECT 7.675 0.64 7.705 0.949 ;
      RECT 7.685 1.485 7.695 2.18 ;
      RECT 7.68 1.512 7.685 2.18 ;
      RECT 7.675 1.562 7.68 2.18 ;
      RECT 7.665 0.606 7.675 0.914 ;
      RECT 7.625 1.63 7.675 2.18 ;
      RECT 7.65 0.583 7.665 0.89 ;
      RECT 7.625 0.455 7.65 0.853 ;
      RECT 7.62 0.455 7.625 0.825 ;
      RECT 7.59 1.73 7.625 2.18 ;
      RECT 7.615 0.455 7.62 0.818 ;
      RECT 7.61 0.455 7.615 0.808 ;
      RECT 7.595 0.455 7.61 0.793 ;
      RECT 7.58 0.455 7.595 0.765 ;
      RECT 7.545 1.835 7.59 2.18 ;
      RECT 7.565 0.455 7.58 0.738 ;
      RECT 7.535 0.455 7.565 0.723 ;
      RECT 7.53 1.907 7.545 2.18 ;
      RECT 7.455 0.99 7.495 1.25 ;
      RECT 7.23 0.937 7.235 1.195 ;
      RECT 3.185 0.415 3.445 0.675 ;
      RECT 3.185 0.44 3.46 0.655 ;
      RECT 5.575 0.265 5.58 0.41 ;
      RECT 7.445 0.985 7.455 1.25 ;
      RECT 7.425 0.977 7.445 1.25 ;
      RECT 7.407 0.973 7.425 1.25 ;
      RECT 7.321 0.962 7.407 1.25 ;
      RECT 7.235 0.945 7.321 1.25 ;
      RECT 7.18 0.932 7.23 1.18 ;
      RECT 7.146 0.924 7.18 1.155 ;
      RECT 7.06 0.913 7.146 1.12 ;
      RECT 7.025 0.89 7.06 1.085 ;
      RECT 7.015 0.852 7.025 1.071 ;
      RECT 7.01 0.825 7.015 1.067 ;
      RECT 7.005 0.812 7.01 1.064 ;
      RECT 6.995 0.792 7.005 1.06 ;
      RECT 6.99 0.767 6.995 1.056 ;
      RECT 6.965 0.722 6.99 1.05 ;
      RECT 6.955 0.663 6.965 1.042 ;
      RECT 6.945 0.631 6.955 1.033 ;
      RECT 6.925 0.583 6.945 1.013 ;
      RECT 6.92 0.543 6.925 0.983 ;
      RECT 6.905 0.517 6.92 0.957 ;
      RECT 6.9 0.495 6.905 0.933 ;
      RECT 6.885 0.467 6.9 0.909 ;
      RECT 6.87 0.44 6.885 0.873 ;
      RECT 6.855 0.417 6.87 0.835 ;
      RECT 6.85 0.407 6.855 0.81 ;
      RECT 6.84 0.4 6.85 0.793 ;
      RECT 6.825 0.387 6.84 0.763 ;
      RECT 6.82 0.377 6.825 0.738 ;
      RECT 6.815 0.372 6.82 0.725 ;
      RECT 6.805 0.365 6.815 0.705 ;
      RECT 6.8 0.358 6.805 0.69 ;
      RECT 6.775 0.351 6.8 0.648 ;
      RECT 6.76 0.341 6.775 0.598 ;
      RECT 6.75 0.336 6.76 0.568 ;
      RECT 6.74 0.332 6.75 0.543 ;
      RECT 6.725 0.329 6.74 0.533 ;
      RECT 6.675 0.326 6.725 0.518 ;
      RECT 6.655 0.324 6.675 0.503 ;
      RECT 6.606 0.322 6.655 0.498 ;
      RECT 6.52 0.318 6.606 0.493 ;
      RECT 6.481 0.315 6.52 0.489 ;
      RECT 6.395 0.311 6.481 0.484 ;
      RECT 6.345 0.308 6.395 0.478 ;
      RECT 6.296 0.305 6.345 0.473 ;
      RECT 6.21 0.302 6.296 0.468 ;
      RECT 6.206 0.3 6.21 0.465 ;
      RECT 6.12 0.297 6.206 0.46 ;
      RECT 6.071 0.293 6.12 0.453 ;
      RECT 5.985 0.29 6.071 0.448 ;
      RECT 5.961 0.287 5.985 0.444 ;
      RECT 5.875 0.285 5.961 0.439 ;
      RECT 5.81 0.281 5.875 0.432 ;
      RECT 5.807 0.28 5.81 0.429 ;
      RECT 5.721 0.277 5.807 0.426 ;
      RECT 5.635 0.271 5.721 0.419 ;
      RECT 5.605 0.267 5.635 0.415 ;
      RECT 5.58 0.265 5.605 0.413 ;
      RECT 5.525 0.262 5.575 0.41 ;
      RECT 5.445 0.261 5.525 0.41 ;
      RECT 5.39 0.263 5.445 0.413 ;
      RECT 5.375 0.264 5.39 0.417 ;
      RECT 5.32 0.272 5.375 0.427 ;
      RECT 5.29 0.28 5.32 0.44 ;
      RECT 5.271 0.281 5.29 0.446 ;
      RECT 5.185 0.284 5.271 0.451 ;
      RECT 5.115 0.289 5.185 0.46 ;
      RECT 5.096 0.292 5.115 0.466 ;
      RECT 5.01 0.296 5.096 0.471 ;
      RECT 4.97 0.3 5.01 0.478 ;
      RECT 4.961 0.302 4.97 0.481 ;
      RECT 4.875 0.306 4.961 0.486 ;
      RECT 4.872 0.309 4.875 0.49 ;
      RECT 4.786 0.312 4.872 0.494 ;
      RECT 4.7 0.318 4.786 0.502 ;
      RECT 4.676 0.322 4.7 0.506 ;
      RECT 4.59 0.326 4.676 0.511 ;
      RECT 4.545 0.331 4.59 0.518 ;
      RECT 4.465 0.336 4.545 0.525 ;
      RECT 4.385 0.342 4.465 0.54 ;
      RECT 4.36 0.346 4.385 0.553 ;
      RECT 4.295 0.349 4.36 0.565 ;
      RECT 4.24 0.354 4.295 0.58 ;
      RECT 4.21 0.357 4.24 0.598 ;
      RECT 4.2 0.359 4.21 0.611 ;
      RECT 4.14 0.374 4.2 0.621 ;
      RECT 4.125 0.391 4.14 0.63 ;
      RECT 4.12 0.4 4.125 0.63 ;
      RECT 4.11 0.41 4.12 0.63 ;
      RECT 4.1 0.427 4.11 0.63 ;
      RECT 4.08 0.437 4.1 0.631 ;
      RECT 4.035 0.447 4.08 0.632 ;
      RECT 4 0.456 4.035 0.634 ;
      RECT 3.935 0.461 4 0.636 ;
      RECT 3.855 0.462 3.935 0.639 ;
      RECT 3.851 0.46 3.855 0.64 ;
      RECT 3.765 0.457 3.851 0.642 ;
      RECT 3.718 0.454 3.765 0.644 ;
      RECT 3.632 0.45 3.718 0.647 ;
      RECT 3.546 0.446 3.632 0.65 ;
      RECT 3.46 0.442 3.546 0.654 ;
      RECT 6.845 2.065 6.875 2.345 ;
      RECT 6.595 1.955 6.615 2.345 ;
      RECT 6.55 1.955 6.615 2.215 ;
      RECT 6.38 0.58 6.415 0.84 ;
      RECT 6.155 0.58 6.215 0.84 ;
      RECT 6.835 2.045 6.845 2.345 ;
      RECT 6.83 2.005 6.835 2.345 ;
      RECT 6.815 1.96 6.83 2.345 ;
      RECT 6.81 1.925 6.815 2.345 ;
      RECT 6.805 1.905 6.81 2.345 ;
      RECT 6.775 1.832 6.805 2.345 ;
      RECT 6.755 1.73 6.775 2.345 ;
      RECT 6.745 1.66 6.755 2.345 ;
      RECT 6.7 1.6 6.745 2.345 ;
      RECT 6.615 1.561 6.7 2.345 ;
      RECT 6.61 1.552 6.615 1.925 ;
      RECT 6.6 1.551 6.61 1.908 ;
      RECT 6.575 1.532 6.6 1.878 ;
      RECT 6.57 1.507 6.575 1.857 ;
      RECT 6.56 1.485 6.57 1.848 ;
      RECT 6.555 1.456 6.56 1.838 ;
      RECT 6.515 1.382 6.555 1.81 ;
      RECT 6.495 1.283 6.515 1.775 ;
      RECT 6.48 1.219 6.495 1.758 ;
      RECT 6.45 1.143 6.48 1.73 ;
      RECT 6.43 1.058 6.45 1.703 ;
      RECT 6.39 0.954 6.43 1.61 ;
      RECT 6.385 0.875 6.39 1.518 ;
      RECT 6.38 0.858 6.385 1.495 ;
      RECT 6.375 0.58 6.38 1.475 ;
      RECT 6.345 0.58 6.375 1.413 ;
      RECT 6.34 0.58 6.345 1.345 ;
      RECT 6.33 0.58 6.34 1.31 ;
      RECT 6.32 0.58 6.33 1.275 ;
      RECT 6.255 0.58 6.32 1.13 ;
      RECT 6.25 0.58 6.255 1 ;
      RECT 6.22 0.58 6.25 0.933 ;
      RECT 6.215 0.58 6.22 0.858 ;
      RECT 5.395 1.505 5.675 1.785 ;
      RECT 5.435 1.485 5.695 1.745 ;
      RECT 5.425 1.495 5.695 1.745 ;
      RECT 5.435 1.422 5.65 1.785 ;
      RECT 5.49 1.345 5.645 1.785 ;
      RECT 5.495 1.13 5.645 1.785 ;
      RECT 5.485 0.932 5.635 1.183 ;
      RECT 5.475 0.932 5.635 1.05 ;
      RECT 5.47 0.81 5.63 0.953 ;
      RECT 5.455 0.81 5.63 0.858 ;
      RECT 5.45 0.52 5.625 0.835 ;
      RECT 5.435 0.52 5.625 0.805 ;
      RECT 5.395 0.52 5.655 0.78 ;
      RECT 5.305 1.99 5.385 2.25 ;
      RECT 4.71 0.71 4.715 0.975 ;
      RECT 4.59 0.71 4.715 0.97 ;
      RECT 5.265 1.955 5.305 2.25 ;
      RECT 5.22 1.877 5.265 2.25 ;
      RECT 5.2 1.805 5.22 2.25 ;
      RECT 5.19 1.757 5.2 2.25 ;
      RECT 5.155 1.69 5.19 2.25 ;
      RECT 5.125 1.59 5.155 2.25 ;
      RECT 5.105 1.515 5.125 2.05 ;
      RECT 5.095 1.465 5.105 2.005 ;
      RECT 5.09 1.442 5.095 1.978 ;
      RECT 5.085 1.427 5.09 1.965 ;
      RECT 5.08 1.412 5.085 1.943 ;
      RECT 5.075 1.397 5.08 1.925 ;
      RECT 5.05 1.352 5.075 1.88 ;
      RECT 5.04 1.3 5.05 1.823 ;
      RECT 5.03 1.27 5.04 1.79 ;
      RECT 5.02 1.235 5.03 1.758 ;
      RECT 4.985 1.167 5.02 1.69 ;
      RECT 4.98 1.106 4.985 1.625 ;
      RECT 4.97 1.094 4.98 1.605 ;
      RECT 4.965 1.082 4.97 1.585 ;
      RECT 4.96 1.074 4.965 1.573 ;
      RECT 4.955 1.066 4.96 1.553 ;
      RECT 4.945 1.054 4.955 1.525 ;
      RECT 4.935 1.038 4.945 1.495 ;
      RECT 4.91 1.01 4.935 1.433 ;
      RECT 4.9 0.981 4.91 1.378 ;
      RECT 4.885 0.96 4.9 1.338 ;
      RECT 4.88 0.944 4.885 1.31 ;
      RECT 4.875 0.932 4.88 1.3 ;
      RECT 4.87 0.927 4.875 1.273 ;
      RECT 4.865 0.92 4.87 1.26 ;
      RECT 4.85 0.903 4.865 1.233 ;
      RECT 4.84 0.71 4.85 1.193 ;
      RECT 4.83 0.71 4.84 1.16 ;
      RECT 4.82 0.71 4.83 1.135 ;
      RECT 4.75 0.71 4.82 1.07 ;
      RECT 4.74 0.71 4.75 1.018 ;
      RECT 4.725 0.71 4.74 1 ;
      RECT 4.715 0.71 4.725 0.985 ;
      RECT 4.545 1.58 4.805 1.84 ;
      RECT 3.08 1.615 3.085 1.822 ;
      RECT 2.715 1.505 2.79 1.82 ;
      RECT 2.53 1.56 2.685 1.82 ;
      RECT 2.715 1.505 2.82 1.785 ;
      RECT 4.53 1.677 4.545 1.838 ;
      RECT 4.505 1.685 4.53 1.843 ;
      RECT 4.48 1.692 4.505 1.848 ;
      RECT 4.417 1.703 4.48 1.857 ;
      RECT 4.331 1.722 4.417 1.874 ;
      RECT 4.245 1.744 4.331 1.893 ;
      RECT 4.23 1.757 4.245 1.904 ;
      RECT 4.19 1.765 4.23 1.911 ;
      RECT 4.17 1.77 4.19 1.918 ;
      RECT 4.132 1.771 4.17 1.921 ;
      RECT 4.046 1.774 4.132 1.922 ;
      RECT 3.96 1.778 4.046 1.923 ;
      RECT 3.911 1.78 3.96 1.925 ;
      RECT 3.825 1.78 3.911 1.927 ;
      RECT 3.785 1.775 3.825 1.929 ;
      RECT 3.775 1.769 3.785 1.93 ;
      RECT 3.735 1.764 3.775 1.927 ;
      RECT 3.725 1.757 3.735 1.923 ;
      RECT 3.71 1.753 3.725 1.921 ;
      RECT 3.693 1.749 3.71 1.919 ;
      RECT 3.607 1.739 3.693 1.911 ;
      RECT 3.521 1.721 3.607 1.897 ;
      RECT 3.435 1.704 3.521 1.883 ;
      RECT 3.41 1.692 3.435 1.874 ;
      RECT 3.34 1.682 3.41 1.867 ;
      RECT 3.295 1.67 3.34 1.858 ;
      RECT 3.235 1.657 3.295 1.85 ;
      RECT 3.23 1.649 3.235 1.845 ;
      RECT 3.195 1.644 3.23 1.843 ;
      RECT 3.14 1.635 3.195 1.836 ;
      RECT 3.1 1.624 3.14 1.828 ;
      RECT 3.085 1.617 3.1 1.824 ;
      RECT 3.065 1.61 3.08 1.821 ;
      RECT 3.05 1.6 3.065 1.819 ;
      RECT 3.035 1.587 3.05 1.816 ;
      RECT 3.01 1.57 3.035 1.812 ;
      RECT 2.995 1.552 3.01 1.809 ;
      RECT 2.97 1.505 2.995 1.807 ;
      RECT 2.946 1.505 2.97 1.804 ;
      RECT 2.86 1.505 2.946 1.796 ;
      RECT 2.82 1.505 2.86 1.788 ;
      RECT 2.685 1.552 2.715 1.82 ;
      RECT 4.365 1.135 4.625 1.395 ;
      RECT 4.325 1.135 4.625 1.273 ;
      RECT 4.29 1.135 4.625 1.258 ;
      RECT 4.235 1.135 4.625 1.238 ;
      RECT 4.155 0.945 4.435 1.225 ;
      RECT 4.155 1.127 4.505 1.225 ;
      RECT 4.155 1.07 4.49 1.225 ;
      RECT 4.155 1.017 4.44 1.225 ;
      RECT 1.985 0.945 2.18 1.73 ;
      RECT 1.92 1.47 1.98 1.73 ;
      RECT 3.29 0.99 3.55 1.25 ;
      RECT 1.975 0.945 2.18 1.225 ;
      RECT 3.285 1 3.55 1.185 ;
      RECT 3 0.975 3.01 1.125 ;
      RECT 3.275 1 3.285 1.184 ;
      RECT 3.265 0.999 3.275 1.181 ;
      RECT 3.256 0.998 3.265 1.179 ;
      RECT 3.17 0.994 3.256 1.169 ;
      RECT 3.096 0.986 3.17 1.151 ;
      RECT 3.01 0.979 3.096 1.134 ;
      RECT 2.95 0.975 3 1.124 ;
      RECT 2.915 0.974 2.95 1.121 ;
      RECT 2.86 0.974 2.915 1.123 ;
      RECT 2.825 0.974 2.86 1.127 ;
      RECT 2.739 0.973 2.825 1.134 ;
      RECT 2.653 0.972 2.739 1.144 ;
      RECT 2.567 0.971 2.653 1.155 ;
      RECT 2.481 0.971 2.567 1.165 ;
      RECT 2.395 0.97 2.481 1.175 ;
      RECT 2.36 0.97 2.395 1.215 ;
      RECT 2.355 0.97 2.36 1.258 ;
      RECT 2.33 0.97 2.355 1.275 ;
      RECT 2.255 0.97 2.33 1.29 ;
      RECT 2.23 0.945 2.255 1.305 ;
      RECT 2.205 0.945 2.23 1.355 ;
      RECT 2.18 0.945 2.205 1.433 ;
      RECT 1.98 1.352 1.985 1.73 ;
      RECT 1.315 1.304 1.33 1.76 ;
      RECT 1.31 1.376 1.416 1.758 ;
      RECT 1.33 0.47 1.465 1.756 ;
      RECT 1.315 1.32 1.47 1.755 ;
      RECT 1.315 1.37 1.475 1.753 ;
      RECT 1.3 1.435 1.475 1.752 ;
      RECT 1.31 1.427 1.48 1.749 ;
      RECT 1.29 1.475 1.48 1.744 ;
      RECT 1.29 1.475 1.495 1.741 ;
      RECT 1.285 1.475 1.495 1.738 ;
      RECT 1.26 1.475 1.52 1.735 ;
      RECT 1.33 0.47 1.49 1.123 ;
      RECT 1.325 0.47 1.49 1.095 ;
      RECT 1.32 0.47 1.49 0.923 ;
      RECT 1.32 0.47 1.51 0.863 ;
      RECT 1.275 0.47 1.535 0.73 ;
      RECT 0.755 0.945 1.035 1.225 ;
      RECT 0.745 0.96 1.035 1.22 ;
      RECT 0.7 1.022 1.035 1.218 ;
      RECT 0.775 0.937 0.94 1.225 ;
      RECT 0.775 0.922 0.896 1.225 ;
      RECT 0.81 0.915 0.896 1.225 ;
      RECT 0.275 2.065 0.555 2.345 ;
      RECT 0.235 2.027 0.53 2.138 ;
      RECT 0.22 1.977 0.51 2.033 ;
      RECT 0.165 1.74 0.425 2 ;
      RECT 0.165 1.942 0.505 2 ;
      RECT 0.165 1.882 0.5 2 ;
      RECT 0.165 1.832 0.48 2 ;
      RECT 0.165 1.812 0.475 2 ;
      RECT 0.165 1.79 0.47 2 ;
      RECT 0.165 1.775 0.44 2 ;
    LAYER via1 ;
      RECT 10.605 0.57 10.755 0.72 ;
      RECT 9.655 2.075 9.805 2.225 ;
      RECT 9.205 0.575 9.355 0.725 ;
      RECT 9.025 1.565 9.175 1.715 ;
      RECT 8.63 2.08 8.78 2.23 ;
      RECT 8.27 2.035 8.42 2.185 ;
      RECT 8.125 0.525 8.275 0.675 ;
      RECT 7.54 1.975 7.69 2.125 ;
      RECT 7.445 0.51 7.595 0.66 ;
      RECT 7.29 1.045 7.44 1.195 ;
      RECT 6.605 2.01 6.755 2.16 ;
      RECT 6.21 0.635 6.36 0.785 ;
      RECT 5.49 1.54 5.64 1.69 ;
      RECT 5.45 0.575 5.6 0.725 ;
      RECT 5.18 2.045 5.33 2.195 ;
      RECT 4.645 0.765 4.795 0.915 ;
      RECT 4.6 1.635 4.75 1.785 ;
      RECT 4.42 1.19 4.57 1.34 ;
      RECT 3.345 1.045 3.495 1.195 ;
      RECT 3.24 0.47 3.39 0.62 ;
      RECT 2.585 1.615 2.735 1.765 ;
      RECT 1.975 1.525 2.125 1.675 ;
      RECT 1.33 0.525 1.48 0.675 ;
      RECT 1.315 1.53 1.465 1.68 ;
      RECT 0.8 1.015 0.95 1.165 ;
      RECT 0.22 1.795 0.37 1.945 ;
    LAYER met1 ;
      RECT 9.6 2.02 9.64 2.28 ;
      RECT 9.64 2 9.645 2.01 ;
      RECT 10.97 1.245 10.98 1.466 ;
      RECT 10.9 1.24 10.97 1.591 ;
      RECT 10.89 1.24 10.9 1.718 ;
      RECT 10.865 1.24 10.89 1.765 ;
      RECT 10.84 1.24 10.865 1.843 ;
      RECT 10.82 1.24 10.84 1.913 ;
      RECT 10.795 1.24 10.82 1.953 ;
      RECT 10.785 1.24 10.795 1.973 ;
      RECT 10.775 1.242 10.785 1.981 ;
      RECT 10.77 1.247 10.775 1.438 ;
      RECT 10.77 1.447 10.775 1.982 ;
      RECT 10.765 1.492 10.77 1.983 ;
      RECT 10.755 1.557 10.765 1.984 ;
      RECT 10.745 1.652 10.755 1.986 ;
      RECT 10.74 1.705 10.745 1.988 ;
      RECT 10.735 1.725 10.74 1.989 ;
      RECT 10.68 1.75 10.735 1.995 ;
      RECT 10.64 1.785 10.68 2.004 ;
      RECT 10.63 1.802 10.64 2.009 ;
      RECT 10.621 1.808 10.63 2.011 ;
      RECT 10.535 1.846 10.621 2.022 ;
      RECT 10.53 1.885 10.535 2.032 ;
      RECT 10.455 1.892 10.53 2.042 ;
      RECT 10.435 1.902 10.455 2.053 ;
      RECT 10.405 1.909 10.435 2.061 ;
      RECT 10.38 1.916 10.405 2.068 ;
      RECT 10.356 1.922 10.38 2.073 ;
      RECT 10.27 1.935 10.356 2.085 ;
      RECT 10.192 1.942 10.27 2.103 ;
      RECT 10.106 1.937 10.192 2.121 ;
      RECT 10.02 1.932 10.106 2.141 ;
      RECT 9.94 1.926 10.02 2.158 ;
      RECT 9.875 1.922 9.94 2.187 ;
      RECT 9.87 1.636 9.875 1.66 ;
      RECT 9.86 1.912 9.875 2.215 ;
      RECT 9.865 1.63 9.87 1.7 ;
      RECT 9.86 1.624 9.865 1.77 ;
      RECT 9.855 1.618 9.86 1.848 ;
      RECT 9.855 1.895 9.86 2.28 ;
      RECT 9.847 1.615 9.855 2.28 ;
      RECT 9.761 1.613 9.847 2.28 ;
      RECT 9.675 1.611 9.761 2.28 ;
      RECT 9.665 1.612 9.675 2.28 ;
      RECT 9.66 1.617 9.665 2.28 ;
      RECT 9.65 1.63 9.66 2.28 ;
      RECT 9.645 1.652 9.65 2.28 ;
      RECT 9.64 2.012 9.645 2.28 ;
      RECT 10.27 1.48 10.275 1.7 ;
      RECT 10.775 0.515 10.81 0.775 ;
      RECT 10.76 0.515 10.775 0.783 ;
      RECT 10.731 0.515 10.76 0.805 ;
      RECT 10.645 0.515 10.731 0.865 ;
      RECT 10.625 0.515 10.645 0.93 ;
      RECT 10.565 0.515 10.625 1.095 ;
      RECT 10.56 0.515 10.565 1.243 ;
      RECT 10.555 0.515 10.56 1.255 ;
      RECT 10.55 0.515 10.555 1.281 ;
      RECT 10.52 0.701 10.55 1.361 ;
      RECT 10.515 0.749 10.52 1.45 ;
      RECT 10.51 0.763 10.515 1.465 ;
      RECT 10.505 0.782 10.51 1.495 ;
      RECT 10.5 0.797 10.505 1.511 ;
      RECT 10.495 0.812 10.5 1.533 ;
      RECT 10.49 0.832 10.495 1.555 ;
      RECT 10.48 0.852 10.49 1.588 ;
      RECT 10.465 0.894 10.48 1.65 ;
      RECT 10.46 0.925 10.465 1.69 ;
      RECT 10.455 0.937 10.46 1.695 ;
      RECT 10.45 0.949 10.455 1.7 ;
      RECT 10.445 0.962 10.45 1.7 ;
      RECT 10.44 0.98 10.445 1.7 ;
      RECT 10.435 1 10.44 1.7 ;
      RECT 10.43 1.012 10.435 1.7 ;
      RECT 10.425 1.025 10.43 1.7 ;
      RECT 10.405 1.06 10.425 1.7 ;
      RECT 10.355 1.162 10.405 1.7 ;
      RECT 10.35 1.247 10.355 1.7 ;
      RECT 10.345 1.255 10.35 1.7 ;
      RECT 10.34 1.272 10.345 1.7 ;
      RECT 10.335 1.287 10.34 1.7 ;
      RECT 10.3 1.352 10.335 1.7 ;
      RECT 10.285 1.417 10.3 1.7 ;
      RECT 10.28 1.447 10.285 1.7 ;
      RECT 10.275 1.472 10.28 1.7 ;
      RECT 10.26 1.482 10.27 1.7 ;
      RECT 10.245 1.495 10.26 1.693 ;
      RECT 9.99 1.085 10.06 1.295 ;
      RECT 9.78 1.062 9.785 1.255 ;
      RECT 7.235 0.99 7.495 1.25 ;
      RECT 10.07 1.272 10.075 1.275 ;
      RECT 10.06 1.09 10.07 1.29 ;
      RECT 9.961 1.083 9.99 1.295 ;
      RECT 9.875 1.075 9.961 1.295 ;
      RECT 9.86 1.069 9.875 1.293 ;
      RECT 9.84 1.068 9.86 1.28 ;
      RECT 9.835 1.067 9.84 1.263 ;
      RECT 9.785 1.064 9.835 1.258 ;
      RECT 9.755 1.061 9.78 1.253 ;
      RECT 9.735 1.059 9.755 1.248 ;
      RECT 9.72 1.057 9.735 1.245 ;
      RECT 9.69 1.055 9.72 1.243 ;
      RECT 9.625 1.051 9.69 1.235 ;
      RECT 9.595 1.046 9.625 1.23 ;
      RECT 9.575 1.044 9.595 1.228 ;
      RECT 9.545 1.041 9.575 1.223 ;
      RECT 9.485 1.037 9.545 1.215 ;
      RECT 9.48 1.034 9.485 1.21 ;
      RECT 9.41 1.032 9.48 1.205 ;
      RECT 9.381 1.028 9.41 1.198 ;
      RECT 9.295 1.023 9.381 1.19 ;
      RECT 9.261 1.018 9.295 1.182 ;
      RECT 9.175 1.01 9.261 1.174 ;
      RECT 9.136 1.003 9.175 1.166 ;
      RECT 9.05 0.998 9.136 1.158 ;
      RECT 8.985 0.992 9.05 1.148 ;
      RECT 8.965 0.987 8.985 1.143 ;
      RECT 8.956 0.984 8.965 1.142 ;
      RECT 8.87 0.98 8.956 1.136 ;
      RECT 8.83 0.976 8.87 1.128 ;
      RECT 8.81 0.972 8.83 1.126 ;
      RECT 8.75 0.972 8.81 1.123 ;
      RECT 8.73 0.975 8.75 1.121 ;
      RECT 8.709 0.975 8.73 1.121 ;
      RECT 8.623 0.977 8.709 1.125 ;
      RECT 8.537 0.979 8.623 1.131 ;
      RECT 8.451 0.981 8.537 1.138 ;
      RECT 8.365 0.984 8.451 1.144 ;
      RECT 8.331 0.985 8.365 1.149 ;
      RECT 8.245 0.988 8.331 1.154 ;
      RECT 8.216 0.995 8.245 1.159 ;
      RECT 8.13 0.995 8.216 1.164 ;
      RECT 8.097 0.995 8.13 1.169 ;
      RECT 8.011 0.997 8.097 1.174 ;
      RECT 7.925 0.999 8.011 1.181 ;
      RECT 7.861 1.001 7.925 1.187 ;
      RECT 7.775 1.003 7.861 1.193 ;
      RECT 7.772 1.005 7.775 1.196 ;
      RECT 7.686 1.006 7.772 1.2 ;
      RECT 7.6 1.009 7.686 1.207 ;
      RECT 7.581 1.011 7.6 1.211 ;
      RECT 7.495 1.013 7.581 1.216 ;
      RECT 7.225 1.025 7.235 1.22 ;
      RECT 9.46 0.605 9.645 0.815 ;
      RECT 9.455 0.606 9.65 0.813 ;
      RECT 9.45 0.611 9.66 0.808 ;
      RECT 9.445 0.587 9.45 0.805 ;
      RECT 9.415 0.584 9.445 0.798 ;
      RECT 9.41 0.58 9.415 0.789 ;
      RECT 9.375 0.611 9.66 0.784 ;
      RECT 9.15 0.52 9.41 0.78 ;
      RECT 9.45 0.589 9.455 0.808 ;
      RECT 9.455 0.59 9.46 0.813 ;
      RECT 9.15 0.602 9.53 0.78 ;
      RECT 9.15 0.6 9.515 0.78 ;
      RECT 9.15 0.595 9.505 0.78 ;
      RECT 9.105 1.51 9.155 1.795 ;
      RECT 9.05 1.48 9.055 1.795 ;
      RECT 9.02 1.46 9.025 1.795 ;
      RECT 9.17 1.51 9.23 1.77 ;
      RECT 9.165 1.51 9.17 1.778 ;
      RECT 9.155 1.51 9.165 1.79 ;
      RECT 9.07 1.5 9.105 1.795 ;
      RECT 9.065 1.487 9.07 1.795 ;
      RECT 9.055 1.482 9.065 1.795 ;
      RECT 9.035 1.472 9.05 1.795 ;
      RECT 9.025 1.465 9.035 1.795 ;
      RECT 9.015 1.457 9.02 1.795 ;
      RECT 8.985 1.447 9.015 1.795 ;
      RECT 8.97 1.435 8.985 1.795 ;
      RECT 8.955 1.425 8.97 1.79 ;
      RECT 8.935 1.415 8.955 1.765 ;
      RECT 8.925 1.407 8.935 1.742 ;
      RECT 8.895 1.39 8.925 1.732 ;
      RECT 8.89 1.367 8.895 1.723 ;
      RECT 8.885 1.354 8.89 1.721 ;
      RECT 8.87 1.33 8.885 1.715 ;
      RECT 8.865 1.306 8.87 1.709 ;
      RECT 8.855 1.295 8.865 1.704 ;
      RECT 8.85 1.285 8.855 1.7 ;
      RECT 8.845 1.277 8.85 1.697 ;
      RECT 8.835 1.272 8.845 1.693 ;
      RECT 8.83 1.267 8.835 1.689 ;
      RECT 8.745 1.265 8.83 1.664 ;
      RECT 8.715 1.265 8.745 1.63 ;
      RECT 8.7 1.265 8.715 1.613 ;
      RECT 8.645 1.265 8.7 1.558 ;
      RECT 8.64 1.27 8.645 1.507 ;
      RECT 8.63 1.275 8.64 1.497 ;
      RECT 8.625 1.285 8.63 1.483 ;
      RECT 8.575 2.025 8.835 2.285 ;
      RECT 8.495 2.04 8.835 2.261 ;
      RECT 8.475 2.04 8.835 2.256 ;
      RECT 8.451 2.04 8.835 2.254 ;
      RECT 8.365 2.04 8.835 2.249 ;
      RECT 8.215 1.98 8.475 2.245 ;
      RECT 8.17 2.04 8.835 2.24 ;
      RECT 8.165 2.047 8.835 2.235 ;
      RECT 8.18 2.035 8.495 2.245 ;
      RECT 8.07 0.47 8.33 0.73 ;
      RECT 8.07 0.527 8.335 0.723 ;
      RECT 8.07 0.557 8.34 0.655 ;
      RECT 8.13 0.988 8.245 0.99 ;
      RECT 8.216 0.985 8.245 0.99 ;
      RECT 7.24 1.989 7.265 2.229 ;
      RECT 7.225 1.992 7.315 2.223 ;
      RECT 7.22 1.997 7.401 2.218 ;
      RECT 7.215 2.005 7.465 2.216 ;
      RECT 7.215 2.005 7.475 2.215 ;
      RECT 7.21 2.012 7.485 2.208 ;
      RECT 7.21 2.012 7.571 2.197 ;
      RECT 7.205 2.047 7.571 2.193 ;
      RECT 7.205 2.047 7.58 2.182 ;
      RECT 7.485 1.92 7.745 2.18 ;
      RECT 7.195 2.097 7.745 2.178 ;
      RECT 7.465 1.965 7.485 2.213 ;
      RECT 7.401 1.968 7.465 2.217 ;
      RECT 7.315 1.973 7.401 2.222 ;
      RECT 7.245 1.984 7.745 2.18 ;
      RECT 7.265 1.978 7.315 2.227 ;
      RECT 7.39 0.455 7.4 0.717 ;
      RECT 7.38 0.512 7.39 0.72 ;
      RECT 7.355 0.517 7.38 0.726 ;
      RECT 7.33 0.521 7.355 0.738 ;
      RECT 7.32 0.524 7.33 0.748 ;
      RECT 7.315 0.525 7.32 0.753 ;
      RECT 7.31 0.526 7.315 0.758 ;
      RECT 7.305 0.527 7.31 0.76 ;
      RECT 7.28 0.53 7.305 0.763 ;
      RECT 7.25 0.536 7.28 0.766 ;
      RECT 7.185 0.547 7.25 0.769 ;
      RECT 7.14 0.555 7.185 0.773 ;
      RECT 7.125 0.555 7.14 0.781 ;
      RECT 7.12 0.556 7.125 0.788 ;
      RECT 7.115 0.558 7.12 0.791 ;
      RECT 7.11 0.562 7.115 0.794 ;
      RECT 7.1 0.57 7.11 0.798 ;
      RECT 7.095 0.583 7.1 0.803 ;
      RECT 7.09 0.591 7.095 0.805 ;
      RECT 7.085 0.597 7.09 0.805 ;
      RECT 7.08 0.601 7.085 0.808 ;
      RECT 7.075 0.603 7.08 0.811 ;
      RECT 7.07 0.606 7.075 0.814 ;
      RECT 7.06 0.611 7.07 0.818 ;
      RECT 7.055 0.617 7.06 0.823 ;
      RECT 7.045 0.623 7.055 0.827 ;
      RECT 7.03 0.63 7.045 0.833 ;
      RECT 7.001 0.644 7.03 0.843 ;
      RECT 6.915 0.679 7.001 0.875 ;
      RECT 6.895 0.712 6.915 0.904 ;
      RECT 6.875 0.725 6.895 0.915 ;
      RECT 6.855 0.737 6.875 0.926 ;
      RECT 6.805 0.759 6.855 0.946 ;
      RECT 6.79 0.777 6.805 0.963 ;
      RECT 6.785 0.783 6.79 0.966 ;
      RECT 6.78 0.787 6.785 0.969 ;
      RECT 6.775 0.791 6.78 0.973 ;
      RECT 6.77 0.793 6.775 0.976 ;
      RECT 6.76 0.8 6.77 0.979 ;
      RECT 6.755 0.805 6.76 0.983 ;
      RECT 6.75 0.807 6.755 0.986 ;
      RECT 6.745 0.811 6.75 0.989 ;
      RECT 6.74 0.813 6.745 0.993 ;
      RECT 6.725 0.818 6.74 0.998 ;
      RECT 6.72 0.823 6.725 1.001 ;
      RECT 6.715 0.831 6.72 1.004 ;
      RECT 6.71 0.833 6.715 1.007 ;
      RECT 6.705 0.835 6.71 1.01 ;
      RECT 6.695 0.837 6.705 1.016 ;
      RECT 6.66 0.851 6.695 1.028 ;
      RECT 6.65 0.866 6.66 1.038 ;
      RECT 6.575 0.895 6.65 1.062 ;
      RECT 6.57 0.92 6.575 1.085 ;
      RECT 6.555 0.924 6.57 1.091 ;
      RECT 6.545 0.932 6.555 1.096 ;
      RECT 6.515 0.945 6.545 1.1 ;
      RECT 6.505 0.96 6.515 1.105 ;
      RECT 6.495 0.965 6.505 1.108 ;
      RECT 6.49 0.967 6.495 1.11 ;
      RECT 6.475 0.97 6.49 1.113 ;
      RECT 6.47 0.972 6.475 1.116 ;
      RECT 6.45 0.977 6.47 1.12 ;
      RECT 6.42 0.982 6.45 1.128 ;
      RECT 6.395 0.989 6.42 1.136 ;
      RECT 6.39 0.994 6.395 1.141 ;
      RECT 6.36 0.997 6.39 1.145 ;
      RECT 6.32 1 6.36 1.155 ;
      RECT 6.285 0.997 6.32 1.167 ;
      RECT 6.275 0.993 6.285 1.174 ;
      RECT 6.25 0.989 6.275 1.18 ;
      RECT 6.245 0.985 6.25 1.185 ;
      RECT 6.205 0.982 6.245 1.185 ;
      RECT 6.19 0.967 6.205 1.186 ;
      RECT 6.167 0.955 6.19 1.186 ;
      RECT 6.081 0.955 6.167 1.187 ;
      RECT 5.995 0.955 6.081 1.189 ;
      RECT 5.975 0.955 5.995 1.186 ;
      RECT 5.97 0.96 5.975 1.181 ;
      RECT 5.965 0.965 5.97 1.179 ;
      RECT 5.955 0.975 5.965 1.177 ;
      RECT 5.95 0.981 5.955 1.17 ;
      RECT 5.945 0.983 5.95 1.155 ;
      RECT 5.94 0.987 5.945 1.145 ;
      RECT 7.4 0.455 7.65 0.715 ;
      RECT 5.125 1.99 5.385 2.25 ;
      RECT 7.42 1.48 7.425 1.69 ;
      RECT 7.425 1.485 7.435 1.685 ;
      RECT 7.375 1.48 7.42 1.705 ;
      RECT 7.365 1.48 7.375 1.725 ;
      RECT 7.346 1.48 7.365 1.73 ;
      RECT 7.26 1.48 7.346 1.727 ;
      RECT 7.23 1.482 7.26 1.725 ;
      RECT 7.175 1.492 7.23 1.723 ;
      RECT 7.11 1.506 7.175 1.721 ;
      RECT 7.105 1.514 7.11 1.72 ;
      RECT 7.09 1.517 7.105 1.718 ;
      RECT 7.025 1.527 7.09 1.714 ;
      RECT 6.977 1.541 7.025 1.715 ;
      RECT 6.891 1.558 6.977 1.729 ;
      RECT 6.805 1.579 6.891 1.746 ;
      RECT 6.785 1.592 6.805 1.756 ;
      RECT 6.74 1.6 6.785 1.763 ;
      RECT 6.705 1.608 6.74 1.771 ;
      RECT 6.671 1.616 6.705 1.779 ;
      RECT 6.585 1.63 6.671 1.791 ;
      RECT 6.55 1.647 6.585 1.803 ;
      RECT 6.541 1.656 6.55 1.807 ;
      RECT 6.455 1.674 6.541 1.824 ;
      RECT 6.396 1.701 6.455 1.851 ;
      RECT 6.31 1.728 6.396 1.879 ;
      RECT 6.29 1.75 6.31 1.899 ;
      RECT 6.23 1.765 6.29 1.915 ;
      RECT 6.22 1.777 6.23 1.928 ;
      RECT 6.215 1.782 6.22 1.931 ;
      RECT 6.205 1.785 6.215 1.934 ;
      RECT 6.2 1.787 6.205 1.937 ;
      RECT 6.17 1.795 6.2 1.944 ;
      RECT 6.155 1.802 6.17 1.952 ;
      RECT 6.145 1.807 6.155 1.956 ;
      RECT 6.14 1.81 6.145 1.959 ;
      RECT 6.13 1.812 6.14 1.962 ;
      RECT 6.095 1.822 6.13 1.971 ;
      RECT 6.02 1.845 6.095 1.993 ;
      RECT 6 1.863 6.02 2.011 ;
      RECT 5.97 1.87 6 2.021 ;
      RECT 5.95 1.878 5.97 2.031 ;
      RECT 5.94 1.884 5.95 2.038 ;
      RECT 5.921 1.889 5.94 2.044 ;
      RECT 5.835 1.909 5.921 2.064 ;
      RECT 5.82 1.929 5.835 2.083 ;
      RECT 5.775 1.941 5.82 2.094 ;
      RECT 5.71 1.962 5.775 2.117 ;
      RECT 5.67 1.982 5.71 2.138 ;
      RECT 5.66 1.992 5.67 2.148 ;
      RECT 5.61 2.004 5.66 2.159 ;
      RECT 5.59 2.02 5.61 2.171 ;
      RECT 5.56 2.03 5.59 2.177 ;
      RECT 5.55 2.035 5.56 2.179 ;
      RECT 5.481 2.036 5.55 2.185 ;
      RECT 5.395 2.038 5.481 2.195 ;
      RECT 5.385 2.039 5.395 2.2 ;
      RECT 6.655 2.065 6.845 2.275 ;
      RECT 6.645 2.07 6.855 2.268 ;
      RECT 6.63 2.07 6.855 2.233 ;
      RECT 6.55 1.955 6.81 2.215 ;
      RECT 5.465 1.485 5.65 1.78 ;
      RECT 5.455 1.485 5.65 1.778 ;
      RECT 5.44 1.485 5.655 1.773 ;
      RECT 5.44 1.485 5.66 1.77 ;
      RECT 5.435 1.485 5.66 1.768 ;
      RECT 5.43 1.74 5.66 1.758 ;
      RECT 5.435 1.485 5.695 1.745 ;
      RECT 5.395 0.52 5.655 0.78 ;
      RECT 5.205 0.445 5.291 0.778 ;
      RECT 5.18 0.449 5.335 0.774 ;
      RECT 5.291 0.441 5.335 0.774 ;
      RECT 5.291 0.442 5.34 0.773 ;
      RECT 5.205 0.447 5.355 0.772 ;
      RECT 5.18 0.455 5.395 0.771 ;
      RECT 5.175 0.45 5.355 0.766 ;
      RECT 5.165 0.465 5.395 0.673 ;
      RECT 5.165 0.517 5.595 0.673 ;
      RECT 5.165 0.51 5.575 0.673 ;
      RECT 5.165 0.497 5.545 0.673 ;
      RECT 5.165 0.485 5.485 0.673 ;
      RECT 5.165 0.47 5.46 0.673 ;
      RECT 4.365 1.1 4.5 1.395 ;
      RECT 4.625 1.123 4.63 1.31 ;
      RECT 5.345 1.02 5.49 1.255 ;
      RECT 5.505 1.02 5.51 1.245 ;
      RECT 5.54 1.031 5.545 1.225 ;
      RECT 5.535 1.023 5.54 1.23 ;
      RECT 5.515 1.02 5.535 1.235 ;
      RECT 5.51 1.02 5.515 1.243 ;
      RECT 5.5 1.02 5.505 1.248 ;
      RECT 5.49 1.02 5.5 1.253 ;
      RECT 5.32 1.022 5.345 1.255 ;
      RECT 5.27 1.029 5.32 1.255 ;
      RECT 5.265 1.034 5.27 1.255 ;
      RECT 5.226 1.039 5.265 1.256 ;
      RECT 5.14 1.051 5.226 1.257 ;
      RECT 5.131 1.061 5.14 1.257 ;
      RECT 5.045 1.07 5.131 1.259 ;
      RECT 5.021 1.08 5.045 1.261 ;
      RECT 4.935 1.091 5.021 1.262 ;
      RECT 4.905 1.102 4.935 1.264 ;
      RECT 4.875 1.107 4.905 1.266 ;
      RECT 4.85 1.113 4.875 1.269 ;
      RECT 4.835 1.118 4.85 1.27 ;
      RECT 4.79 1.124 4.835 1.27 ;
      RECT 4.785 1.129 4.79 1.271 ;
      RECT 4.765 1.129 4.785 1.273 ;
      RECT 4.745 1.127 4.765 1.278 ;
      RECT 4.71 1.126 4.745 1.285 ;
      RECT 4.68 1.125 4.71 1.295 ;
      RECT 4.63 1.124 4.68 1.305 ;
      RECT 4.54 1.121 4.625 1.395 ;
      RECT 4.515 1.115 4.54 1.395 ;
      RECT 4.5 1.105 4.515 1.395 ;
      RECT 4.315 1.1 4.365 1.315 ;
      RECT 4.305 1.105 4.315 1.305 ;
      RECT 4.545 1.58 4.805 1.84 ;
      RECT 4.545 1.58 4.835 1.733 ;
      RECT 4.545 1.58 4.87 1.718 ;
      RECT 4.8 1.5 4.99 1.71 ;
      RECT 4.79 1.505 5 1.703 ;
      RECT 4.755 1.575 5 1.703 ;
      RECT 4.785 1.517 4.805 1.84 ;
      RECT 4.77 1.565 5 1.703 ;
      RECT 4.775 1.537 4.805 1.84 ;
      RECT 3.855 0.605 3.925 1.71 ;
      RECT 4.59 0.71 4.85 0.97 ;
      RECT 4.17 0.756 4.185 0.965 ;
      RECT 4.506 0.769 4.59 0.92 ;
      RECT 4.42 0.766 4.506 0.92 ;
      RECT 4.381 0.764 4.42 0.92 ;
      RECT 4.295 0.762 4.381 0.92 ;
      RECT 4.235 0.76 4.295 0.931 ;
      RECT 4.2 0.758 4.235 0.949 ;
      RECT 4.185 0.756 4.2 0.96 ;
      RECT 4.155 0.756 4.17 0.973 ;
      RECT 4.145 0.756 4.155 0.978 ;
      RECT 4.12 0.755 4.145 0.983 ;
      RECT 4.105 0.75 4.12 0.989 ;
      RECT 4.1 0.743 4.105 0.994 ;
      RECT 4.075 0.734 4.1 1 ;
      RECT 4.03 0.713 4.075 1.013 ;
      RECT 4.02 0.697 4.03 1.023 ;
      RECT 4.005 0.69 4.02 1.033 ;
      RECT 3.995 0.683 4.005 1.05 ;
      RECT 3.99 0.68 3.995 1.08 ;
      RECT 3.985 0.678 3.99 1.11 ;
      RECT 3.98 0.676 3.985 1.147 ;
      RECT 3.965 0.672 3.98 1.214 ;
      RECT 3.965 1.505 3.975 1.705 ;
      RECT 3.96 0.668 3.965 1.34 ;
      RECT 3.96 1.492 3.965 1.71 ;
      RECT 3.955 0.666 3.96 1.425 ;
      RECT 3.955 1.482 3.96 1.71 ;
      RECT 3.94 0.637 3.955 1.71 ;
      RECT 3.925 0.61 3.94 1.71 ;
      RECT 3.85 0.605 3.855 0.96 ;
      RECT 3.85 1.015 3.855 1.71 ;
      RECT 3.835 0.605 3.85 0.938 ;
      RECT 3.845 1.037 3.85 1.71 ;
      RECT 3.835 1.077 3.845 1.71 ;
      RECT 3.8 0.605 3.835 0.88 ;
      RECT 3.83 1.112 3.835 1.71 ;
      RECT 3.815 1.167 3.83 1.71 ;
      RECT 3.81 1.232 3.815 1.71 ;
      RECT 3.795 1.28 3.81 1.71 ;
      RECT 3.77 0.605 3.8 0.835 ;
      RECT 3.79 1.335 3.795 1.71 ;
      RECT 3.775 1.395 3.79 1.71 ;
      RECT 3.77 1.443 3.775 1.708 ;
      RECT 3.765 0.605 3.77 0.828 ;
      RECT 3.765 1.475 3.77 1.703 ;
      RECT 3.74 0.605 3.765 0.82 ;
      RECT 3.73 0.61 3.74 0.81 ;
      RECT 3.945 1.885 3.965 2.125 ;
      RECT 3.175 1.815 3.18 2.025 ;
      RECT 4.455 1.888 4.465 2.083 ;
      RECT 4.45 1.878 4.455 2.086 ;
      RECT 4.37 1.875 4.45 2.109 ;
      RECT 4.366 1.875 4.37 2.131 ;
      RECT 4.28 1.875 4.366 2.141 ;
      RECT 4.265 1.875 4.28 2.149 ;
      RECT 4.236 1.876 4.265 2.147 ;
      RECT 4.15 1.881 4.236 2.143 ;
      RECT 4.137 1.885 4.15 2.139 ;
      RECT 4.051 1.885 4.137 2.135 ;
      RECT 3.965 1.885 4.051 2.129 ;
      RECT 3.881 1.885 3.945 2.123 ;
      RECT 3.795 1.885 3.881 2.118 ;
      RECT 3.775 1.885 3.795 2.114 ;
      RECT 3.715 1.88 3.775 2.111 ;
      RECT 3.687 1.874 3.715 2.108 ;
      RECT 3.601 1.869 3.687 2.104 ;
      RECT 3.515 1.863 3.601 2.098 ;
      RECT 3.44 1.845 3.515 2.093 ;
      RECT 3.405 1.822 3.44 2.089 ;
      RECT 3.395 1.812 3.405 2.088 ;
      RECT 3.34 1.81 3.395 2.087 ;
      RECT 3.265 1.81 3.34 2.083 ;
      RECT 3.255 1.81 3.265 2.078 ;
      RECT 3.24 1.81 3.255 2.07 ;
      RECT 3.19 1.812 3.24 2.048 ;
      RECT 3.18 1.815 3.19 2.028 ;
      RECT 3.17 1.82 3.175 2.023 ;
      RECT 3.165 1.825 3.17 2.018 ;
      RECT 3.29 0.99 3.55 1.25 ;
      RECT 3.29 1.005 3.57 1.215 ;
      RECT 3.29 1.01 3.58 1.21 ;
      RECT 1.275 0.47 1.535 0.73 ;
      RECT 1.265 0.5 1.535 0.71 ;
      RECT 3.185 0.415 3.445 0.675 ;
      RECT 3.18 0.49 3.185 0.676 ;
      RECT 3.155 0.495 3.18 0.678 ;
      RECT 3.14 0.502 3.155 0.681 ;
      RECT 3.08 0.52 3.14 0.686 ;
      RECT 3.05 0.54 3.08 0.693 ;
      RECT 3.025 0.548 3.05 0.698 ;
      RECT 3 0.556 3.025 0.7 ;
      RECT 2.982 0.56 3 0.699 ;
      RECT 2.896 0.558 2.982 0.699 ;
      RECT 2.81 0.556 2.896 0.699 ;
      RECT 2.724 0.554 2.81 0.698 ;
      RECT 2.638 0.552 2.724 0.698 ;
      RECT 2.552 0.55 2.638 0.698 ;
      RECT 2.466 0.548 2.552 0.698 ;
      RECT 2.38 0.546 2.466 0.697 ;
      RECT 2.362 0.545 2.38 0.697 ;
      RECT 2.276 0.544 2.362 0.697 ;
      RECT 2.19 0.542 2.276 0.697 ;
      RECT 2.104 0.541 2.19 0.696 ;
      RECT 2.018 0.54 2.104 0.696 ;
      RECT 1.932 0.538 2.018 0.696 ;
      RECT 1.846 0.537 1.932 0.696 ;
      RECT 1.76 0.535 1.846 0.695 ;
      RECT 1.736 0.533 1.76 0.695 ;
      RECT 1.65 0.526 1.736 0.695 ;
      RECT 1.621 0.518 1.65 0.695 ;
      RECT 1.535 0.51 1.621 0.695 ;
      RECT 1.255 0.507 1.265 0.705 ;
      RECT 2.76 1.47 2.765 1.82 ;
      RECT 2.53 1.56 2.67 1.82 ;
      RECT 3.005 1.245 3.05 1.455 ;
      RECT 3.06 1.256 3.07 1.45 ;
      RECT 3.05 1.248 3.06 1.455 ;
      RECT 2.985 1.245 3.005 1.46 ;
      RECT 2.955 1.245 2.985 1.483 ;
      RECT 2.945 1.245 2.955 1.508 ;
      RECT 2.94 1.245 2.945 1.518 ;
      RECT 2.885 1.245 2.94 1.558 ;
      RECT 2.88 1.245 2.885 1.598 ;
      RECT 2.875 1.247 2.88 1.603 ;
      RECT 2.86 1.257 2.875 1.614 ;
      RECT 2.815 1.315 2.86 1.65 ;
      RECT 2.805 1.37 2.815 1.684 ;
      RECT 2.79 1.397 2.805 1.7 ;
      RECT 2.78 1.424 2.79 1.82 ;
      RECT 2.765 1.447 2.78 1.82 ;
      RECT 2.755 1.487 2.76 1.82 ;
      RECT 2.75 1.497 2.755 1.82 ;
      RECT 2.745 1.512 2.75 1.82 ;
      RECT 2.735 1.517 2.745 1.82 ;
      RECT 2.67 1.54 2.735 1.82 ;
      RECT 2.17 1.035 2.36 1.245 ;
      RECT 0.745 0.96 1.005 1.22 ;
      RECT 1.095 0.955 1.19 1.165 ;
      RECT 1.07 0.97 1.08 1.165 ;
      RECT 2.36 1.042 2.37 1.24 ;
      RECT 2.16 1.042 2.17 1.24 ;
      RECT 2.145 1.057 2.16 1.23 ;
      RECT 2.14 1.065 2.145 1.223 ;
      RECT 2.13 1.068 2.14 1.22 ;
      RECT 2.095 1.067 2.13 1.218 ;
      RECT 2.066 1.063 2.095 1.215 ;
      RECT 1.98 1.058 2.066 1.212 ;
      RECT 1.92 1.052 1.98 1.208 ;
      RECT 1.891 1.048 1.92 1.205 ;
      RECT 1.805 1.04 1.891 1.202 ;
      RECT 1.796 1.034 1.805 1.2 ;
      RECT 1.71 1.029 1.796 1.198 ;
      RECT 1.687 1.024 1.71 1.195 ;
      RECT 1.601 1.018 1.687 1.192 ;
      RECT 1.515 1.009 1.601 1.187 ;
      RECT 1.505 1.004 1.515 1.185 ;
      RECT 1.486 1.003 1.505 1.184 ;
      RECT 1.4 0.998 1.486 1.18 ;
      RECT 1.38 0.993 1.4 1.176 ;
      RECT 1.32 0.988 1.38 1.173 ;
      RECT 1.295 0.978 1.32 1.171 ;
      RECT 1.29 0.971 1.295 1.17 ;
      RECT 1.28 0.962 1.29 1.169 ;
      RECT 1.276 0.955 1.28 1.169 ;
      RECT 1.19 0.955 1.276 1.167 ;
      RECT 1.08 0.962 1.095 1.165 ;
      RECT 1.065 0.972 1.07 1.165 ;
      RECT 1.045 0.975 1.065 1.162 ;
      RECT 1.015 0.975 1.045 1.158 ;
      RECT 1.005 0.975 1.015 1.158 ;
      RECT 1.92 1.47 2.18 1.73 ;
      RECT 1.85 1.48 2.18 1.69 ;
      RECT 1.84 1.487 2.18 1.685 ;
      RECT 1.26 1.475 1.52 1.735 ;
      RECT 1.26 1.515 1.625 1.725 ;
      RECT 1.26 1.517 1.63 1.724 ;
      RECT 1.26 1.525 1.635 1.721 ;
      RECT 0.185 0.6 0.285 2.125 ;
      RECT 0.375 1.74 0.425 2 ;
      RECT 0.37 0.613 0.375 0.8 ;
      RECT 0.365 1.721 0.375 2 ;
      RECT 0.365 0.61 0.37 0.808 ;
      RECT 0.35 0.604 0.365 0.815 ;
      RECT 0.36 1.709 0.365 2.083 ;
      RECT 0.35 1.697 0.36 2.12 ;
      RECT 0.34 0.6 0.35 0.822 ;
      RECT 0.34 1.682 0.35 2.125 ;
      RECT 0.335 0.6 0.34 0.83 ;
      RECT 0.315 1.652 0.34 2.125 ;
      RECT 0.295 0.6 0.335 0.878 ;
      RECT 0.305 1.612 0.315 2.125 ;
      RECT 0.295 1.567 0.305 2.125 ;
      RECT 0.29 0.6 0.295 0.948 ;
      RECT 0.29 1.525 0.295 2.125 ;
      RECT 0.285 0.6 0.29 1.425 ;
      RECT 0.285 1.507 0.29 2.125 ;
      RECT 0.175 0.603 0.185 2.125 ;
      RECT 0.16 0.61 0.175 2.121 ;
      RECT 0.155 0.62 0.16 2.116 ;
      RECT 0.15 0.82 0.155 2.008 ;
      RECT 0.145 0.905 0.15 1.56 ;
      RECT 0 -0.235 11.96 0.245 ;
      RECT 0 2.485 11.96 2.965 ;
      RECT 6.155 0.58 6.415 0.84 ;
    LAYER mcon ;
      RECT 11.645 -0.08 11.815 0.09 ;
      RECT 11.645 2.64 11.815 2.81 ;
      RECT 11.185 -0.08 11.355 0.09 ;
      RECT 11.185 2.64 11.355 2.81 ;
      RECT 10.79 1.26 10.96 1.43 ;
      RECT 10.725 -0.08 10.895 0.09 ;
      RECT 10.725 2.64 10.895 2.81 ;
      RECT 10.58 0.6 10.75 0.77 ;
      RECT 10.265 -0.08 10.435 0.09 ;
      RECT 10.265 1.51 10.435 1.68 ;
      RECT 10.265 2.64 10.435 2.81 ;
      RECT 9.88 1.105 10.05 1.275 ;
      RECT 9.805 -0.08 9.975 0.09 ;
      RECT 9.805 2.64 9.975 2.81 ;
      RECT 9.665 1.67 9.835 1.84 ;
      RECT 9.645 2.07 9.815 2.24 ;
      RECT 9.47 0.625 9.64 0.795 ;
      RECT 9.345 -0.08 9.515 0.09 ;
      RECT 9.345 2.64 9.515 2.81 ;
      RECT 8.975 1.605 9.145 1.775 ;
      RECT 8.885 -0.08 9.055 0.09 ;
      RECT 8.885 2.64 9.055 2.81 ;
      RECT 8.65 1.29 8.82 1.46 ;
      RECT 8.585 2.07 8.755 2.24 ;
      RECT 8.425 -0.08 8.595 0.09 ;
      RECT 8.425 2.64 8.595 2.81 ;
      RECT 8.185 2.055 8.355 2.225 ;
      RECT 8.145 0.54 8.315 0.71 ;
      RECT 7.965 -0.08 8.135 0.09 ;
      RECT 7.965 2.64 8.135 2.81 ;
      RECT 7.505 -0.08 7.675 0.09 ;
      RECT 7.505 2.64 7.675 2.81 ;
      RECT 7.245 1.04 7.415 1.21 ;
      RECT 7.245 1.5 7.415 1.67 ;
      RECT 7.245 2.015 7.415 2.185 ;
      RECT 7.13 0.575 7.3 0.745 ;
      RECT 7.045 -0.08 7.215 0.09 ;
      RECT 7.045 2.64 7.215 2.81 ;
      RECT 6.665 2.085 6.835 2.255 ;
      RECT 6.585 -0.08 6.755 0.09 ;
      RECT 6.585 2.64 6.755 2.81 ;
      RECT 6.185 0.615 6.355 0.785 ;
      RECT 6.125 -0.08 6.295 0.09 ;
      RECT 6.125 2.64 6.295 2.81 ;
      RECT 5.97 0.99 6.14 1.16 ;
      RECT 5.665 -0.08 5.835 0.09 ;
      RECT 5.665 2.64 5.835 2.81 ;
      RECT 5.47 1.59 5.64 1.76 ;
      RECT 5.355 1.04 5.525 1.21 ;
      RECT 5.205 -0.08 5.375 0.09 ;
      RECT 5.205 2.64 5.375 2.81 ;
      RECT 5.185 0.49 5.355 0.66 ;
      RECT 4.81 1.52 4.98 1.69 ;
      RECT 4.745 -0.08 4.915 0.09 ;
      RECT 4.745 2.64 4.915 2.81 ;
      RECT 4.325 1.12 4.495 1.29 ;
      RECT 4.285 -0.08 4.455 0.09 ;
      RECT 4.285 2.64 4.455 2.81 ;
      RECT 4.275 1.895 4.445 2.065 ;
      RECT 3.825 -0.08 3.995 0.09 ;
      RECT 3.825 2.64 3.995 2.81 ;
      RECT 3.785 1.52 3.955 1.69 ;
      RECT 3.75 0.625 3.92 0.795 ;
      RECT 3.39 1.025 3.56 1.195 ;
      RECT 3.365 -0.08 3.535 0.09 ;
      RECT 3.365 2.64 3.535 2.81 ;
      RECT 3.185 1.835 3.355 2.005 ;
      RECT 2.905 -0.08 3.075 0.09 ;
      RECT 2.905 2.64 3.075 2.81 ;
      RECT 2.88 1.265 3.05 1.435 ;
      RECT 2.445 -0.08 2.615 0.09 ;
      RECT 2.445 2.64 2.615 2.81 ;
      RECT 2.18 1.055 2.35 1.225 ;
      RECT 1.985 -0.08 2.155 0.09 ;
      RECT 1.985 2.64 2.155 2.81 ;
      RECT 1.86 1.5 2.03 1.67 ;
      RECT 1.525 -0.08 1.695 0.09 ;
      RECT 1.525 2.64 1.695 2.81 ;
      RECT 1.445 1.535 1.615 1.705 ;
      RECT 1.275 0.52 1.445 0.69 ;
      RECT 1.1 0.975 1.27 1.145 ;
      RECT 1.065 -0.08 1.235 0.09 ;
      RECT 1.065 2.64 1.235 2.81 ;
      RECT 0.605 -0.08 0.775 0.09 ;
      RECT 0.605 2.64 0.775 2.81 ;
      RECT 0.18 0.625 0.35 0.795 ;
      RECT 0.175 1.94 0.345 2.11 ;
      RECT 0.145 -0.08 0.315 0.09 ;
      RECT 0.145 2.64 0.315 2.81 ;
    LAYER li ;
      RECT 11.05 -0.08 11.22 0.59 ;
      RECT 10.09 -0.08 10.26 0.59 ;
      RECT 9.13 -0.08 9.3 0.59 ;
      RECT 8.61 -0.08 8.78 0.59 ;
      RECT 7.65 -0.08 7.82 0.59 ;
      RECT 6.65 -0.08 6.82 0.59 ;
      RECT 5.69 -0.08 5.86 0.59 ;
      RECT 4.21 -0.08 4.38 0.59 ;
      RECT 2.29 -0.08 2.46 0.59 ;
      RECT 0.81 -0.08 0.98 0.59 ;
      RECT 0 -0.08 11.96 0.09 ;
      RECT 0 2.64 11.96 2.81 ;
      RECT 10.09 2.14 10.26 2.81 ;
      RECT 7.65 2.14 7.82 2.81 ;
      RECT 5.69 2.14 5.86 2.81 ;
      RECT 4.73 2.14 4.9 2.81 ;
      RECT 2.77 2.14 2.94 2.81 ;
      RECT 1.77 2.14 1.94 2.81 ;
      RECT 0.81 2.14 0.98 2.81 ;
      RECT 11.375 1.747 11.39 1.798 ;
      RECT 11.37 1.727 11.375 1.845 ;
      RECT 11.355 1.717 11.37 1.913 ;
      RECT 11.33 1.697 11.355 1.968 ;
      RECT 11.29 1.682 11.33 1.988 ;
      RECT 11.245 1.676 11.29 2.016 ;
      RECT 11.175 1.666 11.245 2.033 ;
      RECT 11.155 1.658 11.175 2.033 ;
      RECT 11.095 1.652 11.155 2.025 ;
      RECT 11.036 1.643 11.095 2.013 ;
      RECT 10.95 1.632 11.036 1.996 ;
      RECT 10.928 1.623 10.95 1.984 ;
      RECT 10.842 1.616 10.928 1.971 ;
      RECT 10.756 1.603 10.842 1.952 ;
      RECT 10.67 1.591 10.756 1.932 ;
      RECT 10.64 1.58 10.67 1.919 ;
      RECT 10.59 1.566 10.64 1.911 ;
      RECT 10.57 1.555 10.59 1.903 ;
      RECT 10.521 1.544 10.57 1.895 ;
      RECT 10.435 1.523 10.521 1.88 ;
      RECT 10.39 1.51 10.435 1.865 ;
      RECT 10.345 1.51 10.39 1.845 ;
      RECT 10.29 1.51 10.345 1.78 ;
      RECT 10.265 1.51 10.29 1.703 ;
      RECT 10.79 1.247 10.96 1.43 ;
      RECT 10.79 1.247 10.975 1.388 ;
      RECT 10.79 1.247 10.98 1.33 ;
      RECT 10.85 1.015 10.985 1.306 ;
      RECT 10.85 1.019 10.99 1.289 ;
      RECT 10.795 1.182 10.99 1.289 ;
      RECT 10.82 1.027 10.96 1.43 ;
      RECT 10.82 1.031 11 1.23 ;
      RECT 10.805 1.117 11 1.23 ;
      RECT 10.815 1.047 10.96 1.43 ;
      RECT 10.815 1.05 11.01 1.143 ;
      RECT 10.81 1.067 11.01 1.143 ;
      RECT 10.58 0.287 10.75 0.77 ;
      RECT 10.575 0.282 10.725 0.76 ;
      RECT 10.575 0.289 10.755 0.754 ;
      RECT 10.565 0.283 10.725 0.733 ;
      RECT 10.565 0.299 10.77 0.692 ;
      RECT 10.535 0.284 10.725 0.655 ;
      RECT 10.535 0.314 10.78 0.595 ;
      RECT 10.53 0.286 10.725 0.593 ;
      RECT 10.51 0.295 10.755 0.55 ;
      RECT 10.485 0.311 10.77 0.462 ;
      RECT 10.485 0.33 10.795 0.453 ;
      RECT 10.48 0.367 10.795 0.405 ;
      RECT 10.485 0.347 10.8 0.373 ;
      RECT 10.58 0.281 10.69 0.77 ;
      RECT 10.666 0.28 10.69 0.77 ;
      RECT 9.9 1.065 9.905 1.276 ;
      RECT 10.5 1.065 10.505 1.25 ;
      RECT 10.565 1.105 10.57 1.218 ;
      RECT 10.56 1.097 10.565 1.224 ;
      RECT 10.555 1.087 10.56 1.232 ;
      RECT 10.55 1.077 10.555 1.241 ;
      RECT 10.545 1.067 10.55 1.245 ;
      RECT 10.505 1.065 10.545 1.248 ;
      RECT 10.477 1.064 10.5 1.252 ;
      RECT 10.391 1.061 10.477 1.259 ;
      RECT 10.305 1.057 10.391 1.27 ;
      RECT 10.285 1.055 10.305 1.276 ;
      RECT 10.267 1.054 10.285 1.279 ;
      RECT 10.181 1.052 10.267 1.286 ;
      RECT 10.095 1.047 10.181 1.299 ;
      RECT 10.076 1.044 10.095 1.304 ;
      RECT 9.99 1.042 10.076 1.295 ;
      RECT 9.98 1.042 9.99 1.288 ;
      RECT 9.905 1.055 9.98 1.282 ;
      RECT 9.89 1.066 9.9 1.276 ;
      RECT 9.88 1.068 9.89 1.275 ;
      RECT 9.87 1.072 9.88 1.271 ;
      RECT 9.865 1.075 9.87 1.265 ;
      RECT 9.855 1.077 9.865 1.259 ;
      RECT 9.85 1.08 9.855 1.253 ;
      RECT 9.83 1.666 9.835 1.87 ;
      RECT 9.815 1.653 9.83 1.963 ;
      RECT 9.8 1.634 9.815 2.24 ;
      RECT 9.765 1.6 9.8 2.24 ;
      RECT 9.761 1.57 9.765 2.24 ;
      RECT 9.675 1.452 9.761 2.24 ;
      RECT 9.665 1.327 9.675 2.24 ;
      RECT 9.65 1.295 9.665 2.24 ;
      RECT 9.645 1.27 9.65 2.24 ;
      RECT 9.64 1.26 9.645 2.196 ;
      RECT 9.625 1.232 9.64 2.101 ;
      RECT 9.61 1.198 9.625 2 ;
      RECT 9.605 1.176 9.61 1.953 ;
      RECT 9.6 1.165 9.605 1.923 ;
      RECT 9.595 1.155 9.6 1.889 ;
      RECT 9.585 1.142 9.595 1.857 ;
      RECT 9.56 1.118 9.585 1.783 ;
      RECT 9.555 1.098 9.56 1.708 ;
      RECT 9.55 1.092 9.555 1.683 ;
      RECT 9.545 1.087 9.55 1.648 ;
      RECT 9.54 1.082 9.545 1.623 ;
      RECT 9.535 1.08 9.54 1.603 ;
      RECT 9.53 1.08 9.535 1.588 ;
      RECT 9.525 1.08 9.53 1.548 ;
      RECT 9.515 1.08 9.525 1.52 ;
      RECT 9.505 1.08 9.515 1.465 ;
      RECT 9.49 1.08 9.505 1.403 ;
      RECT 9.485 1.079 9.49 1.348 ;
      RECT 9.47 1.078 9.485 1.328 ;
      RECT 9.41 1.076 9.47 1.302 ;
      RECT 9.375 1.077 9.41 1.282 ;
      RECT 9.37 1.079 9.375 1.272 ;
      RECT 9.36 1.098 9.37 1.262 ;
      RECT 9.355 1.125 9.36 1.193 ;
      RECT 9.47 0.55 9.64 0.795 ;
      RECT 9.505 0.321 9.64 0.795 ;
      RECT 9.505 0.323 9.65 0.79 ;
      RECT 9.505 0.325 9.675 0.778 ;
      RECT 9.505 0.328 9.7 0.76 ;
      RECT 9.505 0.333 9.75 0.733 ;
      RECT 9.505 0.338 9.77 0.698 ;
      RECT 9.485 0.34 9.78 0.673 ;
      RECT 9.475 0.435 9.78 0.673 ;
      RECT 9.505 0.32 9.615 0.795 ;
      RECT 9.515 0.317 9.61 0.795 ;
      RECT 9.035 1.582 9.225 1.94 ;
      RECT 9.035 1.594 9.26 1.939 ;
      RECT 9.035 1.622 9.28 1.937 ;
      RECT 9.035 1.647 9.285 1.936 ;
      RECT 9.035 1.705 9.3 1.935 ;
      RECT 9.02 1.578 9.18 1.92 ;
      RECT 9 1.587 9.225 1.873 ;
      RECT 8.975 1.598 9.26 1.81 ;
      RECT 8.975 1.682 9.295 1.81 ;
      RECT 8.975 1.657 9.29 1.81 ;
      RECT 9.035 1.573 9.18 1.94 ;
      RECT 9.121 1.572 9.18 1.94 ;
      RECT 9.121 1.571 9.165 1.94 ;
      RECT 8.82 1.087 8.825 1.465 ;
      RECT 8.815 1.055 8.82 1.465 ;
      RECT 8.81 1.027 8.815 1.465 ;
      RECT 8.805 1.007 8.81 1.465 ;
      RECT 8.75 0.99 8.805 1.465 ;
      RECT 8.71 0.975 8.75 1.465 ;
      RECT 8.655 0.962 8.71 1.465 ;
      RECT 8.62 0.953 8.655 1.465 ;
      RECT 8.616 0.951 8.62 1.464 ;
      RECT 8.53 0.947 8.616 1.447 ;
      RECT 8.445 0.939 8.53 1.41 ;
      RECT 8.435 0.935 8.445 1.383 ;
      RECT 8.425 0.935 8.435 1.365 ;
      RECT 8.415 0.937 8.425 1.348 ;
      RECT 8.41 0.942 8.415 1.334 ;
      RECT 8.405 0.946 8.41 1.321 ;
      RECT 8.395 0.951 8.405 1.305 ;
      RECT 8.38 0.965 8.395 1.28 ;
      RECT 8.375 0.971 8.38 1.26 ;
      RECT 8.37 0.973 8.375 1.253 ;
      RECT 8.365 0.977 8.37 1.128 ;
      RECT 8.545 1.777 8.79 2.24 ;
      RECT 8.465 1.75 8.785 2.236 ;
      RECT 8.395 1.785 8.79 2.229 ;
      RECT 8.185 2.04 8.79 2.225 ;
      RECT 8.365 1.808 8.79 2.225 ;
      RECT 8.205 2 8.79 2.225 ;
      RECT 8.355 1.82 8.79 2.225 ;
      RECT 8.24 1.937 8.79 2.225 ;
      RECT 8.295 1.862 8.79 2.225 ;
      RECT 8.545 1.727 8.785 2.24 ;
      RECT 8.575 1.72 8.785 2.24 ;
      RECT 8.565 1.722 8.785 2.24 ;
      RECT 8.575 1.717 8.705 2.24 ;
      RECT 8.13 0.28 8.216 0.719 ;
      RECT 8.125 0.28 8.216 0.717 ;
      RECT 8.125 0.28 8.285 0.716 ;
      RECT 8.125 0.28 8.315 0.713 ;
      RECT 8.11 0.287 8.315 0.704 ;
      RECT 8.11 0.287 8.32 0.7 ;
      RECT 8.105 0.297 8.32 0.693 ;
      RECT 8.1 0.302 8.32 0.668 ;
      RECT 8.1 0.302 8.335 0.65 ;
      RECT 8.125 0.28 8.355 0.565 ;
      RECT 8.095 0.307 8.355 0.563 ;
      RECT 8.105 0.3 8.36 0.501 ;
      RECT 8.095 0.422 8.365 0.484 ;
      RECT 8.08 0.317 8.36 0.435 ;
      RECT 8.075 0.327 8.36 0.335 ;
      RECT 8.155 1.098 8.16 1.175 ;
      RECT 8.145 1.092 8.155 1.365 ;
      RECT 8.135 1.084 8.145 1.386 ;
      RECT 8.125 1.075 8.135 1.408 ;
      RECT 8.12 1.07 8.125 1.425 ;
      RECT 8.08 1.07 8.12 1.465 ;
      RECT 8.06 1.07 8.08 1.52 ;
      RECT 8.055 1.07 8.06 1.548 ;
      RECT 8.045 1.07 8.055 1.563 ;
      RECT 8.01 1.07 8.045 1.605 ;
      RECT 8.005 1.07 8.01 1.648 ;
      RECT 7.995 1.07 8.005 1.663 ;
      RECT 7.98 1.07 7.995 1.683 ;
      RECT 7.965 1.07 7.98 1.71 ;
      RECT 7.96 1.071 7.965 1.728 ;
      RECT 7.94 1.072 7.96 1.735 ;
      RECT 7.885 1.073 7.94 1.755 ;
      RECT 7.875 1.074 7.885 1.769 ;
      RECT 7.87 1.077 7.875 1.768 ;
      RECT 7.83 1.15 7.87 1.766 ;
      RECT 7.815 1.23 7.83 1.764 ;
      RECT 7.79 1.285 7.815 1.762 ;
      RECT 7.775 1.35 7.79 1.761 ;
      RECT 7.73 1.382 7.775 1.758 ;
      RECT 7.645 1.405 7.73 1.753 ;
      RECT 7.62 1.425 7.645 1.748 ;
      RECT 7.55 1.43 7.62 1.744 ;
      RECT 7.53 1.432 7.55 1.741 ;
      RECT 7.445 1.443 7.53 1.735 ;
      RECT 7.44 1.454 7.445 1.73 ;
      RECT 7.43 1.456 7.44 1.73 ;
      RECT 7.395 1.46 7.43 1.728 ;
      RECT 7.345 1.47 7.395 1.715 ;
      RECT 7.325 1.478 7.345 1.7 ;
      RECT 7.245 1.49 7.325 1.683 ;
      RECT 7.41 1.04 7.58 1.25 ;
      RECT 7.526 1.036 7.58 1.25 ;
      RECT 7.331 1.04 7.58 1.241 ;
      RECT 7.331 1.04 7.585 1.23 ;
      RECT 7.245 1.04 7.585 1.221 ;
      RECT 7.245 1.048 7.595 1.165 ;
      RECT 7.245 1.06 7.6 1.078 ;
      RECT 7.245 1.067 7.605 1.07 ;
      RECT 7.44 1.038 7.58 1.25 ;
      RECT 7.195 1.983 7.44 2.315 ;
      RECT 7.19 1.975 7.195 2.312 ;
      RECT 7.16 1.995 7.44 2.293 ;
      RECT 7.14 2.027 7.44 2.266 ;
      RECT 7.19 1.98 7.367 2.312 ;
      RECT 7.19 1.977 7.281 2.312 ;
      RECT 7.13 0.325 7.3 0.745 ;
      RECT 7.125 0.325 7.3 0.743 ;
      RECT 7.125 0.325 7.325 0.733 ;
      RECT 7.125 0.325 7.345 0.708 ;
      RECT 7.12 0.325 7.345 0.703 ;
      RECT 7.12 0.325 7.355 0.693 ;
      RECT 7.12 0.325 7.36 0.688 ;
      RECT 7.12 0.33 7.365 0.683 ;
      RECT 7.12 0.362 7.38 0.673 ;
      RECT 7.12 0.432 7.405 0.656 ;
      RECT 7.1 0.432 7.405 0.648 ;
      RECT 7.1 0.492 7.415 0.625 ;
      RECT 7.1 0.532 7.425 0.57 ;
      RECT 7.085 0.325 7.36 0.55 ;
      RECT 7.075 0.34 7.365 0.448 ;
      RECT 6.665 1.73 6.835 2.255 ;
      RECT 6.66 1.73 6.835 2.248 ;
      RECT 6.65 1.73 6.84 2.213 ;
      RECT 6.645 1.74 6.84 2.185 ;
      RECT 6.64 1.76 6.84 2.168 ;
      RECT 6.65 1.735 6.845 2.158 ;
      RECT 6.635 1.78 6.845 2.15 ;
      RECT 6.63 1.8 6.845 2.135 ;
      RECT 6.625 1.83 6.845 2.125 ;
      RECT 6.615 1.875 6.845 2.1 ;
      RECT 6.645 1.745 6.85 2.083 ;
      RECT 6.61 1.927 6.85 2.078 ;
      RECT 6.645 1.755 6.855 2.048 ;
      RECT 6.605 1.96 6.855 2.045 ;
      RECT 6.6 1.985 6.855 2.025 ;
      RECT 6.64 1.772 6.865 1.965 ;
      RECT 6.635 1.794 6.875 1.858 ;
      RECT 6.585 1.041 6.6 1.31 ;
      RECT 6.54 1.025 6.585 1.355 ;
      RECT 6.535 1.013 6.54 1.405 ;
      RECT 6.525 1.009 6.535 1.438 ;
      RECT 6.52 1.006 6.525 1.466 ;
      RECT 6.505 1.008 6.52 1.508 ;
      RECT 6.5 1.012 6.505 1.548 ;
      RECT 6.48 1.017 6.5 1.6 ;
      RECT 6.476 1.022 6.48 1.657 ;
      RECT 6.39 1.041 6.476 1.694 ;
      RECT 6.38 1.062 6.39 1.73 ;
      RECT 6.375 1.07 6.38 1.731 ;
      RECT 6.37 1.112 6.375 1.732 ;
      RECT 6.355 1.2 6.37 1.733 ;
      RECT 6.345 1.35 6.355 1.735 ;
      RECT 6.34 1.395 6.345 1.737 ;
      RECT 6.305 1.437 6.34 1.74 ;
      RECT 6.3 1.455 6.305 1.743 ;
      RECT 6.223 1.461 6.3 1.749 ;
      RECT 6.137 1.475 6.223 1.762 ;
      RECT 6.051 1.489 6.137 1.776 ;
      RECT 5.965 1.503 6.051 1.789 ;
      RECT 5.905 1.515 5.965 1.801 ;
      RECT 5.88 1.522 5.905 1.808 ;
      RECT 5.866 1.525 5.88 1.813 ;
      RECT 5.78 1.533 5.866 1.829 ;
      RECT 5.775 1.54 5.78 1.844 ;
      RECT 5.751 1.54 5.775 1.851 ;
      RECT 5.665 1.543 5.751 1.879 ;
      RECT 5.58 1.547 5.665 1.923 ;
      RECT 5.515 1.551 5.58 1.96 ;
      RECT 5.49 1.554 5.515 1.976 ;
      RECT 5.415 1.567 5.49 1.98 ;
      RECT 5.39 1.585 5.415 1.984 ;
      RECT 5.38 1.592 5.39 1.986 ;
      RECT 5.365 1.595 5.38 1.987 ;
      RECT 5.305 1.607 5.365 1.991 ;
      RECT 5.295 1.621 5.305 1.995 ;
      RECT 5.24 1.631 5.295 1.983 ;
      RECT 5.215 1.652 5.24 1.966 ;
      RECT 5.195 1.672 5.215 1.957 ;
      RECT 5.19 1.685 5.195 1.952 ;
      RECT 5.175 1.697 5.19 1.948 ;
      RECT 6.41 0.352 6.415 0.375 ;
      RECT 6.405 0.343 6.41 0.415 ;
      RECT 6.4 0.341 6.405 0.458 ;
      RECT 6.395 0.332 6.4 0.493 ;
      RECT 6.39 0.322 6.395 0.565 ;
      RECT 6.385 0.312 6.39 0.63 ;
      RECT 6.38 0.309 6.385 0.67 ;
      RECT 6.355 0.303 6.38 0.76 ;
      RECT 6.32 0.291 6.355 0.785 ;
      RECT 6.31 0.282 6.32 0.785 ;
      RECT 6.175 0.28 6.185 0.768 ;
      RECT 6.165 0.28 6.175 0.735 ;
      RECT 6.16 0.28 6.165 0.71 ;
      RECT 6.155 0.28 6.16 0.698 ;
      RECT 6.15 0.28 6.155 0.68 ;
      RECT 6.14 0.28 6.15 0.645 ;
      RECT 6.135 0.282 6.14 0.623 ;
      RECT 6.13 0.288 6.135 0.608 ;
      RECT 6.125 0.294 6.13 0.593 ;
      RECT 6.11 0.306 6.125 0.566 ;
      RECT 6.105 0.317 6.11 0.534 ;
      RECT 6.1 0.327 6.105 0.518 ;
      RECT 6.09 0.335 6.1 0.487 ;
      RECT 6.085 0.345 6.09 0.461 ;
      RECT 6.08 0.402 6.085 0.444 ;
      RECT 6.185 0.28 6.31 0.785 ;
      RECT 5.9 0.967 6.16 1.265 ;
      RECT 5.895 0.974 6.16 1.263 ;
      RECT 5.9 0.969 6.175 1.258 ;
      RECT 5.89 0.982 6.175 1.255 ;
      RECT 5.89 0.987 6.18 1.248 ;
      RECT 5.885 0.995 6.18 1.245 ;
      RECT 5.885 1.012 6.185 1.043 ;
      RECT 5.9 0.964 6.131 1.265 ;
      RECT 5.955 0.963 6.131 1.265 ;
      RECT 5.955 0.96 6.045 1.265 ;
      RECT 5.955 0.957 6.041 1.265 ;
      RECT 5.645 1.23 5.65 1.243 ;
      RECT 5.64 1.197 5.645 1.248 ;
      RECT 5.635 1.152 5.64 1.255 ;
      RECT 5.63 1.107 5.635 1.263 ;
      RECT 5.625 1.075 5.63 1.271 ;
      RECT 5.62 1.035 5.625 1.272 ;
      RECT 5.605 1.015 5.62 1.274 ;
      RECT 5.53 0.997 5.605 1.286 ;
      RECT 5.52 0.99 5.53 1.297 ;
      RECT 5.515 0.99 5.52 1.299 ;
      RECT 5.485 0.996 5.515 1.303 ;
      RECT 5.445 1.009 5.485 1.303 ;
      RECT 5.42 1.02 5.445 1.289 ;
      RECT 5.405 1.026 5.42 1.272 ;
      RECT 5.395 1.028 5.405 1.263 ;
      RECT 5.39 1.029 5.395 1.258 ;
      RECT 5.385 1.03 5.39 1.253 ;
      RECT 5.38 1.031 5.385 1.25 ;
      RECT 5.355 1.036 5.38 1.24 ;
      RECT 5.345 1.052 5.355 1.227 ;
      RECT 5.34 1.072 5.345 1.222 ;
      RECT 5.35 0.465 5.355 0.661 ;
      RECT 5.335 0.429 5.35 0.663 ;
      RECT 5.325 0.411 5.335 0.668 ;
      RECT 5.315 0.397 5.325 0.672 ;
      RECT 5.27 0.381 5.315 0.682 ;
      RECT 5.265 0.371 5.27 0.691 ;
      RECT 5.22 0.36 5.265 0.697 ;
      RECT 5.215 0.348 5.22 0.704 ;
      RECT 5.2 0.343 5.215 0.708 ;
      RECT 5.185 0.335 5.2 0.713 ;
      RECT 5.175 0.328 5.185 0.718 ;
      RECT 5.165 0.325 5.175 0.723 ;
      RECT 5.155 0.325 5.165 0.724 ;
      RECT 5.15 0.322 5.155 0.723 ;
      RECT 5.115 0.317 5.14 0.722 ;
      RECT 5.091 0.313 5.115 0.721 ;
      RECT 5.005 0.304 5.091 0.718 ;
      RECT 4.99 0.296 5.005 0.715 ;
      RECT 4.968 0.295 4.99 0.714 ;
      RECT 4.882 0.295 4.968 0.712 ;
      RECT 4.796 0.295 4.882 0.71 ;
      RECT 4.71 0.295 4.796 0.707 ;
      RECT 4.7 0.295 4.71 0.698 ;
      RECT 4.67 0.295 4.7 0.658 ;
      RECT 4.66 0.305 4.67 0.613 ;
      RECT 4.655 0.345 4.66 0.598 ;
      RECT 4.65 0.36 4.655 0.585 ;
      RECT 4.62 0.44 4.65 0.547 ;
      RECT 5.14 0.32 5.15 0.723 ;
      RECT 4.965 1.085 4.98 1.69 ;
      RECT 4.97 1.08 4.98 1.69 ;
      RECT 5.135 1.08 5.14 1.263 ;
      RECT 5.125 1.08 5.135 1.293 ;
      RECT 5.11 1.08 5.125 1.353 ;
      RECT 5.105 1.08 5.11 1.398 ;
      RECT 5.1 1.08 5.105 1.428 ;
      RECT 5.095 1.08 5.1 1.448 ;
      RECT 5.085 1.08 5.095 1.483 ;
      RECT 5.07 1.08 5.085 1.515 ;
      RECT 5.025 1.08 5.07 1.543 ;
      RECT 5.02 1.08 5.025 1.573 ;
      RECT 5.015 1.08 5.02 1.585 ;
      RECT 5.01 1.08 5.015 1.593 ;
      RECT 5 1.08 5.01 1.608 ;
      RECT 4.995 1.08 5 1.63 ;
      RECT 4.985 1.08 4.995 1.653 ;
      RECT 4.98 1.08 4.985 1.673 ;
      RECT 4.945 1.095 4.965 1.69 ;
      RECT 4.92 1.112 4.945 1.69 ;
      RECT 4.915 1.122 4.92 1.69 ;
      RECT 4.885 1.137 4.915 1.69 ;
      RECT 4.81 1.179 4.885 1.69 ;
      RECT 4.805 1.21 4.81 1.673 ;
      RECT 4.8 1.214 4.805 1.655 ;
      RECT 4.795 1.218 4.8 1.618 ;
      RECT 4.79 1.402 4.795 1.585 ;
      RECT 4.275 1.591 4.361 2.156 ;
      RECT 4.23 1.593 4.395 2.15 ;
      RECT 4.361 1.59 4.395 2.15 ;
      RECT 4.275 1.592 4.48 2.144 ;
      RECT 4.23 1.602 4.49 2.14 ;
      RECT 4.205 1.594 4.48 2.136 ;
      RECT 4.2 1.597 4.48 2.131 ;
      RECT 4.175 1.612 4.49 2.125 ;
      RECT 4.175 1.637 4.53 2.12 ;
      RECT 4.135 1.645 4.53 2.095 ;
      RECT 4.135 1.672 4.545 2.093 ;
      RECT 4.135 1.702 4.555 2.08 ;
      RECT 4.13 1.847 4.555 2.068 ;
      RECT 4.135 1.776 4.575 2.065 ;
      RECT 4.135 1.833 4.58 1.873 ;
      RECT 4.325 1.112 4.495 1.29 ;
      RECT 4.275 1.051 4.325 1.275 ;
      RECT 4.01 1.031 4.275 1.26 ;
      RECT 3.97 1.095 4.445 1.26 ;
      RECT 3.97 1.085 4.4 1.26 ;
      RECT 3.97 1.082 4.39 1.26 ;
      RECT 3.97 1.07 4.38 1.26 ;
      RECT 3.97 1.055 4.325 1.26 ;
      RECT 4.01 1.027 4.211 1.26 ;
      RECT 4.02 1.005 4.211 1.26 ;
      RECT 4.045 0.99 4.125 1.26 ;
      RECT 3.8 1.52 3.92 1.965 ;
      RECT 3.785 1.52 3.92 1.964 ;
      RECT 3.74 1.542 3.92 1.959 ;
      RECT 3.7 1.591 3.92 1.953 ;
      RECT 3.7 1.591 3.925 1.928 ;
      RECT 3.7 1.591 3.945 1.818 ;
      RECT 3.695 1.621 3.945 1.815 ;
      RECT 3.785 1.52 3.955 1.71 ;
      RECT 3.445 0.305 3.45 0.75 ;
      RECT 3.255 0.305 3.275 0.715 ;
      RECT 3.225 0.305 3.23 0.69 ;
      RECT 3.905 0.612 3.92 0.8 ;
      RECT 3.9 0.597 3.905 0.806 ;
      RECT 3.88 0.57 3.9 0.809 ;
      RECT 3.83 0.537 3.88 0.818 ;
      RECT 3.8 0.517 3.83 0.822 ;
      RECT 3.781 0.505 3.8 0.818 ;
      RECT 3.695 0.477 3.781 0.808 ;
      RECT 3.685 0.452 3.695 0.798 ;
      RECT 3.615 0.42 3.685 0.79 ;
      RECT 3.59 0.38 3.615 0.782 ;
      RECT 3.57 0.362 3.59 0.776 ;
      RECT 3.56 0.352 3.57 0.773 ;
      RECT 3.55 0.345 3.56 0.771 ;
      RECT 3.53 0.332 3.55 0.768 ;
      RECT 3.52 0.322 3.53 0.765 ;
      RECT 3.51 0.315 3.52 0.763 ;
      RECT 3.46 0.307 3.51 0.757 ;
      RECT 3.45 0.305 3.46 0.751 ;
      RECT 3.42 0.305 3.445 0.748 ;
      RECT 3.391 0.305 3.42 0.743 ;
      RECT 3.305 0.305 3.391 0.733 ;
      RECT 3.275 0.305 3.305 0.72 ;
      RECT 3.23 0.305 3.255 0.703 ;
      RECT 3.215 0.305 3.225 0.685 ;
      RECT 3.195 0.312 3.215 0.67 ;
      RECT 3.19 0.327 3.195 0.658 ;
      RECT 3.185 0.332 3.19 0.598 ;
      RECT 3.18 0.337 3.185 0.44 ;
      RECT 3.175 0.34 3.18 0.358 ;
      RECT 3.44 1.025 3.526 1.346 ;
      RECT 3.44 1.025 3.56 1.339 ;
      RECT 3.39 1.025 3.56 1.335 ;
      RECT 3.39 1.027 3.646 1.333 ;
      RECT 3.39 1.029 3.67 1.327 ;
      RECT 3.39 1.036 3.68 1.326 ;
      RECT 3.39 1.045 3.685 1.323 ;
      RECT 3.39 1.051 3.69 1.318 ;
      RECT 3.39 1.095 3.695 1.315 ;
      RECT 3.39 1.187 3.7 1.312 ;
      RECT 2.915 1.63 2.95 1.95 ;
      RECT 3.5 1.815 3.505 1.997 ;
      RECT 3.455 1.697 3.5 2.016 ;
      RECT 3.44 1.674 3.455 2.039 ;
      RECT 3.43 1.664 3.44 2.049 ;
      RECT 3.41 1.659 3.43 2.062 ;
      RECT 3.385 1.657 3.41 2.083 ;
      RECT 3.366 1.656 3.385 2.095 ;
      RECT 3.28 1.653 3.366 2.095 ;
      RECT 3.21 1.648 3.28 2.083 ;
      RECT 3.135 1.644 3.21 2.058 ;
      RECT 3.07 1.64 3.135 2.025 ;
      RECT 3 1.637 3.07 1.985 ;
      RECT 2.97 1.633 3 1.96 ;
      RECT 2.95 1.631 2.97 1.953 ;
      RECT 2.866 1.629 2.915 1.951 ;
      RECT 2.78 1.626 2.866 1.952 ;
      RECT 2.705 1.625 2.78 1.954 ;
      RECT 2.62 1.625 2.705 1.98 ;
      RECT 2.543 1.626 2.62 2.005 ;
      RECT 2.457 1.627 2.543 2.005 ;
      RECT 2.371 1.627 2.457 2.005 ;
      RECT 2.285 1.628 2.371 2.005 ;
      RECT 2.265 1.629 2.285 1.997 ;
      RECT 2.25 1.635 2.265 1.982 ;
      RECT 2.215 1.655 2.25 1.962 ;
      RECT 2.205 1.675 2.215 1.944 ;
      RECT 3.175 0.98 3.18 1.25 ;
      RECT 3.17 0.971 3.175 1.255 ;
      RECT 3.16 0.961 3.17 1.267 ;
      RECT 3.155 0.95 3.16 1.278 ;
      RECT 3.135 0.944 3.155 1.296 ;
      RECT 3.09 0.941 3.135 1.345 ;
      RECT 3.075 0.94 3.09 1.39 ;
      RECT 3.07 0.94 3.075 1.403 ;
      RECT 3.06 0.94 3.07 1.415 ;
      RECT 3.055 0.941 3.06 1.43 ;
      RECT 3.035 0.949 3.055 1.435 ;
      RECT 3.005 0.965 3.035 1.435 ;
      RECT 2.995 0.977 3 1.435 ;
      RECT 2.96 0.992 2.995 1.435 ;
      RECT 2.93 1.012 2.96 1.435 ;
      RECT 2.92 1.037 2.93 1.435 ;
      RECT 2.915 1.065 2.92 1.435 ;
      RECT 2.91 1.095 2.915 1.435 ;
      RECT 2.905 1.112 2.91 1.435 ;
      RECT 2.895 1.14 2.905 1.435 ;
      RECT 2.885 1.175 2.895 1.435 ;
      RECT 2.88 1.21 2.885 1.435 ;
      RECT 3 0.975 3.005 1.435 ;
      RECT 2.515 1.077 2.7 1.25 ;
      RECT 2.475 0.995 2.66 1.248 ;
      RECT 2.436 1 2.66 1.244 ;
      RECT 2.35 1.009 2.66 1.239 ;
      RECT 2.266 1.025 2.665 1.234 ;
      RECT 2.18 1.045 2.69 1.228 ;
      RECT 2.18 1.065 2.695 1.228 ;
      RECT 2.266 1.035 2.69 1.234 ;
      RECT 2.35 1.01 2.665 1.239 ;
      RECT 2.515 0.992 2.66 1.25 ;
      RECT 2.515 0.987 2.615 1.25 ;
      RECT 2.601 0.981 2.615 1.25 ;
      RECT 1.99 0.305 1.995 0.704 ;
      RECT 1.735 0.305 1.77 0.702 ;
      RECT 1.33 0.34 1.335 0.696 ;
      RECT 2.075 0.343 2.08 0.598 ;
      RECT 2.07 0.341 2.075 0.604 ;
      RECT 2.065 0.34 2.07 0.611 ;
      RECT 2.04 0.333 2.065 0.635 ;
      RECT 2.035 0.326 2.04 0.659 ;
      RECT 2.03 0.322 2.035 0.668 ;
      RECT 2.02 0.317 2.03 0.681 ;
      RECT 2.015 0.314 2.02 0.69 ;
      RECT 2.01 0.312 2.015 0.695 ;
      RECT 1.995 0.308 2.01 0.705 ;
      RECT 1.98 0.302 1.99 0.704 ;
      RECT 1.942 0.3 1.98 0.704 ;
      RECT 1.856 0.302 1.942 0.704 ;
      RECT 1.77 0.304 1.856 0.703 ;
      RECT 1.699 0.305 1.735 0.702 ;
      RECT 1.613 0.307 1.699 0.702 ;
      RECT 1.527 0.309 1.613 0.701 ;
      RECT 1.441 0.311 1.527 0.701 ;
      RECT 1.355 0.314 1.441 0.7 ;
      RECT 1.345 0.32 1.355 0.699 ;
      RECT 1.335 0.332 1.345 0.697 ;
      RECT 1.275 0.367 1.33 0.693 ;
      RECT 1.27 0.397 1.275 0.455 ;
      RECT 2.015 1.477 2.03 1.67 ;
      RECT 2.01 1.445 2.015 1.67 ;
      RECT 2 1.42 2.01 1.67 ;
      RECT 1.995 1.392 2 1.67 ;
      RECT 1.965 1.315 1.995 1.67 ;
      RECT 1.94 1.197 1.965 1.67 ;
      RECT 1.935 1.135 1.94 1.67 ;
      RECT 1.925 1.122 1.935 1.67 ;
      RECT 1.905 1.112 1.925 1.67 ;
      RECT 1.89 1.095 1.905 1.67 ;
      RECT 1.86 1.083 1.89 1.67 ;
      RECT 1.855 1.082 1.86 1.615 ;
      RECT 1.85 1.082 1.855 1.573 ;
      RECT 1.835 1.081 1.85 1.525 ;
      RECT 1.82 1.081 1.835 1.463 ;
      RECT 1.8 1.081 1.82 1.423 ;
      RECT 1.795 1.081 1.8 1.408 ;
      RECT 1.77 1.08 1.795 1.403 ;
      RECT 1.7 1.079 1.77 1.39 ;
      RECT 1.685 1.078 1.7 1.375 ;
      RECT 1.655 1.077 1.685 1.358 ;
      RECT 1.65 1.077 1.655 1.343 ;
      RECT 1.6 1.076 1.65 1.323 ;
      RECT 1.535 1.075 1.6 1.278 ;
      RECT 1.53 1.075 1.535 1.25 ;
      RECT 1.615 1.612 1.62 1.869 ;
      RECT 1.595 1.531 1.615 1.886 ;
      RECT 1.575 1.525 1.595 1.915 ;
      RECT 1.515 1.512 1.575 1.935 ;
      RECT 1.47 1.496 1.515 1.936 ;
      RECT 1.386 1.484 1.47 1.924 ;
      RECT 1.3 1.471 1.386 1.908 ;
      RECT 1.29 1.464 1.3 1.9 ;
      RECT 1.245 1.461 1.29 1.84 ;
      RECT 1.225 1.457 1.245 1.755 ;
      RECT 1.21 1.455 1.225 1.708 ;
      RECT 1.18 1.452 1.21 1.678 ;
      RECT 1.145 1.448 1.18 1.655 ;
      RECT 1.102 1.443 1.145 1.643 ;
      RECT 1.016 1.434 1.102 1.652 ;
      RECT 0.93 1.423 1.016 1.664 ;
      RECT 0.865 1.414 0.93 1.673 ;
      RECT 0.845 1.405 0.865 1.678 ;
      RECT 0.84 1.398 0.845 1.68 ;
      RECT 0.8 1.383 0.84 1.677 ;
      RECT 0.78 1.362 0.8 1.672 ;
      RECT 0.765 1.35 0.78 1.665 ;
      RECT 0.76 1.342 0.765 1.658 ;
      RECT 0.745 1.322 0.76 1.651 ;
      RECT 0.74 1.185 0.745 1.645 ;
      RECT 0.66 1.074 0.74 1.617 ;
      RECT 0.651 1.067 0.66 1.583 ;
      RECT 0.565 1.061 0.651 1.508 ;
      RECT 0.54 1.052 0.565 1.42 ;
      RECT 0.51 1.047 0.54 1.395 ;
      RECT 0.445 1.056 0.51 1.38 ;
      RECT 0.425 1.072 0.445 1.355 ;
      RECT 0.415 1.078 0.425 1.303 ;
      RECT 0.395 1.1 0.415 1.185 ;
      RECT 1.05 1.065 1.22 1.25 ;
      RECT 1.05 1.065 1.255 1.248 ;
      RECT 1.1 0.975 1.27 1.239 ;
      RECT 1.05 1.132 1.275 1.232 ;
      RECT 1.065 1.01 1.27 1.239 ;
      RECT 0.265 1.743 0.33 2.186 ;
      RECT 0.205 1.768 0.33 2.184 ;
      RECT 0.205 1.768 0.385 2.178 ;
      RECT 0.19 1.793 0.385 2.177 ;
      RECT 0.33 1.73 0.405 2.174 ;
      RECT 0.265 1.755 0.485 2.168 ;
      RECT 0.19 1.794 0.53 2.162 ;
      RECT 0.175 1.821 0.53 2.153 ;
      RECT 0.19 1.814 0.55 2.145 ;
      RECT 0.175 1.823 0.555 2.128 ;
      RECT 0.17 1.84 0.555 1.955 ;
      RECT 0.175 0.562 0.21 0.8 ;
      RECT 0.175 0.562 0.24 0.799 ;
      RECT 0.175 0.562 0.355 0.795 ;
      RECT 0.175 0.562 0.41 0.773 ;
      RECT 0.185 0.505 0.465 0.673 ;
      RECT 0.29 0.345 0.32 0.796 ;
      RECT 0.32 0.34 0.5 0.553 ;
      RECT 0.19 0.481 0.5 0.553 ;
      RECT 0.24 0.377 0.29 0.797 ;
      RECT 0.21 0.433 0.5 0.553 ;
  END
END scs130hd_mpr2at_8

MACRO scs130hd_mpr2ca_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130hd_mpr2ca_8 0 0 ;
  SIZE 6.9 BY 5.44 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT 4.775 1.025 5.105 1.355 ;
      RECT 4.775 1.04 5.575 1.34 ;
      RECT 4.775 2.045 5.105 2.375 ;
      RECT 4.775 2.06 5.575 2.36 ;
      RECT 4.78 1.995 5.08 2.375 ;
      RECT 4.095 4.085 4.425 4.415 ;
      RECT 4.095 4.1 4.895 4.4 ;
      RECT 4.1 4.08 4.4 4.415 ;
      RECT 4.075 1.365 4.405 1.695 ;
      RECT 3.605 1.38 4.405 1.68 ;
      RECT 4.1 1.35 4.4 1.695 ;
      RECT 3.415 3.065 3.745 3.395 ;
      RECT 3.415 3.08 4.215 3.38 ;
      RECT 3.05 4.085 3.38 4.415 ;
      RECT 2.58 4.1 3.38 4.4 ;
      RECT 2.735 0.68 3.065 1.01 ;
      RECT 2.265 0.7 2.625 1 ;
      RECT 2.625 0.695 3.065 0.995 ;
      RECT 2.345 4.78 2.645 5.195 ;
      RECT 2.375 4.765 2.705 5.095 ;
      RECT 1.905 4.78 2.705 5.08 ;
    LAYER via2 ;
      RECT 4.84 1.09 5.04 1.29 ;
      RECT 4.84 2.11 5.04 2.31 ;
      RECT 4.16 4.15 4.36 4.35 ;
      RECT 4.14 1.43 4.34 1.63 ;
      RECT 3.48 3.13 3.68 3.33 ;
      RECT 3.115 4.15 3.315 4.35 ;
      RECT 2.8 0.745 3 0.945 ;
      RECT 2.44 4.83 2.64 5.03 ;
    LAYER met2 ;
      RECT 6.5 3.07 6.76 3.39 ;
      RECT 6.56 1.03 6.7 3.39 ;
      RECT 6.5 1.03 6.76 1.35 ;
      RECT 5.48 4.09 5.74 4.41 ;
      RECT 4.86 4.18 5.74 4.32 ;
      RECT 4.86 2.025 5 4.32 ;
      RECT 4.8 2.025 5.08 2.395 ;
      RECT 4.12 4.065 4.4 4.435 ;
      RECT 4.18 2.14 4.32 4.435 ;
      RECT 4.18 2.14 4.66 2.28 ;
      RECT 4.52 0.35 4.66 2.28 ;
      RECT 4.46 0.35 4.72 0.67 ;
      RECT 3.44 3.045 3.72 3.415 ;
      RECT 3.5 0.69 3.64 3.415 ;
      RECT 3.44 0.69 3.7 1.01 ;
      RECT 3.075 4.065 3.355 4.435 ;
      RECT 3.075 4.09 3.36 4.41 ;
      RECT 4.8 1.005 5.08 1.375 ;
      RECT 4.1 1.345 4.38 1.715 ;
      RECT 2.76 0.66 3.04 1.03 ;
      RECT 2.4 4.745 2.68 5.115 ;
    LAYER via1 ;
      RECT 6.555 1.115 6.705 1.265 ;
      RECT 6.555 3.155 6.705 3.305 ;
      RECT 5.535 4.175 5.685 4.325 ;
      RECT 4.855 1.115 5.005 1.265 ;
      RECT 4.855 2.135 5.005 2.285 ;
      RECT 4.515 0.435 4.665 0.585 ;
      RECT 4.175 1.455 4.325 1.605 ;
      RECT 4.175 4.175 4.325 4.325 ;
      RECT 3.495 0.775 3.645 0.925 ;
      RECT 3.495 3.155 3.645 3.305 ;
      RECT 3.155 4.175 3.305 4.325 ;
      RECT 2.815 0.77 2.965 0.92 ;
      RECT 2.475 4.855 2.625 5.005 ;
    LAYER met1 ;
      RECT 6.47 1.06 6.79 1.32 ;
      RECT 6.195 1.12 6.79 1.26 ;
      RECT 4.09 1.4 4.41 1.66 ;
      RECT 6.065 1.415 6.355 1.645 ;
      RECT 4.09 1.46 6.355 1.6 ;
      RECT 5.45 4.12 5.77 4.38 ;
      RECT 5.45 4.18 6.045 4.32 ;
      RECT 4.77 1.06 5.09 1.32 ;
      RECT 0.03 1.075 0.32 1.305 ;
      RECT 0.03 1.12 5.09 1.26 ;
      RECT 4.86 0.78 5 1.32 ;
      RECT 4.86 0.78 5.34 0.92 ;
      RECT 5.2 0.395 5.34 0.92 ;
      RECT 5.125 0.395 5.415 0.625 ;
      RECT 4.77 2.08 5.09 2.34 ;
      RECT 4.105 2.095 4.395 2.325 ;
      RECT 1.895 2.095 2.185 2.325 ;
      RECT 1.895 2.14 5.09 2.28 ;
      RECT 3.07 4.12 3.39 4.38 ;
      RECT 4.785 4.135 5.075 4.365 ;
      RECT 2.405 4.135 2.695 4.365 ;
      RECT 2.405 4.18 3.39 4.32 ;
      RECT 4.86 3.84 5 4.365 ;
      RECT 3.16 3.84 3.3 4.38 ;
      RECT 3.16 3.84 5 3.98 ;
      RECT 2.065 0.735 2.355 0.965 ;
      RECT 2.14 0.44 2.28 0.965 ;
      RECT 4.43 0.38 4.75 0.64 ;
      RECT 4.33 0.395 4.75 0.625 ;
      RECT 2.14 0.44 4.75 0.58 ;
      RECT 3.41 0.72 3.73 0.98 ;
      RECT 3.41 0.78 4.005 0.92 ;
      RECT 2.39 4.8 2.71 5.06 ;
      RECT 1.46 4.86 3.81 5 ;
      RECT 3.67 4.135 3.81 5 ;
      RECT 1.46 4.135 1.6 5 ;
      RECT 3.595 4.135 3.885 4.365 ;
      RECT 1.385 4.135 1.675 4.365 ;
      RECT 3.41 3.1 3.73 3.36 ;
      RECT 0.705 3.115 0.995 3.345 ;
      RECT 0.705 3.16 3.73 3.3 ;
      RECT 2.735 0.68 3.065 1.01 ;
      RECT 2.73 0.715 3.065 0.975 ;
      RECT 3.08 0.735 3.195 0.965 ;
      RECT 2.73 0.73 3.08 0.96 ;
      RECT 2.73 0.78 3.21 0.92 ;
      RECT 2.615 0.78 2.625 0.92 ;
      RECT 2.625 0.775 3.195 0.915 ;
      RECT 0 -0.24 6.9 0.24 ;
      RECT 0 2.48 6.9 2.96 ;
      RECT 0 5.2 6.9 5.68 ;
      RECT 6.145 3.1 6.79 3.36 ;
      RECT 4.09 4.12 4.41 4.38 ;
    LAYER mcon ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.585 5.355 6.755 5.525 ;
      RECT 6.545 1.105 6.715 1.275 ;
      RECT 6.205 3.145 6.375 3.315 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 1.445 6.295 1.615 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.125 5.355 6.295 5.525 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.665 5.355 5.835 5.525 ;
      RECT 5.525 4.165 5.695 4.335 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.205 5.355 5.375 5.525 ;
      RECT 5.185 0.425 5.355 0.595 ;
      RECT 4.845 4.165 5.015 4.335 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.745 5.355 4.915 5.525 ;
      RECT 4.39 0.425 4.56 0.595 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.285 5.355 4.455 5.525 ;
      RECT 4.165 2.125 4.335 2.295 ;
      RECT 4.165 4.165 4.335 4.335 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 3.825 5.355 3.995 5.525 ;
      RECT 3.655 4.165 3.825 4.335 ;
      RECT 3.485 0.765 3.655 0.935 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.365 5.355 3.535 5.525 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.905 5.355 3.075 5.525 ;
      RECT 2.465 4.165 2.635 4.335 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.445 5.355 2.615 5.525 ;
      RECT 2.125 0.765 2.295 0.935 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 1.985 5.355 2.155 5.525 ;
      RECT 1.955 2.125 2.125 2.295 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.525 5.355 1.695 5.525 ;
      RECT 1.445 4.165 1.615 4.335 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.065 5.355 1.235 5.525 ;
      RECT 0.765 3.145 0.935 3.315 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 0.09 1.105 0.26 1.275 ;
    LAYER li ;
      RECT 0.085 -0.085 0.345 0.905 ;
      RECT 6.535 -0.085 6.805 0.895 ;
      RECT 5.625 -0.085 5.865 0.895 ;
      RECT 4.755 -0.085 5.005 0.625 ;
      RECT 2.375 -0.085 2.705 0.545 ;
      RECT 0 -0.085 6.9 0.085 ;
      RECT 3.355 1.98 3.62 3.585 ;
      RECT 1.195 2.13 1.525 3.525 ;
      RECT 2.195 2.635 2.475 3.475 ;
      RECT 4.17 2.635 4.545 3.185 ;
      RECT 0 2.635 6.9 2.805 ;
      RECT 6.475 1.495 6.805 2.805 ;
      RECT 4.735 2.09 4.99 2.805 ;
      RECT 3.305 1.98 3.91 2.805 ;
      RECT 2.435 2.09 2.65 2.805 ;
      RECT 1.005 2.13 1.62 2.805 ;
      RECT 1.425 1.765 1.62 2.805 ;
      RECT 0.085 2.125 0.345 2.805 ;
      RECT 3.735 1.71 3.92 2.08 ;
      RECT 3.735 1.71 4.065 1.955 ;
      RECT 1.425 1.765 1.755 1.955 ;
      RECT 0 5.355 6.9 5.525 ;
      RECT 5.435 4.845 5.885 5.525 ;
      RECT 3.345 4.955 3.675 5.525 ;
      RECT 1.275 4.895 1.525 5.525 ;
      RECT 3.855 4.935 5.16 5.185 ;
      RECT 3.855 4.615 4.035 5.185 ;
      RECT 3.305 4.615 4.035 4.785 ;
      RECT 3.305 3.775 3.475 4.785 ;
      RECT 4.14 3.815 5.885 3.995 ;
      RECT 5.555 2.975 5.885 3.995 ;
      RECT 3.305 3.775 4.365 3.945 ;
      RECT 5.555 3.145 6.375 3.315 ;
      RECT 4.715 2.975 5.045 3.185 ;
      RECT 4.715 2.975 5.885 3.145 ;
      RECT 5.615 1.495 5.945 2.45 ;
      RECT 5.615 1.495 6.295 1.665 ;
      RECT 6.125 0.255 6.295 1.665 ;
      RECT 6.035 0.255 6.365 0.895 ;
      RECT 5.16 1.765 5.435 2.465 ;
      RECT 5.265 0.255 5.435 2.465 ;
      RECT 5.605 1.075 5.955 1.325 ;
      RECT 5.265 1.105 5.955 1.275 ;
      RECT 5.175 0.255 5.435 0.735 ;
      RECT 4.505 3.405 5.385 3.645 ;
      RECT 5.155 3.315 5.385 3.645 ;
      RECT 3.855 3.405 5.385 3.605 ;
      RECT 4.77 3.355 5.385 3.645 ;
      RECT 3.855 3.275 4.025 3.605 ;
      RECT 4.74 4.165 4.99 4.765 ;
      RECT 4.74 4.165 5.215 4.365 ;
      RECT 4.235 1.385 4.99 1.885 ;
      RECT 3.305 1.19 3.565 1.81 ;
      RECT 4.22 1.33 4.235 1.635 ;
      RECT 4.205 1.315 4.225 1.6 ;
      RECT 4.865 0.99 5.095 1.59 ;
      RECT 4.18 1.26 4.2 1.575 ;
      RECT 4.16 1.385 5.095 1.56 ;
      RECT 4.135 1.385 5.095 1.55 ;
      RECT 4.065 1.385 5.095 1.54 ;
      RECT 4.045 1.385 5.095 1.51 ;
      RECT 4.025 0.295 4.195 1.48 ;
      RECT 3.995 1.385 5.095 1.45 ;
      RECT 3.96 1.385 5.095 1.425 ;
      RECT 3.93 1.38 4.32 1.39 ;
      RECT 3.93 1.37 4.295 1.39 ;
      RECT 3.93 1.365 4.28 1.39 ;
      RECT 3.93 1.355 4.265 1.39 ;
      RECT 3.305 1.19 4.195 1.36 ;
      RECT 3.305 1.345 4.255 1.36 ;
      RECT 3.305 1.34 4.245 1.36 ;
      RECT 4.2 1.285 4.21 1.59 ;
      RECT 3.305 1.32 4.23 1.36 ;
      RECT 3.305 1.3 4.215 1.36 ;
      RECT 3.305 0.295 4.195 0.465 ;
      RECT 4.365 0.79 4.695 1.215 ;
      RECT 4.365 0.305 4.585 1.215 ;
      RECT 4.28 4.165 4.49 4.765 ;
      RECT 4.14 4.165 4.49 4.365 ;
      RECT 2.86 1.765 3.135 2.465 ;
      RECT 3.08 0.255 3.135 2.465 ;
      RECT 2.965 1.06 3.135 2.465 ;
      RECT 2.965 0.255 3.135 1.055 ;
      RECT 2.875 0.255 3.135 0.73 ;
      RECT 1.005 1.425 1.255 1.96 ;
      RECT 1.975 1.425 2.69 1.89 ;
      RECT 1.005 1.425 2.795 1.595 ;
      RECT 2.565 1.06 2.795 1.595 ;
      RECT 1.56 0.305 1.815 1.595 ;
      RECT 2.565 0.995 2.625 1.89 ;
      RECT 2.625 0.99 2.795 1.055 ;
      RECT 1.025 0.305 1.815 0.57 ;
      RECT 1.985 4.115 2.66 4.365 ;
      RECT 2.395 3.755 2.66 4.365 ;
      RECT 2.145 4.535 2.475 5.085 ;
      RECT 1.085 4.535 2.475 4.725 ;
      RECT 1.085 3.695 1.255 4.725 ;
      RECT 0.965 4.115 1.255 4.445 ;
      RECT 1.085 3.695 2.025 3.865 ;
      RECT 1.725 3.145 2.025 3.865 ;
      RECT 1.985 0.725 2.395 1.245 ;
      RECT 1.985 0.305 2.185 1.245 ;
      RECT 0.595 0.485 0.765 2.465 ;
      RECT 0.595 0.995 1.39 1.245 ;
      RECT 0.595 0.485 0.845 1.245 ;
      RECT 0.515 0.485 0.845 0.905 ;
      RECT 0.545 4.895 1.105 5.185 ;
      RECT 0.545 2.975 0.795 5.185 ;
      RECT 0.545 2.975 1.005 3.525 ;
      RECT 6.465 1.075 6.815 1.325 ;
      RECT 5.405 4.165 5.855 4.675 ;
      RECT 4.085 2.125 4.565 2.465 ;
      RECT 3.645 4.115 3.97 4.445 ;
      RECT 3.305 0.635 3.855 1.02 ;
      RECT 1.79 2.125 2.265 2.465 ;
      RECT 1.425 4.115 1.765 4.365 ;
      RECT 0.085 1.075 0.425 1.955 ;
  END
END scs130hd_mpr2ca_8

MACRO scs130hd_mpr2ct_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130hd_mpr2ct_8 0 0 ;
  SIZE 7.36 BY 5.44 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT 5.115 4.08 5.445 4.41 ;
      RECT 5.115 4.095 5.915 4.395 ;
      RECT 5.17 4.055 5.47 4.395 ;
      RECT 4.765 2.045 5.095 2.375 ;
      RECT 4.765 2.06 5.565 2.36 ;
      RECT 4.78 2.015 5.08 2.375 ;
      RECT 4.425 1.365 4.755 1.695 ;
      RECT 4.425 1.38 5.225 1.68 ;
      RECT 4.51 1.355 4.81 1.68 ;
      RECT 4.075 4.08 4.405 4.41 ;
      RECT 3.605 4.095 4.405 4.395 ;
      RECT 4.1 4.035 4.4 4.41 ;
      RECT 3.745 2.445 4.075 2.775 ;
      RECT 1.705 2.445 2.035 2.775 ;
      RECT 1.705 2.46 4.075 2.76 ;
      RECT 3.395 1.705 3.725 2.035 ;
      RECT 2.935 1.72 3.735 2.02 ;
      RECT 3.065 0.515 3.395 0.845 ;
      RECT 2.595 0.53 3.395 0.83 ;
      RECT 3.055 0.525 3.395 0.83 ;
      RECT 3.065 4.77 3.395 5.1 ;
      RECT 2.595 4.785 3.395 5.085 ;
      RECT 2.975 4.745 3.275 5.085 ;
      RECT 2.385 4.08 2.715 4.41 ;
      RECT 1.915 4.095 2.715 4.395 ;
    LAYER via2 ;
      RECT 5.18 4.145 5.38 4.345 ;
      RECT 4.83 2.11 5.03 2.31 ;
      RECT 4.49 1.43 4.69 1.63 ;
      RECT 4.14 4.145 4.34 4.345 ;
      RECT 3.81 2.51 4.01 2.71 ;
      RECT 3.46 1.77 3.66 1.97 ;
      RECT 3.13 0.58 3.33 0.78 ;
      RECT 3.13 4.835 3.33 5.035 ;
      RECT 2.45 4.145 2.65 4.345 ;
      RECT 1.77 2.51 1.97 2.71 ;
    LAYER met2 ;
      RECT 6.16 4.77 6.42 5.09 ;
      RECT 6.22 1.03 6.36 5.09 ;
      RECT 6.16 1.03 6.42 1.35 ;
      RECT 5.48 3.07 5.74 3.39 ;
      RECT 5.54 2.05 5.68 3.39 ;
      RECT 5.48 2.05 5.74 2.37 ;
      RECT 4.46 4.77 4.72 5.09 ;
      RECT 4.52 3.5 4.66 5.09 ;
      RECT 3.84 3.5 4.66 3.64 ;
      RECT 3.84 1.03 3.98 3.64 ;
      RECT 3.77 2.425 4.05 2.795 ;
      RECT 3.78 1.03 4.04 1.35 ;
      RECT 1.73 2.425 2.01 2.795 ;
      RECT 1.8 0.69 1.94 2.795 ;
      RECT 1.74 0.69 2 1.01 ;
      RECT 1.06 3.07 1.32 3.39 ;
      RECT 1.12 1.03 1.26 3.39 ;
      RECT 1.06 1.03 1.32 1.35 ;
      RECT 5.14 4.06 5.42 4.43 ;
      RECT 4.79 2.025 5.07 2.395 ;
      RECT 4.45 1.345 4.73 1.715 ;
      RECT 4.1 4.06 4.38 4.43 ;
      RECT 3.42 1.685 3.7 2.055 ;
      RECT 3.09 0.495 3.37 0.865 ;
      RECT 3.09 4.75 3.37 5.12 ;
      RECT 2.41 4.06 2.69 4.43 ;
    LAYER via1 ;
      RECT 6.215 1.115 6.365 1.265 ;
      RECT 6.215 4.855 6.365 5.005 ;
      RECT 5.535 2.135 5.685 2.285 ;
      RECT 5.535 3.155 5.685 3.305 ;
      RECT 5.195 4.175 5.345 4.325 ;
      RECT 4.855 2.135 5.005 2.285 ;
      RECT 4.515 1.455 4.665 1.605 ;
      RECT 4.515 4.855 4.665 5.005 ;
      RECT 4.165 4.175 4.315 4.325 ;
      RECT 3.835 1.115 3.985 1.265 ;
      RECT 3.495 1.795 3.645 1.945 ;
      RECT 3.155 0.605 3.305 0.755 ;
      RECT 3.155 4.855 3.305 5.005 ;
      RECT 2.475 4.175 2.625 4.325 ;
      RECT 1.795 0.775 1.945 0.925 ;
      RECT 1.115 1.115 1.265 1.265 ;
      RECT 1.115 3.155 1.265 3.305 ;
    LAYER met1 ;
      RECT 5.45 2.08 5.77 2.34 ;
      RECT 6.485 2.095 6.775 2.325 ;
      RECT 5.45 2.14 6.775 2.28 ;
      RECT 5.11 4.12 5.43 4.38 ;
      RECT 6.485 4.135 6.775 4.365 ;
      RECT 6.56 3.84 6.7 4.365 ;
      RECT 5.2 3.84 5.34 4.38 ;
      RECT 5.2 3.84 6.7 3.98 ;
      RECT 6.13 1.06 6.45 1.32 ;
      RECT 5.855 1.12 6.45 1.26 ;
      RECT 3.07 4.8 3.39 5.06 ;
      RECT 2.065 4.815 2.355 5.045 ;
      RECT 2.065 4.86 3.98 5 ;
      RECT 3.84 4.52 3.98 5 ;
      RECT 3.84 4.52 5.85 4.66 ;
      RECT 5.71 4.135 5.85 4.66 ;
      RECT 5.635 4.135 5.925 4.365 ;
      RECT 5.45 3.1 5.77 3.36 ;
      RECT 3.305 3.115 3.595 3.345 ;
      RECT 3.305 3.16 5.77 3.3 ;
      RECT 4.77 2.08 5.09 2.34 ;
      RECT 2.405 2.095 2.695 2.325 ;
      RECT 2.405 2.14 5.09 2.28 ;
      RECT 4.43 4.8 4.75 5.06 ;
      RECT 4.43 4.86 5.025 5 ;
      RECT 4.43 1.4 4.75 1.66 ;
      RECT 4.155 1.46 4.75 1.6 ;
      RECT 3.75 1.06 4.07 1.32 ;
      RECT 3.475 1.12 4.07 1.26 ;
      RECT 3.41 1.74 3.73 2 ;
      RECT 0.535 1.755 0.825 1.985 ;
      RECT 0.535 1.8 3.73 1.94 ;
      RECT 2.99 1.08 3.13 1.94 ;
      RECT 2.915 1.08 3.205 1.31 ;
      RECT 3.07 0.55 3.39 0.81 ;
      RECT 3.07 0.565 3.575 0.795 ;
      RECT 2.98 0.61 3.575 0.75 ;
      RECT 2.39 4.12 2.71 4.38 ;
      RECT 0.025 4.135 0.315 4.365 ;
      RECT 0.025 4.18 2.71 4.32 ;
      RECT 2.405 1.08 2.695 1.31 ;
      RECT 1.8 1.125 2.695 1.265 ;
      RECT 1.8 0.72 1.94 1.265 ;
      RECT 1.71 0.72 2.03 0.98 ;
      RECT 1.03 1.06 1.35 1.32 ;
      RECT 0.755 1.12 1.35 1.26 ;
      RECT 1.03 3.1 1.35 3.36 ;
      RECT 0.755 3.16 1.35 3.3 ;
      RECT 0 -0.24 7.36 0.24 ;
      RECT 0 2.48 7.36 2.96 ;
      RECT 0 5.2 7.36 5.68 ;
      RECT 5.805 4.8 6.45 5.06 ;
      RECT 3.755 4.12 4.4 4.38 ;
    LAYER mcon ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 7.045 5.355 7.215 5.525 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.585 5.355 6.755 5.525 ;
      RECT 6.545 2.125 6.715 2.295 ;
      RECT 6.545 4.165 6.715 4.335 ;
      RECT 6.205 1.105 6.375 1.275 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.125 5.355 6.295 5.525 ;
      RECT 5.865 4.845 6.035 5.015 ;
      RECT 5.695 4.165 5.865 4.335 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.665 5.355 5.835 5.525 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 5.205 5.355 5.375 5.525 ;
      RECT 5.185 4.165 5.355 4.335 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.745 5.355 4.915 5.525 ;
      RECT 4.505 1.445 4.675 1.615 ;
      RECT 4.505 4.845 4.675 5.015 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.285 5.355 4.455 5.525 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 1.105 3.995 1.275 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 3.825 5.355 3.995 5.525 ;
      RECT 3.815 4.165 3.985 4.335 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.365 3.145 3.535 3.315 ;
      RECT 3.365 5.355 3.535 5.525 ;
      RECT 3.345 0.595 3.515 0.765 ;
      RECT 2.975 1.11 3.145 1.28 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.905 5.355 3.075 5.525 ;
      RECT 2.465 1.11 2.635 1.28 ;
      RECT 2.465 2.125 2.635 2.295 ;
      RECT 2.465 4.165 2.635 4.335 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.445 5.355 2.615 5.525 ;
      RECT 2.125 4.845 2.295 5.015 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 1.985 5.355 2.155 5.525 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.525 5.355 1.695 5.525 ;
      RECT 1.105 1.105 1.275 1.275 ;
      RECT 1.105 3.145 1.275 3.315 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.065 5.355 1.235 5.525 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.595 1.785 0.765 1.955 ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 0.085 4.165 0.255 4.335 ;
    LAYER li ;
      RECT 4.225 -0.085 4.515 0.92 ;
      RECT 1.025 -0.085 1.255 0.905 ;
      RECT 0.145 -0.085 0.355 0.905 ;
      RECT 3.775 -0.085 4.045 0.895 ;
      RECT 2.865 -0.085 3.105 0.895 ;
      RECT 2.415 -0.085 2.655 0.895 ;
      RECT 1.475 -0.085 1.745 0.895 ;
      RECT 6.895 -0.085 7.225 0.475 ;
      RECT 6.055 -0.085 6.385 0.475 ;
      RECT 0 -0.085 7.36 0.085 ;
      RECT 6.535 2.635 6.815 3.945 ;
      RECT 5.605 2.635 5.865 3.945 ;
      RECT 5.155 2.635 5.435 3.945 ;
      RECT 4.225 2.635 4.485 3.945 ;
      RECT 3.795 2.635 4.055 3.945 ;
      RECT 2.845 2.635 3.125 3.945 ;
      RECT 1.495 1.495 1.755 3.945 ;
      RECT 0.545 2.635 0.825 3.945 ;
      RECT 0 2.635 7.36 2.805 ;
      RECT 6.135 1.785 6.305 2.805 ;
      RECT 5.295 2.125 5.465 2.805 ;
      RECT 3.715 1.495 4.045 2.805 ;
      RECT 1.475 1.495 1.805 2.805 ;
      RECT 1.025 1.495 1.255 2.805 ;
      RECT 0.145 1.495 0.355 2.805 ;
      RECT 0 5.355 7.36 5.525 ;
      RECT 6.505 4.555 6.815 5.525 ;
      RECT 5.125 4.555 5.435 5.525 ;
      RECT 2.845 4.555 3.155 5.525 ;
      RECT 0.545 4.555 0.855 5.525 ;
      RECT 6.895 1.785 7.275 2.465 ;
      RECT 7.105 0.655 7.275 2.465 ;
      RECT 5.025 0.655 5.255 1.325 ;
      RECT 5.025 0.655 7.275 0.825 ;
      RECT 6.555 0.335 6.725 0.825 ;
      RECT 6.545 1.445 6.715 2.295 ;
      RECT 5.63 1.445 6.935 1.615 ;
      RECT 6.69 0.995 6.935 1.615 ;
      RECT 5.63 1.075 5.8 1.615 ;
      RECT 5.425 1.075 5.8 1.245 ;
      RECT 5.605 4.555 6.3 5.185 ;
      RECT 6.13 2.975 6.3 5.185 ;
      RECT 6.035 2.975 6.365 3.955 ;
      RECT 5.635 1.785 5.965 2.465 ;
      RECT 4.725 1.785 5.125 2.465 ;
      RECT 4.725 1.785 5.965 1.955 ;
      RECT 4.225 1.365 4.545 2.465 ;
      RECT 4.225 1.365 4.675 1.615 ;
      RECT 4.225 1.365 4.855 1.535 ;
      RECT 4.685 0.315 4.855 1.535 ;
      RECT 4.685 0.315 5.64 0.485 ;
      RECT 4.225 4.555 4.92 5.185 ;
      RECT 4.75 2.975 4.92 5.185 ;
      RECT 4.655 2.975 4.985 3.955 ;
      RECT 4.245 4.115 4.58 4.365 ;
      RECT 3.7 4.115 4.035 4.365 ;
      RECT 3.7 4.165 4.58 4.335 ;
      RECT 3.36 4.555 4.055 5.185 ;
      RECT 3.36 2.975 3.53 5.185 ;
      RECT 3.295 2.975 3.625 3.955 ;
      RECT 2.855 1.495 3.185 2.45 ;
      RECT 2.855 1.495 3.535 1.665 ;
      RECT 3.365 0.255 3.535 1.665 ;
      RECT 3.275 0.255 3.605 0.895 ;
      RECT 2.855 4.115 3.19 4.385 ;
      RECT 2.465 4.165 3.19 4.335 ;
      RECT 2.335 1.495 2.665 2.45 ;
      RECT 1.985 1.495 2.665 1.665 ;
      RECT 1.985 0.255 2.155 1.665 ;
      RECT 1.915 0.255 2.245 0.895 ;
      RECT 2.125 4.165 2.295 5.015 ;
      RECT 1.4 4.115 1.735 4.365 ;
      RECT 1.4 4.165 2.295 4.335 ;
      RECT 1.465 1.075 1.815 1.325 ;
      RECT 0.945 1.075 1.275 1.325 ;
      RECT 0.945 1.105 1.815 1.275 ;
      RECT 1.06 4.555 1.755 5.185 ;
      RECT 1.06 2.975 1.23 5.185 ;
      RECT 0.995 2.975 1.325 3.955 ;
      RECT 0.555 4.115 0.89 4.385 ;
      RECT 0.085 4.165 0.89 4.335 ;
      RECT 0.525 1.485 0.855 2.465 ;
      RECT 0.525 0.255 0.775 2.465 ;
      RECT 0.525 0.255 0.855 0.885 ;
      RECT 6.47 4.115 6.805 4.385 ;
      RECT 5.97 1.075 6.52 1.275 ;
      RECT 5.625 4.115 5.96 4.365 ;
      RECT 5.09 4.115 5.425 4.385 ;
      RECT 3.705 1.075 4.055 1.325 ;
      RECT 2.845 1.075 3.195 1.325 ;
      RECT 2.325 1.075 2.675 1.325 ;
  END
END scs130hd_mpr2ct_8

MACRO scs130hd_mpr2ea_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130hd_mpr2ea_8 0 0 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT 4.87 2.035 5.2 2.365 ;
      RECT 3.665 2.05 5.2 2.35 ;
      RECT 3.665 0.93 3.965 2.35 ;
      RECT 3.41 0.915 3.74 1.245 ;
      RECT 8.89 1.475 9.22 2.205 ;
      RECT 8.41 0.35 8.74 1.08 ;
      RECT 6.81 1.075 7.14 1.805 ;
      RECT 5.25 0.515 5.58 1.245 ;
      RECT 4.37 0.515 4.7 1.245 ;
      RECT 2.69 0.915 3.02 1.645 ;
      RECT 1.69 0.355 2.02 1.085 ;
      RECT 0.25 1.075 0.58 1.805 ;
    LAYER via2 ;
      RECT 8.955 1.54 9.155 1.74 ;
      RECT 8.475 0.815 8.675 1.015 ;
      RECT 6.875 1.54 7.075 1.74 ;
      RECT 5.315 0.98 5.515 1.18 ;
      RECT 4.935 2.1 5.135 2.3 ;
      RECT 4.435 0.98 4.635 1.18 ;
      RECT 3.475 0.98 3.675 1.18 ;
      RECT 2.755 0.98 2.955 1.18 ;
      RECT 1.755 0.42 1.955 0.62 ;
      RECT 0.315 1.54 0.515 1.74 ;
    LAYER met2 ;
      RECT 6.955 0.895 7.235 1.265 ;
      RECT 5.885 0.92 6.145 1.24 ;
      RECT 8.435 0.73 8.715 1.1 ;
      RECT 9.045 0.64 9.305 0.96 ;
      RECT 5.945 0.08 6.085 1.24 ;
      RECT 7.025 0.08 7.165 1.265 ;
      RECT 8.145 0.73 9.305 0.87 ;
      RECT 8.145 0.08 8.285 0.87 ;
      RECT 5.945 0.08 8.285 0.22 ;
      RECT 8.915 1.455 9.195 1.825 ;
      RECT 8.925 1.2 9.185 1.825 ;
      RECT 5.975 2.22 8.15 2.385 ;
      RECT 8.005 1.1 8.15 2.385 ;
      RECT 4.895 2.015 5.175 2.385 ;
      RECT 4.895 2.13 6.115 2.27 ;
      RECT 7.725 1.1 8.15 1.24 ;
      RECT 7.725 0.92 7.985 1.24 ;
      RECT 1.065 2.5 4.725 2.64 ;
      RECT 4.585 1.685 4.725 2.64 ;
      RECT 1.065 1.57 1.205 2.64 ;
      RECT 7.605 1.76 7.865 2.08 ;
      RECT 4.585 1.685 7.115 1.825 ;
      RECT 6.835 1.455 7.115 1.825 ;
      RECT 1.065 1.57 1.515 1.825 ;
      RECT 1.235 1.455 1.515 1.825 ;
      RECT 7.605 1.57 7.805 2.08 ;
      RECT 6.835 1.57 7.805 1.71 ;
      RECT 7.405 0.36 7.545 1.71 ;
      RECT 7.345 0.36 7.605 0.68 ;
      RECT 1.245 0.92 1.505 1.24 ;
      RECT 1.245 1.01 2.285 1.15 ;
      RECT 2.145 0.22 2.285 1.15 ;
      RECT 4.905 0.36 5.165 0.68 ;
      RECT 2.145 0.22 5.105 0.36 ;
      RECT 4.285 1.2 4.545 1.52 ;
      RECT 4.285 1.2 4.605 1.43 ;
      RECT 4.395 0.895 4.675 1.265 ;
      RECT 3.985 1.76 4.305 2.08 ;
      RECT 3.985 0.64 4.125 2.08 ;
      RECT 3.925 0.64 4.185 0.96 ;
      RECT 1.485 2.04 1.745 2.36 ;
      RECT 1.485 2.13 3.165 2.27 ;
      RECT 3.025 1.85 3.165 2.27 ;
      RECT 3.025 1.85 3.465 2.08 ;
      RECT 3.205 1.76 3.465 2.08 ;
      RECT 2.525 0.92 2.925 1.43 ;
      RECT 2.715 0.895 2.995 1.265 ;
      RECT 2.465 0.92 2.995 1.24 ;
      RECT 5.275 0.895 5.555 1.265 ;
      RECT 3.435 0.895 3.715 1.265 ;
      RECT 1.715 0.335 1.995 0.705 ;
      RECT 0.275 1.455 0.555 1.825 ;
    LAYER via1 ;
      RECT 9.1 0.725 9.25 0.875 ;
      RECT 8.98 1.285 9.13 1.435 ;
      RECT 7.78 1.005 7.93 1.155 ;
      RECT 7.66 1.845 7.81 1.995 ;
      RECT 7.4 0.445 7.55 0.595 ;
      RECT 5.94 1.005 6.09 1.155 ;
      RECT 5.34 1.005 5.49 1.155 ;
      RECT 4.96 0.445 5.11 0.595 ;
      RECT 4.34 1.285 4.49 1.435 ;
      RECT 4.1 1.845 4.25 1.995 ;
      RECT 3.98 0.725 4.13 0.875 ;
      RECT 3.5 1.005 3.65 1.155 ;
      RECT 3.26 1.845 3.41 1.995 ;
      RECT 2.52 1.005 2.67 1.155 ;
      RECT 1.78 0.445 1.93 0.595 ;
      RECT 1.54 2.125 1.69 2.275 ;
      RECT 1.3 1.005 1.45 1.155 ;
      RECT 1.3 1.565 1.45 1.715 ;
      RECT 0.34 1.565 0.49 1.715 ;
    LAYER met1 ;
      RECT 8.31 0.965 8.6 1.195 ;
      RECT 8.31 0.965 8.765 1.15 ;
      RECT 8.625 0.87 9.245 1.01 ;
      RECT 9.015 0.67 9.335 0.93 ;
      RECT 7.405 1.43 9.005 1.57 ;
      RECT 8.895 1.23 9.215 1.49 ;
      RECT 8.895 1.245 9.32 1.475 ;
      RECT 8.865 1.29 9.32 1.475 ;
      RECT 7.07 1.29 7.545 1.475 ;
      RECT 7.07 1.245 7.36 1.475 ;
      RECT 7.695 0.95 8.015 1.21 ;
      RECT 7.695 0.95 8.16 1.195 ;
      RECT 8.02 0.57 8.16 1.195 ;
      RECT 8.02 0.57 8.285 0.71 ;
      RECT 8.55 0.405 8.84 0.635 ;
      RECT 8.145 0.45 8.84 0.59 ;
      RECT 7.59 1.79 7.88 2.315 ;
      RECT 7.575 1.79 7.895 2.05 ;
      RECT 7.315 0.39 7.635 0.65 ;
      RECT 7.315 0.405 7.88 0.635 ;
      RECT 6.59 2.085 6.88 2.315 ;
      RECT 6.785 0.73 6.925 2.27 ;
      RECT 6.83 0.685 7.12 0.915 ;
      RECT 6.425 0.73 7.12 0.87 ;
      RECT 6.425 0.57 6.565 0.87 ;
      RECT 4.965 0.57 6.565 0.71 ;
      RECT 4.875 0.39 5.195 0.65 ;
      RECT 4.875 0.405 5.44 0.65 ;
      RECT 3.985 1.43 6.565 1.57 ;
      RECT 6.35 1.245 6.64 1.475 ;
      RECT 3.91 1.245 4.575 1.475 ;
      RECT 4.255 1.23 4.575 1.57 ;
      RECT 5.255 0.95 5.575 1.21 ;
      RECT 5.255 0.965 5.68 1.195 ;
      RECT 3.895 0.67 4.215 0.93 ;
      RECT 4.39 0.685 4.68 0.915 ;
      RECT 3.895 0.73 4.68 0.87 ;
      RECT 4.015 1.79 4.335 2.05 ;
      RECT 3.175 1.79 3.495 2.05 ;
      RECT 4.015 1.805 4.44 2.035 ;
      RECT 3.175 1.85 4.44 1.99 ;
      RECT 2.71 1.525 3 1.755 ;
      RECT 2.785 0.45 2.925 1.755 ;
      RECT 2.435 0.95 2.925 1.21 ;
      RECT 2.19 0.965 2.925 1.195 ;
      RECT 3.19 0.405 3.48 0.635 ;
      RECT 2.785 0.45 3.48 0.59 ;
      RECT 1.95 1.805 2.24 2.035 ;
      RECT 1.95 1.805 2.405 1.99 ;
      RECT 2.265 1.43 2.405 1.99 ;
      RECT 1.905 1.43 2.405 1.57 ;
      RECT 1.905 0.45 2.045 1.57 ;
      RECT 1.695 0.39 2.015 0.65 ;
      RECT 1.455 2.07 1.775 2.33 ;
      RECT 0.75 2.085 1.04 2.315 ;
      RECT 0.75 2.13 1.775 2.27 ;
      RECT 0.825 2.08 1.085 2.27 ;
      RECT 1.215 0.95 1.535 1.21 ;
      RECT 1.215 0.965 1.76 1.195 ;
      RECT 1.215 1.51 1.535 1.77 ;
      RECT 1.215 1.525 1.76 1.755 ;
      RECT 0.255 1.51 0.575 1.77 ;
      RECT 0.345 0.45 0.485 1.77 ;
      RECT 0.75 0.405 1.04 0.635 ;
      RECT 0.345 0.45 1.04 0.59 ;
      RECT 0 -0.24 9.66 0.24 ;
      RECT 0 2.48 9.66 2.96 ;
      RECT 5.855 0.95 6.175 1.21 ;
      RECT 3.415 0.95 3.735 1.21 ;
    LAYER mcon ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.09 1.275 9.26 1.445 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 8.61 0.435 8.78 0.605 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.37 0.995 8.54 1.165 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 7.89 0.995 8.06 1.165 ;
      RECT 7.65 0.435 7.82 0.605 ;
      RECT 7.65 2.115 7.82 2.285 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.13 1.275 7.3 1.445 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 6.89 0.715 7.06 0.885 ;
      RECT 6.65 2.115 6.82 2.285 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.41 1.275 6.58 1.445 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 5.93 0.995 6.1 1.165 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.45 0.995 5.62 1.165 ;
      RECT 5.21 0.435 5.38 0.605 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.45 0.715 4.62 0.885 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.21 1.835 4.38 2.005 ;
      RECT 3.97 1.275 4.14 1.445 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 3.49 0.995 3.66 1.165 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.25 0.435 3.42 0.605 ;
      RECT 3.25 1.835 3.42 2.005 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.77 1.555 2.94 1.725 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.25 0.995 2.42 1.165 ;
      RECT 2.01 1.835 2.18 2.005 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 1.77 0.435 1.94 0.605 ;
      RECT 1.53 0.995 1.7 1.165 ;
      RECT 1.53 1.555 1.7 1.725 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 0.81 0.435 0.98 0.605 ;
      RECT 0.81 2.115 0.98 2.285 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.33 1.555 0.5 1.725 ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
    LAYER li ;
      RECT 8.13 -0.085 8.3 0.585 ;
      RECT 6.17 -0.085 6.34 0.585 ;
      RECT 3.73 -0.085 3.9 0.585 ;
      RECT 2.77 -0.085 2.94 0.585 ;
      RECT 2.25 -0.085 2.42 0.585 ;
      RECT 1.29 -0.085 1.46 0.585 ;
      RECT 0.33 -0.085 0.5 0.585 ;
      RECT 0 -0.085 9.66 0.085 ;
      RECT 0 2.635 9.66 2.805 ;
      RECT 9.09 2.135 9.26 2.805 ;
      RECT 8.13 2.135 8.3 2.805 ;
      RECT 5.69 2.135 5.86 2.805 ;
      RECT 4.69 2.135 4.86 2.805 ;
      RECT 3.73 2.135 3.9 2.805 ;
      RECT 1.29 2.135 1.46 2.805 ;
      RECT 8.61 0.335 8.78 0.605 ;
      RECT 8.61 0.335 9.34 0.505 ;
      RECT 9.09 1.075 9.26 1.445 ;
      RECT 8.77 1.075 9.26 1.245 ;
      RECT 8.53 1.725 8.86 1.895 ;
      RECT 7.77 1.555 8.78 1.725 ;
      RECT 7.77 1.075 7.94 1.725 ;
      RECT 7.89 0.995 8.06 1.325 ;
      RECT 7.05 1.725 7.38 1.895 ;
      RECT 5.13 1.725 6.42 1.895 ;
      RECT 6.17 1.64 7.3 1.81 ;
      RECT 6.89 0.715 7.3 0.885 ;
      RECT 7.13 0.255 7.3 0.885 ;
      RECT 7.13 1.075 7.3 1.445 ;
      RECT 6.81 1.075 7.3 1.245 ;
      RECT 4.37 1.075 5.7 1.245 ;
      RECT 5.45 0.995 5.62 1.245 ;
      RECT 4.45 0.675 4.62 0.885 ;
      RECT 4.45 0.675 4.94 0.845 ;
      RECT 3.13 1.835 3.42 2.005 ;
      RECT 3.13 1.075 3.3 2.005 ;
      RECT 2.93 1.075 3.3 1.245 ;
      RECT 1.93 1.075 2.42 1.245 ;
      RECT 2.25 0.995 2.42 1.245 ;
      RECT 2.01 1.835 2.42 2.005 ;
      RECT 2.25 1.645 2.42 2.005 ;
      RECT 1.05 1.555 1.7 1.725 ;
      RECT 1.05 0.995 1.22 1.725 ;
      RECT 0.69 2.115 0.98 2.285 ;
      RECT 0.69 1.075 0.86 2.285 ;
      RECT 0.49 1.075 0.86 1.245 ;
      RECT 8.37 0.995 8.54 1.325 ;
      RECT 7.65 0.255 7.82 0.605 ;
      RECT 7.65 1.985 7.82 2.315 ;
      RECT 6.65 1.985 6.82 2.315 ;
      RECT 6.41 0.995 6.58 1.445 ;
      RECT 5.93 0.995 6.1 1.325 ;
      RECT 5.21 0.255 5.38 0.605 ;
      RECT 4.21 1.645 4.38 2.005 ;
      RECT 3.97 0.995 4.14 1.445 ;
      RECT 3.49 0.995 3.66 1.325 ;
      RECT 3.25 0.255 3.42 0.605 ;
      RECT 2.77 1.555 2.94 1.975 ;
      RECT 1.77 0.255 1.94 0.605 ;
      RECT 1.53 0.995 1.7 1.325 ;
      RECT 0.81 0.255 0.98 0.605 ;
      RECT 0.33 1.555 0.5 1.975 ;
  END
END scs130hd_mpr2ea_8

MACRO scs130hd_mpr2et_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130hd_mpr2et_8 0 0 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT 9.305 2.035 9.86 2.365 ;
      RECT 9.305 0.37 9.605 2.365 ;
      RECT 5.37 1.475 5.925 1.805 ;
      RECT 5.625 0.37 5.925 1.805 ;
      RECT 5.625 0.37 9.605 0.67 ;
      RECT 10.49 0.355 11.22 0.685 ;
      RECT 8.27 2.035 9 2.365 ;
      RECT 6.57 2.035 7.3 2.365 ;
      RECT 4.13 0.915 4.86 1.245 ;
      RECT 2.69 1.475 3.42 1.805 ;
      RECT 1.615 0.915 2.345 1.245 ;
      RECT 0.58 0.915 1.31 1.245 ;
      RECT 0.25 2.035 0.98 2.365 ;
    LAYER via2 ;
      RECT 10.555 0.42 10.755 0.62 ;
      RECT 9.595 2.1 9.795 2.3 ;
      RECT 8.595 2.1 8.795 2.3 ;
      RECT 6.635 2.1 6.835 2.3 ;
      RECT 5.435 1.54 5.635 1.74 ;
      RECT 4.195 0.98 4.395 1.18 ;
      RECT 2.755 1.54 2.955 1.74 ;
      RECT 2.015 0.98 2.215 1.18 ;
      RECT 0.795 0.98 0.995 1.18 ;
      RECT 0.315 2.1 0.515 2.3 ;
    LAYER met2 ;
      RECT 9.085 1.48 9.345 1.8 ;
      RECT 9.145 0.36 9.285 1.8 ;
      RECT 9.085 0.36 9.345 0.68 ;
      RECT 8.085 2.04 8.345 2.36 ;
      RECT 8.085 1.455 8.285 2.36 ;
      RECT 8.025 0.36 8.165 1.99 ;
      RECT 8.025 1.455 8.525 1.825 ;
      RECT 7.965 0.36 8.225 0.68 ;
      RECT 7.605 2.04 7.865 2.36 ;
      RECT 7.665 0.45 7.805 2.36 ;
      RECT 7.365 0.45 7.805 0.68 ;
      RECT 7.365 0.36 7.625 0.68 ;
      RECT 7.125 0.92 7.385 1.24 ;
      RECT 6.545 1.01 7.385 1.15 ;
      RECT 6.545 0.07 6.685 1.15 ;
      RECT 3.205 0.36 3.465 0.68 ;
      RECT 3.205 0.45 4.245 0.59 ;
      RECT 4.105 0.07 4.245 0.59 ;
      RECT 4.105 0.07 6.685 0.21 ;
      RECT 6.595 2.015 6.875 2.385 ;
      RECT 6.665 1.57 6.805 2.385 ;
      RECT 6.475 1.455 6.755 1.825 ;
      RECT 6.185 1.57 6.805 1.71 ;
      RECT 6.185 0.36 6.325 1.71 ;
      RECT 6.125 0.36 6.385 0.68 ;
      RECT 5.395 1.455 5.675 1.825 ;
      RECT 5.465 0.36 5.605 1.825 ;
      RECT 5.405 0.36 5.665 0.68 ;
      RECT 5.045 2.04 5.305 2.36 ;
      RECT 5.105 0.45 5.245 2.36 ;
      RECT 4.685 0.36 4.945 0.68 ;
      RECT 4.685 0.45 5.245 0.59 ;
      RECT 2.715 1.455 2.995 1.825 ;
      RECT 4.685 1.48 4.945 1.8 ;
      RECT 2.365 1.48 2.995 1.8 ;
      RECT 2.365 1.57 4.945 1.71 ;
      RECT 4.155 0.895 4.435 1.265 ;
      RECT 4.155 0.92 4.685 1.24 ;
      RECT 1.725 1.48 1.985 1.8 ;
      RECT 1.665 1.01 1.805 1.71 ;
      RECT 1.975 0.895 2.255 1.265 ;
      RECT 3.445 0.92 3.705 1.24 ;
      RECT 1.665 1.01 3.705 1.15 ;
      RECT 1.245 1.48 1.505 1.8 ;
      RECT 1.305 0.36 1.445 1.8 ;
      RECT 1.245 0.36 1.505 0.68 ;
      RECT 0.275 2.015 0.555 2.385 ;
      RECT 0.285 1.76 0.545 2.385 ;
      RECT 10.515 0.335 10.795 0.705 ;
      RECT 9.555 2.015 9.835 2.385 ;
      RECT 8.555 2.015 8.835 2.385 ;
      RECT 0.755 0.895 1.035 1.265 ;
    LAYER via1 ;
      RECT 10.58 0.445 10.73 0.595 ;
      RECT 9.62 2.125 9.77 2.275 ;
      RECT 9.14 0.445 9.29 0.595 ;
      RECT 9.14 1.565 9.29 1.715 ;
      RECT 8.62 2.125 8.77 2.275 ;
      RECT 8.14 2.125 8.29 2.275 ;
      RECT 8.02 0.445 8.17 0.595 ;
      RECT 7.66 2.125 7.81 2.275 ;
      RECT 7.42 0.445 7.57 0.595 ;
      RECT 7.18 1.005 7.33 1.155 ;
      RECT 6.66 2.125 6.81 2.275 ;
      RECT 6.18 0.445 6.33 0.595 ;
      RECT 5.46 0.445 5.61 0.595 ;
      RECT 5.46 1.565 5.61 1.715 ;
      RECT 5.1 2.125 5.25 2.275 ;
      RECT 4.74 0.445 4.89 0.595 ;
      RECT 4.74 1.565 4.89 1.715 ;
      RECT 4.48 1.005 4.63 1.155 ;
      RECT 3.5 1.005 3.65 1.155 ;
      RECT 3.26 0.445 3.41 0.595 ;
      RECT 2.42 1.565 2.57 1.715 ;
      RECT 1.78 1.565 1.93 1.715 ;
      RECT 1.3 0.445 1.45 0.595 ;
      RECT 1.3 1.565 1.45 1.715 ;
      RECT 0.82 1.005 0.97 1.155 ;
      RECT 0.34 1.845 0.49 1.995 ;
    LAYER met1 ;
      RECT 9.535 2.07 9.855 2.33 ;
      RECT 10.825 1.245 10.965 2.105 ;
      RECT 9.625 1.965 10.965 2.105 ;
      RECT 9.625 1.525 9.765 2.33 ;
      RECT 9.55 1.525 9.84 1.755 ;
      RECT 10.75 1.245 11.04 1.475 ;
      RECT 10.27 1.525 10.56 1.755 ;
      RECT 10.465 0.45 10.605 1.71 ;
      RECT 10.495 0.39 10.815 0.65 ;
      RECT 7.095 0.95 7.415 1.21 ;
      RECT 9.79 0.965 10.08 1.195 ;
      RECT 7.185 0.87 10.005 1.01 ;
      RECT 9.055 0.39 9.375 0.65 ;
      RECT 9.55 0.405 9.84 0.635 ;
      RECT 9.055 0.45 9.84 0.59 ;
      RECT 9.055 1.51 9.375 1.77 ;
      RECT 9.055 1.29 9.285 1.77 ;
      RECT 8.55 1.245 8.84 1.475 ;
      RECT 8.55 1.29 9.285 1.43 ;
      RECT 7.575 2.07 7.895 2.33 ;
      RECT 7.11 2.085 7.4 2.315 ;
      RECT 7.11 2.13 7.895 2.27 ;
      RECT 5.87 0.965 6.16 1.195 ;
      RECT 5.87 1.01 6.805 1.15 ;
      RECT 6.665 0.45 6.805 1.15 ;
      RECT 7.335 0.39 7.655 0.65 ;
      RECT 7.11 0.405 7.655 0.635 ;
      RECT 6.665 0.45 7.655 0.59 ;
      RECT 5.015 2.07 5.335 2.33 ;
      RECT 5.015 2.13 6.085 2.27 ;
      RECT 5.945 1.57 6.085 2.27 ;
      RECT 7.11 1.525 7.4 1.755 ;
      RECT 5.945 1.57 7.4 1.71 ;
      RECT 5.375 0.39 5.695 0.65 ;
      RECT 5.15 0.405 5.695 0.635 ;
      RECT 4.395 0.95 4.715 1.21 ;
      RECT 5.39 0.965 5.68 1.195 ;
      RECT 4.15 0.965 4.715 1.195 ;
      RECT 4.15 1.01 5.68 1.15 ;
      RECT 3.67 1.525 3.96 1.755 ;
      RECT 3.865 0.45 4.005 1.71 ;
      RECT 4.655 0.39 4.975 0.65 ;
      RECT 3.67 0.405 3.96 0.635 ;
      RECT 3.67 0.45 4.975 0.59 ;
      RECT 3.265 1.965 4.365 2.105 ;
      RECT 4.15 1.805 4.44 2.035 ;
      RECT 3.19 1.805 3.48 2.035 ;
      RECT 3.43 0.87 3.72 1.24 ;
      RECT 2.665 0.87 3.72 1.01 ;
      RECT 3.175 0.39 3.495 0.65 ;
      RECT 1.215 0.39 1.535 0.65 ;
      RECT 1.215 0.45 3.495 0.59 ;
      RECT 2.335 1.51 2.655 1.77 ;
      RECT 2.335 1.51 3.165 1.65 ;
      RECT 2.95 1.245 3.165 1.65 ;
      RECT 2.95 1.245 3.24 1.475 ;
      RECT 0.735 0.95 1.055 1.21 ;
      RECT 2.145 0.965 2.435 1.195 ;
      RECT 0.735 0.965 1.28 1.195 ;
      RECT 0.735 1.05 1.685 1.19 ;
      RECT 1.545 0.87 1.685 1.19 ;
      RECT 2.045 0.965 2.435 1.15 ;
      RECT 1.545 0.87 2.185 1.01 ;
      RECT 0.255 1.76 0.575 2.175 ;
      RECT 0.335 0.405 0.49 2.175 ;
      RECT 0.27 0.405 0.56 0.635 ;
      RECT 0 -0.24 11.96 0.24 ;
      RECT 0 2.48 11.96 2.96 ;
      RECT 8.535 2.07 8.855 2.33 ;
      RECT 7.935 0.39 8.615 0.65 ;
      RECT 8.055 2.07 8.375 2.33 ;
      RECT 6.575 2.07 6.895 2.33 ;
      RECT 6.095 0.39 6.415 0.65 ;
      RECT 5.375 1.51 5.695 1.77 ;
      RECT 4.655 1.51 4.975 1.77 ;
      RECT 1.695 1.51 2.015 1.77 ;
      RECT 1.215 1.51 1.535 1.77 ;
    LAYER mcon ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.645 2.635 11.815 2.805 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 11.185 2.635 11.355 2.805 ;
      RECT 10.81 1.275 10.98 1.445 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.725 2.635 10.895 2.805 ;
      RECT 10.57 0.435 10.74 0.605 ;
      RECT 10.33 1.555 10.5 1.725 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 10.265 2.635 10.435 2.805 ;
      RECT 9.85 0.995 10.02 1.165 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.805 2.635 9.975 2.805 ;
      RECT 9.61 0.435 9.78 0.605 ;
      RECT 9.61 1.555 9.78 1.725 ;
      RECT 9.61 2.115 9.78 2.285 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 9.345 2.635 9.515 2.805 ;
      RECT 9.13 1.555 9.3 1.725 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.885 2.635 9.055 2.805 ;
      RECT 8.61 1.275 8.78 1.445 ;
      RECT 8.61 2.115 8.78 2.285 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 8.13 0.435 8.3 0.605 ;
      RECT 8.13 2.115 8.3 2.285 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.17 0.435 7.34 0.605 ;
      RECT 7.17 0.995 7.34 1.165 ;
      RECT 7.17 1.555 7.34 1.725 ;
      RECT 7.17 2.115 7.34 2.285 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 6.65 2.115 6.82 2.285 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.17 0.435 6.34 0.605 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 5.93 0.995 6.1 1.165 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.45 0.995 5.62 1.165 ;
      RECT 5.45 1.555 5.62 1.725 ;
      RECT 5.21 0.435 5.38 0.605 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.73 1.555 4.9 1.725 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 4.21 0.995 4.38 1.165 ;
      RECT 4.21 1.835 4.38 2.005 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 3.73 0.435 3.9 0.605 ;
      RECT 3.73 1.555 3.9 1.725 ;
      RECT 3.49 0.995 3.66 1.165 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.25 1.835 3.42 2.005 ;
      RECT 3.01 1.275 3.18 1.445 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.205 0.995 2.375 1.165 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 1.77 1.555 1.94 1.725 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.29 0.435 1.46 0.605 ;
      RECT 1.29 1.555 1.46 1.725 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.05 0.995 1.22 1.165 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.33 0.435 0.5 0.605 ;
      RECT 0.33 1.975 0.5 2.145 ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
    LAYER li ;
      RECT 11.05 -0.085 11.22 0.585 ;
      RECT 10.09 -0.085 10.26 0.585 ;
      RECT 9.13 -0.085 9.3 0.585 ;
      RECT 8.61 -0.085 8.78 0.585 ;
      RECT 7.65 -0.085 7.82 0.585 ;
      RECT 6.65 -0.085 6.82 0.585 ;
      RECT 5.69 -0.085 5.86 0.585 ;
      RECT 4.21 -0.085 4.38 0.585 ;
      RECT 2.29 -0.085 2.46 0.585 ;
      RECT 0.81 -0.085 0.98 0.585 ;
      RECT 0 -0.085 11.96 0.085 ;
      RECT 0 2.635 11.96 2.805 ;
      RECT 10.09 2.135 10.26 2.805 ;
      RECT 7.65 2.135 7.82 2.805 ;
      RECT 5.69 2.135 5.86 2.805 ;
      RECT 4.73 2.135 4.9 2.805 ;
      RECT 2.77 2.135 2.94 2.805 ;
      RECT 1.77 2.135 1.94 2.805 ;
      RECT 0.81 2.135 0.98 2.805 ;
      RECT 10.33 1.725 11.3 1.895 ;
      RECT 10.33 1.555 10.5 1.895 ;
      RECT 9.85 0.995 10.02 1.325 ;
      RECT 9.85 1.075 10.58 1.245 ;
      RECT 9.49 2.115 9.78 2.285 ;
      RECT 9.49 1.075 9.66 2.285 ;
      RECT 9.49 1.555 9.78 1.725 ;
      RECT 9.29 1.075 9.66 1.245 ;
      RECT 8.61 1.175 8.78 1.445 ;
      RECT 8.37 1.175 8.78 1.345 ;
      RECT 8.29 1.075 8.62 1.245 ;
      RECT 8.13 2.115 8.78 2.285 ;
      RECT 8.61 1.645 8.78 2.285 ;
      RECT 8.49 1.725 8.78 2.285 ;
      RECT 7.17 1.415 7.34 1.725 ;
      RECT 7.17 1.415 8.06 1.585 ;
      RECT 7.89 0.995 8.06 1.585 ;
      RECT 7.17 1.075 7.66 1.245 ;
      RECT 7.17 0.995 7.34 1.245 ;
      RECT 5.13 1.725 5.62 1.895 ;
      RECT 6.29 1.075 6.46 1.725 ;
      RECT 5.45 1.555 6.46 1.725 ;
      RECT 6.41 0.995 6.58 1.325 ;
      RECT 5.21 0.335 5.38 0.605 ;
      RECT 4.65 0.335 5.38 0.505 ;
      RECT 4.73 1.075 4.9 1.725 ;
      RECT 4.73 1.075 5.22 1.245 ;
      RECT 3.89 1.075 4.38 1.245 ;
      RECT 4.21 0.995 4.38 1.245 ;
      RECT 3.73 0.335 3.9 0.605 ;
      RECT 3.17 0.335 3.9 0.505 ;
      RECT 3.25 1.725 3.42 2.005 ;
      RECT 2.21 1.725 3.5 1.895 ;
      RECT 2.205 1.075 2.78 1.245 ;
      RECT 2.205 0.995 2.375 1.245 ;
      RECT 1.29 0.335 1.46 0.605 ;
      RECT 1.29 0.335 2.02 0.505 ;
      RECT 1.65 1.555 1.94 1.725 ;
      RECT 1.65 1.075 1.82 1.725 ;
      RECT 1.45 1.075 1.82 1.245 ;
      RECT 1.29 1.555 1.46 1.975 ;
      RECT 0.67 1.64 1.46 1.81 ;
      RECT 0.67 1.415 0.84 1.81 ;
      RECT 0.57 0.995 0.74 1.585 ;
      RECT 0.33 1.075 0.74 1.345 ;
      RECT 10.81 0.995 10.98 1.445 ;
      RECT 10.57 0.255 10.74 0.605 ;
      RECT 9.61 0.255 9.78 0.605 ;
      RECT 9.13 1.555 9.3 1.975 ;
      RECT 8.13 0.255 8.3 0.605 ;
      RECT 7.17 0.255 7.34 0.605 ;
      RECT 7.17 1.985 7.34 2.315 ;
      RECT 6.65 1.645 6.82 2.285 ;
      RECT 6.17 0.255 6.34 0.605 ;
      RECT 5.93 0.995 6.1 1.325 ;
      RECT 5.45 0.995 5.62 1.325 ;
      RECT 4.21 1.645 4.38 2.005 ;
      RECT 3.73 1.555 3.9 1.975 ;
      RECT 3.49 0.995 3.66 1.325 ;
      RECT 3.01 0.995 3.18 1.445 ;
      RECT 1.05 0.995 1.22 1.325 ;
      RECT 0.33 0.255 0.5 0.605 ;
      RECT 0.33 1.785 0.5 2.145 ;
  END
END scs130hd_mpr2et_8

MACRO scs130hd_mpr2xa_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130hd_mpr2xa_8 0 0 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met4 ;
      RECT 2.15 1.475 2.48 1.805 ;
      RECT 2.165 1 2.48 1.805 ;
      RECT 4.31 0.985 4.64 1.34 ;
      RECT 2.165 1 4.64 1.3 ;
    LAYER via3 ;
      RECT 4.375 1.075 4.575 1.275 ;
      RECT 2.215 1.54 2.415 1.74 ;
    LAYER met3 ;
      RECT 4.79 2.01 5.12 2.365 ;
      RECT 2.885 2.05 5.12 2.35 ;
      RECT 2.885 0.915 3.185 2.35 ;
      RECT 2.87 0.915 3.2 1.245 ;
      RECT 3.86 1.02 4.64 1.365 ;
      RECT 4.335 0.985 4.64 1.365 ;
      RECT 4.315 1.015 4.64 1.365 ;
      RECT 2.155 0.915 2.475 1.83 ;
      RECT 2.155 0.915 2.485 1.45 ;
      RECT 7.71 0.355 8.44 0.685 ;
      RECT 6.02 0.37 6.75 0.7 ;
      RECT 4.985 0.355 5.715 0.705 ;
      RECT 3.435 0.38 4.165 0.71 ;
      RECT 0.965 1.475 1.695 1.805 ;
      RECT 0.83 0.355 1.56 0.685 ;
    LAYER via2 ;
      RECT 7.945 0.42 8.145 0.62 ;
      RECT 6.085 0.435 6.285 0.635 ;
      RECT 5.065 0.44 5.265 0.64 ;
      RECT 4.855 2.075 5.055 2.275 ;
      RECT 4.375 1.075 4.575 1.275 ;
      RECT 3.625 0.445 3.825 0.645 ;
      RECT 2.935 0.98 3.135 1.18 ;
      RECT 2.22 0.98 2.42 1.18 ;
      RECT 1.255 1.54 1.455 1.74 ;
      RECT 1.015 0.42 1.215 0.62 ;
    LAYER met2 ;
      RECT 7.915 2.04 8.175 2.36 ;
      RECT 7.975 0.335 8.115 2.36 ;
      RECT 7.8 0.895 8.115 1.265 ;
      RECT 7.87 0.45 8.115 1.265 ;
      RECT 7.905 0.335 8.185 0.705 ;
      RECT 7.225 0.92 7.485 1.24 ;
      RECT 6.565 1.01 7.485 1.15 ;
      RECT 6.565 0.07 6.705 1.15 ;
      RECT 3.025 0.36 3.285 0.68 ;
      RECT 3.205 0.07 3.345 0.59 ;
      RECT 3.205 0.07 6.705 0.21 ;
      RECT 6.055 1.76 6.315 2.08 ;
      RECT 6.115 0.35 6.255 2.08 ;
      RECT 6.045 0.35 6.325 0.72 ;
      RECT 3.445 2.51 5.88 2.65 ;
      RECT 5.74 1.2 5.88 2.65 ;
      RECT 3.445 2.13 3.585 2.65 ;
      RECT 3.145 2.13 3.585 2.36 ;
      RECT 0.805 2.13 3.585 2.27 ;
      RECT 3.145 2.04 3.405 2.36 ;
      RECT 0.805 1.85 0.945 2.27 ;
      RECT 0.295 1.76 0.555 2.08 ;
      RECT 0.295 1.85 0.945 1.99 ;
      RECT 0.355 0.36 0.495 2.08 ;
      RECT 5.68 1.2 5.94 1.52 ;
      RECT 0.295 0.36 0.555 0.68 ;
      RECT 5.305 2.04 5.565 2.36 ;
      RECT 5.365 0.45 5.505 2.36 ;
      RECT 5.025 0.45 5.505 0.725 ;
      RECT 4.825 0.355 5.305 0.7 ;
      RECT 4.815 1.99 5.095 2.36 ;
      RECT 4.885 0.895 5.025 2.36 ;
      RECT 4.825 0.895 5.085 1.52 ;
      RECT 4.815 0.895 5.095 1.265 ;
      RECT 3.745 2.04 4.005 2.36 ;
      RECT 3.745 1.85 3.945 2.36 ;
      RECT 3.55 1.85 3.945 1.99 ;
      RECT 3.55 0.36 3.69 1.99 ;
      RECT 3.55 0.36 3.865 0.73 ;
      RECT 3.49 0.36 3.865 0.68 ;
      RECT 1.215 1.455 1.495 1.825 ;
      RECT 2.665 1.48 2.925 1.8 ;
      RECT 1.045 1.57 2.925 1.71 ;
      RECT 1.045 1.455 1.495 1.71 ;
      RECT 0.985 0.895 1.245 1.52 ;
      RECT 0.975 0.895 1.255 1.265 ;
      RECT 2.055 0.895 2.465 1.265 ;
      RECT 1.465 0.92 1.725 1.24 ;
      RECT 1.465 1.01 2.465 1.15 ;
      RECT 0.975 0.335 1.255 0.705 ;
      RECT 0.975 0.36 1.365 0.68 ;
      RECT 4.335 0.895 4.615 1.36 ;
      RECT 4.095 0.36 4.375 0.705 ;
      RECT 2.895 0.895 3.175 1.265 ;
    LAYER via1 ;
      RECT 7.97 0.445 8.12 0.595 ;
      RECT 7.97 2.125 8.12 2.275 ;
      RECT 7.28 1.005 7.43 1.155 ;
      RECT 6.11 0.445 6.26 0.595 ;
      RECT 6.11 1.845 6.26 1.995 ;
      RECT 5.735 1.285 5.885 1.435 ;
      RECT 5.36 2.125 5.51 2.275 ;
      RECT 4.88 0.445 5.03 0.595 ;
      RECT 4.88 1.285 5.03 1.435 ;
      RECT 4.4 1.005 4.55 1.155 ;
      RECT 4.16 0.445 4.31 0.595 ;
      RECT 3.8 2.125 3.95 2.275 ;
      RECT 3.545 0.445 3.695 0.595 ;
      RECT 3.2 2.125 3.35 2.275 ;
      RECT 3.08 0.445 3.23 0.595 ;
      RECT 2.96 1.005 3.11 1.155 ;
      RECT 2.72 1.565 2.87 1.715 ;
      RECT 1.52 1.005 1.67 1.155 ;
      RECT 1.16 0.445 1.31 0.595 ;
      RECT 1.04 1.285 1.19 1.435 ;
      RECT 0.35 0.445 0.5 0.595 ;
      RECT 0.35 1.845 0.5 1.995 ;
    LAYER met1 ;
      RECT 7.885 0.39 8.205 0.65 ;
      RECT 7.45 0.405 7.74 0.635 ;
      RECT 7.45 0.45 8.205 0.59 ;
      RECT 7.885 2.07 8.205 2.33 ;
      RECT 7.45 2.085 7.74 2.315 ;
      RECT 7.45 2.13 8.205 2.27 ;
      RECT 7.21 1.525 7.5 1.755 ;
      RECT 7.21 1.57 7.785 1.71 ;
      RECT 7.645 1.43 7.905 1.57 ;
      RECT 7.69 1.245 7.98 1.475 ;
      RECT 5.845 1.43 6.945 1.57 ;
      RECT 5.65 1.23 5.97 1.49 ;
      RECT 6.73 1.245 7.02 1.475 ;
      RECT 5.65 1.245 6.06 1.49 ;
      RECT 6.025 0.39 6.345 0.65 ;
      RECT 6.49 0.405 6.78 0.635 ;
      RECT 6.025 0.45 6.78 0.59 ;
      RECT 3.325 1.655 5.505 1.795 ;
      RECT 5.365 0.665 5.505 1.795 ;
      RECT 3.325 1.57 4.62 1.795 ;
      RECT 4.33 1.525 4.62 1.795 ;
      RECT 3.325 1.29 3.66 1.795 ;
      RECT 3.37 1.245 3.66 1.795 ;
      RECT 6.25 0.965 6.54 1.195 ;
      RECT 5.365 0.87 6.465 1.01 ;
      RECT 5.29 0.665 5.58 0.915 ;
      RECT 5.275 2.07 5.595 2.33 ;
      RECT 5.275 2.085 5.79 2.315 ;
      RECT 3.85 0.965 4.14 1.195 ;
      RECT 4 0.57 4.14 1.195 ;
      RECT 4 0.57 4.305 0.71 ;
      RECT 4.795 0.39 5.115 0.65 ;
      RECT 4.075 0.39 4.395 0.65 ;
      RECT 4.57 0.405 5.115 0.635 ;
      RECT 4.075 0.45 5.115 0.59 ;
      RECT 3.715 2.07 4.035 2.33 ;
      RECT 3.61 2.085 4.035 2.315 ;
      RECT 1.69 1.525 1.98 1.755 ;
      RECT 1.69 1.525 2.145 1.71 ;
      RECT 2.005 1.05 2.145 1.71 ;
      RECT 2.125 0.45 2.265 1.19 ;
      RECT 2.995 0.39 3.315 0.65 ;
      RECT 2.17 0.405 2.46 0.635 ;
      RECT 2.125 0.45 3.315 0.59 ;
      RECT 2.875 0.95 3.195 1.21 ;
      RECT 2.41 0.965 2.7 1.195 ;
      RECT 2.41 1.01 3.195 1.15 ;
      RECT 2.635 1.51 2.955 1.77 ;
      RECT 2.635 1.525 3.18 1.755 ;
      RECT 2.17 2.085 2.46 2.315 ;
      RECT 1.285 1.965 2.385 2.105 ;
      RECT 1.21 1.805 1.5 2.035 ;
      RECT 0.49 1.245 0.78 1.475 ;
      RECT 0.565 0.87 0.705 1.475 ;
      RECT 0.565 0.87 1.185 1.01 ;
      RECT 1.045 0.45 1.185 1.01 ;
      RECT 0.805 0.45 1.185 0.71 ;
      RECT 1.075 0.39 1.395 0.65 ;
      RECT 1.69 0.405 1.98 0.635 ;
      RECT 0.805 0.45 1.98 0.59 ;
      RECT 0 -0.24 8.74 0.24 ;
      RECT 0 2.48 8.74 2.96 ;
      RECT 7.195 0.95 7.515 1.21 ;
      RECT 6.025 1.79 6.345 2.05 ;
      RECT 4.795 1.23 5.115 1.49 ;
      RECT 4.315 0.95 4.635 1.21 ;
      RECT 3.46 0.39 3.86 0.65 ;
      RECT 3.115 2.07 3.435 2.33 ;
      RECT 1.435 0.95 1.755 1.21 ;
      RECT 0.955 1.23 1.275 1.49 ;
      RECT 0.265 0.39 0.585 0.65 ;
      RECT 0.265 1.79 0.585 2.05 ;
    LAYER mcon ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 7.75 1.275 7.92 1.445 ;
      RECT 7.51 0.435 7.68 0.605 ;
      RECT 7.51 2.115 7.68 2.285 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.27 0.995 7.44 1.165 ;
      RECT 7.27 1.555 7.44 1.725 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 6.79 1.275 6.96 1.445 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.55 0.435 6.72 0.605 ;
      RECT 6.31 0.995 6.48 1.165 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 6.1 1.835 6.27 2.005 ;
      RECT 5.83 1.275 6 1.445 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.56 2.115 5.73 2.285 ;
      RECT 5.35 0.695 5.52 0.865 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 4.87 1.275 5.04 1.445 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.63 0.435 4.8 0.605 ;
      RECT 4.39 0.995 4.56 1.165 ;
      RECT 4.39 1.555 4.56 1.725 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 3.91 0.995 4.08 1.165 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 3.67 2.115 3.84 2.285 ;
      RECT 3.63 0.435 3.8 0.605 ;
      RECT 3.43 1.275 3.6 1.445 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.19 2.115 3.36 2.285 ;
      RECT 2.95 1.555 3.12 1.725 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.47 0.995 2.64 1.165 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 2.23 0.435 2.4 0.605 ;
      RECT 2.23 2.115 2.4 2.285 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 1.75 0.435 1.92 0.605 ;
      RECT 1.75 1.555 1.92 1.725 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.51 0.995 1.68 1.165 ;
      RECT 1.27 1.835 1.44 2.005 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.03 1.275 1.2 1.445 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.55 1.275 0.72 1.445 ;
      RECT 0.34 0.435 0.51 0.605 ;
      RECT 0.34 1.835 0.51 2.005 ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
    LAYER li ;
      RECT 7.97 -0.085 8.14 0.585 ;
      RECT 7.03 -0.085 7.2 0.585 ;
      RECT 6.07 -0.085 6.24 0.585 ;
      RECT 4.15 -0.085 4.32 0.585 ;
      RECT 3.19 -0.085 3.36 0.585 ;
      RECT 1.27 -0.085 1.44 0.585 ;
      RECT 0 -0.085 8.74 0.085 ;
      RECT 0 2.635 8.74 2.805 ;
      RECT 7.03 2.135 7.2 2.805 ;
      RECT 5.11 2.135 5.28 2.805 ;
      RECT 4.17 2.135 4.34 2.805 ;
      RECT 2.71 2.135 2.88 2.805 ;
      RECT 0.79 2.135 0.96 2.805 ;
      RECT 7.51 2.115 8.025 2.285 ;
      RECT 7.855 1.725 8.025 2.285 ;
      RECT 7.96 1.645 8.13 1.975 ;
      RECT 7.75 1.035 8.025 1.445 ;
      RECT 7.63 1.035 8.025 1.245 ;
      RECT 6.1 1.645 6.27 2.005 ;
      RECT 6.1 1.725 7.44 1.895 ;
      RECT 7.27 1.555 7.44 1.895 ;
      RECT 5.83 1.075 6 1.445 ;
      RECT 5.35 1.075 6 1.345 ;
      RECT 5.27 1.075 6.08 1.245 ;
      RECT 4.63 0.315 4.8 0.605 ;
      RECT 4.63 0.315 5.87 0.485 ;
      RECT 5.35 0.655 5.52 0.865 ;
      RECT 4.99 0.655 5.52 0.825 ;
      RECT 4.39 1.725 4.88 1.895 ;
      RECT 4.39 1.555 4.56 1.895 ;
      RECT 3.67 1.725 3.84 2.285 ;
      RECT 3.56 1.725 3.89 1.895 ;
      RECT 3.63 0.335 3.8 0.605 ;
      RECT 3.67 0.255 3.84 0.585 ;
      RECT 3.535 0.335 3.84 0.555 ;
      RECT 2.11 1.725 2.4 2.285 ;
      RECT 2.23 1.645 2.4 2.285 ;
      RECT 1.87 1.075 2.24 1.245 ;
      RECT 1.87 0.435 2.04 1.245 ;
      RECT 1.75 0.435 2.04 0.605 ;
      RECT 7.51 0.255 7.68 0.605 ;
      RECT 7.27 0.995 7.44 1.325 ;
      RECT 6.79 0.995 6.96 1.445 ;
      RECT 6.55 0.255 6.72 0.605 ;
      RECT 6.31 0.995 6.48 1.325 ;
      RECT 5.56 1.985 5.73 2.315 ;
      RECT 4.87 0.995 5.04 1.445 ;
      RECT 4.39 0.995 4.56 1.325 ;
      RECT 3.91 0.995 4.08 1.325 ;
      RECT 3.43 0.995 3.6 1.445 ;
      RECT 3.19 1.985 3.36 2.315 ;
      RECT 2.95 0.995 3.12 1.725 ;
      RECT 2.47 0.995 2.64 1.325 ;
      RECT 2.23 0.255 2.4 0.605 ;
      RECT 1.75 1.555 1.92 1.975 ;
      RECT 1.51 0.995 1.68 1.325 ;
      RECT 1.27 1.645 1.44 2.005 ;
      RECT 1.03 0.995 1.2 1.445 ;
      RECT 0.55 0.995 0.72 1.445 ;
      RECT 0.34 0.255 0.51 0.605 ;
      RECT 0.34 1.645 0.51 2.005 ;
  END
END scs130hd_mpr2xa_8

MACRO scs130hd_mpr2ya_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN scs130hd_mpr2ya_8 0 0 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT 7.55 0.515 7.88 1.245 ;
      RECT 6.35 1.38 6.68 2.11 ;
      RECT 5.51 0.355 6.24 0.685 ;
      RECT 4.07 0.355 4.8 0.685 ;
      RECT 4.43 1.26 4.76 1.99 ;
      RECT 3.11 0.355 3.44 1.085 ;
      RECT 1.91 0.515 2.24 1.245 ;
      RECT 1.19 0.515 1.52 1.245 ;
    LAYER via2 ;
      RECT 7.615 0.98 7.815 1.18 ;
      RECT 6.415 1.54 6.615 1.74 ;
      RECT 5.575 0.42 5.775 0.62 ;
      RECT 4.495 1.325 4.695 1.525 ;
      RECT 4.135 0.42 4.335 0.62 ;
      RECT 3.175 0.42 3.375 0.62 ;
      RECT 1.975 0.98 2.175 1.18 ;
      RECT 1.255 0.98 1.455 1.18 ;
    LAYER met2 ;
      RECT 7.575 0.94 7.855 1.22 ;
      RECT 7.57 0.94 7.855 1.173 ;
      RECT 7.55 0.94 7.855 1.15 ;
      RECT 7.54 0.94 7.855 1.13 ;
      RECT 7.53 0.94 7.855 1.115 ;
      RECT 7.505 0.94 7.855 1.088 ;
      RECT 7.495 0.94 7.855 1.063 ;
      RECT 7.45 0.795 7.73 1.055 ;
      RECT 7.45 0.89 7.83 1.055 ;
      RECT 7.45 0.835 7.775 1.055 ;
      RECT 7.45 0.827 7.77 1.055 ;
      RECT 7.45 0.817 7.765 1.055 ;
      RECT 7.45 0.805 7.76 1.055 ;
      RECT 6.375 1.5 6.655 1.78 ;
      RECT 6.375 1.5 6.69 1.76 ;
      RECT 6.41 0.92 6.46 1.18 ;
      RECT 6.2 0.92 6.205 1.18 ;
      RECT 5.395 0.475 5.425 0.735 ;
      RECT 5.165 0.475 5.24 0.735 ;
      RECT 6.385 0.87 6.41 1.18 ;
      RECT 6.38 0.827 6.385 1.18 ;
      RECT 6.375 0.81 6.38 1.18 ;
      RECT 6.37 0.797 6.375 1.18 ;
      RECT 6.295 0.68 6.37 1.18 ;
      RECT 6.25 0.497 6.295 1.18 ;
      RECT 6.245 0.425 6.25 1.18 ;
      RECT 6.23 0.4 6.245 1.18 ;
      RECT 6.205 0.362 6.23 1.18 ;
      RECT 6.195 0.342 6.205 0.902 ;
      RECT 6.18 0.334 6.195 0.857 ;
      RECT 6.175 0.326 6.18 0.828 ;
      RECT 6.17 0.323 6.175 0.808 ;
      RECT 6.165 0.32 6.17 0.788 ;
      RECT 6.16 0.317 6.165 0.768 ;
      RECT 6.13 0.306 6.16 0.705 ;
      RECT 6.11 0.291 6.13 0.62 ;
      RECT 6.105 0.283 6.11 0.583 ;
      RECT 6.095 0.277 6.105 0.55 ;
      RECT 6.08 0.269 6.095 0.51 ;
      RECT 6.075 0.262 6.08 0.47 ;
      RECT 6.07 0.259 6.075 0.448 ;
      RECT 6.065 0.256 6.07 0.435 ;
      RECT 6.06 0.255 6.065 0.425 ;
      RECT 6.045 0.249 6.06 0.415 ;
      RECT 6.02 0.236 6.045 0.4 ;
      RECT 5.97 0.211 6.02 0.371 ;
      RECT 5.955 0.19 5.97 0.346 ;
      RECT 5.945 0.183 5.955 0.335 ;
      RECT 5.89 0.164 5.945 0.308 ;
      RECT 5.865 0.142 5.89 0.281 ;
      RECT 5.86 0.135 5.865 0.276 ;
      RECT 5.845 0.135 5.86 0.274 ;
      RECT 5.82 0.127 5.845 0.27 ;
      RECT 5.805 0.125 5.82 0.266 ;
      RECT 5.775 0.125 5.805 0.263 ;
      RECT 5.765 0.125 5.775 0.258 ;
      RECT 5.72 0.125 5.765 0.256 ;
      RECT 5.691 0.125 5.72 0.257 ;
      RECT 5.605 0.125 5.691 0.259 ;
      RECT 5.591 0.126 5.605 0.261 ;
      RECT 5.505 0.127 5.591 0.263 ;
      RECT 5.49 0.128 5.505 0.273 ;
      RECT 5.485 0.129 5.49 0.282 ;
      RECT 5.465 0.132 5.485 0.292 ;
      RECT 5.45 0.14 5.465 0.307 ;
      RECT 5.43 0.158 5.45 0.322 ;
      RECT 5.42 0.17 5.43 0.345 ;
      RECT 5.41 0.179 5.42 0.375 ;
      RECT 5.395 0.191 5.41 0.42 ;
      RECT 5.34 0.224 5.395 0.735 ;
      RECT 5.335 0.252 5.34 0.735 ;
      RECT 5.315 0.267 5.335 0.735 ;
      RECT 5.28 0.327 5.315 0.735 ;
      RECT 5.278 0.377 5.28 0.735 ;
      RECT 5.275 0.385 5.278 0.735 ;
      RECT 5.265 0.4 5.275 0.735 ;
      RECT 5.26 0.412 5.265 0.735 ;
      RECT 5.25 0.437 5.26 0.735 ;
      RECT 5.24 0.465 5.25 0.735 ;
      RECT 3.145 1.97 3.195 2.23 ;
      RECT 6.055 1.52 6.115 1.78 ;
      RECT 6.04 1.52 6.055 1.79 ;
      RECT 6.021 1.52 6.04 1.823 ;
      RECT 5.935 1.52 6.021 1.948 ;
      RECT 5.855 1.52 5.935 2.13 ;
      RECT 5.85 1.757 5.855 2.215 ;
      RECT 5.825 1.827 5.85 2.243 ;
      RECT 5.82 1.897 5.825 2.27 ;
      RECT 5.8 1.969 5.82 2.292 ;
      RECT 5.795 2.036 5.8 2.315 ;
      RECT 5.785 2.065 5.795 2.33 ;
      RECT 5.775 2.087 5.785 2.347 ;
      RECT 5.77 2.097 5.775 2.358 ;
      RECT 5.765 2.105 5.77 2.366 ;
      RECT 5.755 2.113 5.765 2.378 ;
      RECT 5.75 2.125 5.755 2.388 ;
      RECT 5.745 2.133 5.75 2.393 ;
      RECT 5.725 2.151 5.745 2.403 ;
      RECT 5.72 2.168 5.725 2.41 ;
      RECT 5.715 2.176 5.72 2.411 ;
      RECT 5.71 2.187 5.715 2.413 ;
      RECT 5.67 2.225 5.71 2.423 ;
      RECT 5.665 2.26 5.67 2.434 ;
      RECT 5.66 2.265 5.665 2.437 ;
      RECT 5.635 2.275 5.66 2.444 ;
      RECT 5.625 2.289 5.635 2.453 ;
      RECT 5.605 2.301 5.625 2.456 ;
      RECT 5.555 2.32 5.605 2.46 ;
      RECT 5.51 2.335 5.555 2.465 ;
      RECT 5.445 2.338 5.51 2.471 ;
      RECT 5.43 2.336 5.445 2.478 ;
      RECT 5.4 2.335 5.43 2.478 ;
      RECT 5.361 2.334 5.4 2.474 ;
      RECT 5.275 2.331 5.361 2.47 ;
      RECT 5.258 2.329 5.275 2.467 ;
      RECT 5.172 2.327 5.258 2.464 ;
      RECT 5.086 2.324 5.172 2.458 ;
      RECT 5 2.32 5.086 2.453 ;
      RECT 4.922 2.317 5 2.449 ;
      RECT 4.836 2.314 4.922 2.447 ;
      RECT 4.75 2.311 4.836 2.444 ;
      RECT 4.692 2.309 4.75 2.441 ;
      RECT 4.606 2.306 4.692 2.439 ;
      RECT 4.52 2.302 4.606 2.437 ;
      RECT 4.434 2.299 4.52 2.434 ;
      RECT 4.348 2.295 4.434 2.432 ;
      RECT 4.262 2.291 4.348 2.429 ;
      RECT 4.176 2.288 4.262 2.427 ;
      RECT 4.09 2.284 4.176 2.424 ;
      RECT 4.004 2.281 4.09 2.422 ;
      RECT 3.918 2.277 4.004 2.419 ;
      RECT 3.832 2.274 3.918 2.417 ;
      RECT 3.746 2.27 3.832 2.414 ;
      RECT 3.66 2.267 3.746 2.412 ;
      RECT 3.65 2.265 3.66 2.408 ;
      RECT 3.645 2.265 3.65 2.406 ;
      RECT 3.605 2.26 3.645 2.4 ;
      RECT 3.591 2.251 3.605 2.393 ;
      RECT 3.505 2.221 3.591 2.378 ;
      RECT 3.485 2.187 3.505 2.363 ;
      RECT 3.415 2.156 3.485 2.35 ;
      RECT 3.41 2.131 3.415 2.339 ;
      RECT 3.405 2.125 3.41 2.337 ;
      RECT 3.336 1.97 3.405 2.325 ;
      RECT 3.25 1.97 3.336 2.299 ;
      RECT 3.225 1.97 3.25 2.278 ;
      RECT 3.22 1.97 3.225 2.268 ;
      RECT 3.215 1.97 3.22 2.26 ;
      RECT 3.195 1.97 3.215 2.243 ;
      RECT 5.615 0.54 5.875 0.8 ;
      RECT 5.6 0.54 5.875 0.703 ;
      RECT 5.57 0.54 5.875 0.678 ;
      RECT 5.535 0.38 5.815 0.66 ;
      RECT 5.505 1.87 5.565 2.13 ;
      RECT 4.53 0.56 4.585 0.82 ;
      RECT 5.465 1.827 5.505 2.13 ;
      RECT 5.436 1.748 5.465 2.13 ;
      RECT 5.35 1.62 5.436 2.13 ;
      RECT 5.33 1.5 5.35 2.13 ;
      RECT 5.305 1.451 5.33 2.13 ;
      RECT 5.3 1.416 5.305 1.98 ;
      RECT 5.27 1.376 5.3 1.918 ;
      RECT 5.245 1.313 5.27 1.833 ;
      RECT 5.235 1.275 5.245 1.77 ;
      RECT 5.22 1.25 5.235 1.731 ;
      RECT 5.177 1.208 5.22 1.637 ;
      RECT 5.175 1.181 5.177 1.564 ;
      RECT 5.17 1.176 5.175 1.555 ;
      RECT 5.165 1.169 5.17 1.53 ;
      RECT 5.16 1.163 5.165 1.515 ;
      RECT 5.155 1.157 5.16 1.503 ;
      RECT 5.145 1.148 5.155 1.485 ;
      RECT 5.14 1.139 5.145 1.463 ;
      RECT 5.115 1.12 5.14 1.413 ;
      RECT 5.11 1.101 5.115 1.363 ;
      RECT 5.095 1.087 5.11 1.323 ;
      RECT 5.09 1.073 5.095 1.29 ;
      RECT 5.085 1.066 5.09 1.283 ;
      RECT 5.07 1.053 5.085 1.275 ;
      RECT 5.025 1.015 5.07 1.248 ;
      RECT 4.995 0.968 5.025 1.213 ;
      RECT 4.975 0.937 4.995 1.19 ;
      RECT 4.895 0.87 4.975 1.143 ;
      RECT 4.865 0.8 4.895 1.09 ;
      RECT 4.86 0.777 4.865 1.073 ;
      RECT 4.83 0.755 4.86 1.058 ;
      RECT 4.8 0.714 4.83 1.03 ;
      RECT 4.795 0.689 4.8 1.015 ;
      RECT 4.79 0.683 4.795 1.008 ;
      RECT 4.78 0.56 4.79 1 ;
      RECT 4.77 0.56 4.78 0.993 ;
      RECT 4.765 0.56 4.77 0.985 ;
      RECT 4.745 0.56 4.765 0.973 ;
      RECT 4.695 0.56 4.745 0.943 ;
      RECT 4.64 0.56 4.695 0.893 ;
      RECT 4.61 0.56 4.64 0.853 ;
      RECT 4.585 0.56 4.61 0.83 ;
      RECT 4.455 1.285 4.735 1.565 ;
      RECT 4.42 1.2 4.68 1.46 ;
      RECT 4.42 1.282 4.69 1.46 ;
      RECT 2.62 0.655 2.625 1.14 ;
      RECT 2.51 0.84 2.515 1.14 ;
      RECT 2.42 0.88 2.485 1.14 ;
      RECT 4.095 0.38 4.185 1.01 ;
      RECT 4.06 0.43 4.065 1.01 ;
      RECT 4.005 0.455 4.015 1.01 ;
      RECT 3.96 0.455 3.97 1.01 ;
      RECT 4.33 0.38 4.375 0.66 ;
      RECT 3.18 0.11 3.38 0.25 ;
      RECT 4.296 0.38 4.33 0.672 ;
      RECT 4.21 0.38 4.296 0.712 ;
      RECT 4.195 0.38 4.21 0.753 ;
      RECT 4.19 0.38 4.195 0.773 ;
      RECT 4.185 0.38 4.19 0.793 ;
      RECT 4.065 0.422 4.095 1.01 ;
      RECT 4.015 0.442 4.06 1.01 ;
      RECT 4 0.457 4.005 1.01 ;
      RECT 3.97 0.457 4 1.01 ;
      RECT 3.925 0.442 3.96 1.01 ;
      RECT 3.92 0.43 3.925 0.79 ;
      RECT 3.915 0.427 3.92 0.77 ;
      RECT 3.9 0.417 3.915 0.723 ;
      RECT 3.895 0.41 3.9 0.686 ;
      RECT 3.89 0.407 3.895 0.669 ;
      RECT 3.875 0.397 3.89 0.625 ;
      RECT 3.87 0.388 3.875 0.585 ;
      RECT 3.865 0.384 3.87 0.57 ;
      RECT 3.855 0.378 3.865 0.553 ;
      RECT 3.815 0.359 3.855 0.528 ;
      RECT 3.81 0.341 3.815 0.508 ;
      RECT 3.8 0.335 3.81 0.503 ;
      RECT 3.77 0.319 3.8 0.49 ;
      RECT 3.755 0.301 3.77 0.473 ;
      RECT 3.74 0.289 3.755 0.46 ;
      RECT 3.735 0.281 3.74 0.453 ;
      RECT 3.705 0.267 3.735 0.44 ;
      RECT 3.7 0.252 3.705 0.428 ;
      RECT 3.69 0.246 3.7 0.42 ;
      RECT 3.67 0.234 3.69 0.408 ;
      RECT 3.66 0.222 3.67 0.395 ;
      RECT 3.63 0.206 3.66 0.38 ;
      RECT 3.61 0.186 3.63 0.363 ;
      RECT 3.605 0.176 3.61 0.353 ;
      RECT 3.58 0.164 3.605 0.34 ;
      RECT 3.575 0.152 3.58 0.328 ;
      RECT 3.57 0.147 3.575 0.324 ;
      RECT 3.555 0.14 3.57 0.316 ;
      RECT 3.545 0.127 3.555 0.306 ;
      RECT 3.54 0.125 3.545 0.3 ;
      RECT 3.515 0.118 3.54 0.289 ;
      RECT 3.51 0.111 3.515 0.278 ;
      RECT 3.485 0.11 3.51 0.265 ;
      RECT 3.466 0.11 3.485 0.255 ;
      RECT 3.38 0.11 3.466 0.252 ;
      RECT 3.15 0.11 3.18 0.255 ;
      RECT 3.11 0.117 3.15 0.268 ;
      RECT 3.085 0.127 3.11 0.281 ;
      RECT 3.07 0.136 3.085 0.291 ;
      RECT 3.04 0.141 3.07 0.31 ;
      RECT 3.035 0.147 3.04 0.328 ;
      RECT 3.015 0.157 3.035 0.343 ;
      RECT 3.005 0.17 3.015 0.363 ;
      RECT 2.99 0.182 3.005 0.38 ;
      RECT 2.985 0.192 2.99 0.39 ;
      RECT 2.98 0.197 2.985 0.395 ;
      RECT 2.97 0.205 2.98 0.408 ;
      RECT 2.92 0.237 2.97 0.445 ;
      RECT 2.905 0.272 2.92 0.486 ;
      RECT 2.9 0.282 2.905 0.501 ;
      RECT 2.895 0.287 2.9 0.508 ;
      RECT 2.87 0.303 2.895 0.528 ;
      RECT 2.855 0.324 2.87 0.553 ;
      RECT 2.83 0.345 2.855 0.578 ;
      RECT 2.82 0.364 2.83 0.601 ;
      RECT 2.795 0.382 2.82 0.624 ;
      RECT 2.78 0.402 2.795 0.648 ;
      RECT 2.775 0.412 2.78 0.66 ;
      RECT 2.76 0.424 2.775 0.68 ;
      RECT 2.75 0.439 2.76 0.72 ;
      RECT 2.745 0.447 2.75 0.748 ;
      RECT 2.735 0.457 2.745 0.768 ;
      RECT 2.73 0.47 2.735 0.793 ;
      RECT 2.725 0.483 2.73 0.813 ;
      RECT 2.72 0.489 2.725 0.835 ;
      RECT 2.71 0.498 2.72 0.855 ;
      RECT 2.705 0.518 2.71 0.878 ;
      RECT 2.7 0.524 2.705 0.898 ;
      RECT 2.695 0.531 2.7 0.92 ;
      RECT 2.69 0.542 2.695 0.933 ;
      RECT 2.68 0.552 2.69 0.958 ;
      RECT 2.66 0.577 2.68 1.14 ;
      RECT 2.63 0.617 2.66 1.14 ;
      RECT 2.625 0.647 2.63 1.14 ;
      RECT 2.6 0.675 2.62 1.14 ;
      RECT 2.57 0.72 2.6 1.14 ;
      RECT 2.565 0.747 2.57 1.14 ;
      RECT 2.545 0.765 2.565 1.14 ;
      RECT 2.535 0.79 2.545 1.14 ;
      RECT 2.53 0.802 2.535 1.14 ;
      RECT 2.515 0.825 2.53 1.14 ;
      RECT 2.495 0.852 2.51 1.14 ;
      RECT 2.485 0.875 2.495 1.14 ;
      RECT 4.275 1.76 4.355 2.02 ;
      RECT 3.51 0.98 3.58 1.24 ;
      RECT 4.241 1.727 4.275 2.02 ;
      RECT 4.155 1.63 4.241 2.02 ;
      RECT 4.135 1.542 4.155 2.02 ;
      RECT 4.125 1.512 4.135 2.02 ;
      RECT 4.115 1.492 4.125 2.02 ;
      RECT 4.095 1.479 4.115 2.02 ;
      RECT 4.08 1.469 4.095 1.848 ;
      RECT 4.075 1.462 4.08 1.803 ;
      RECT 4.065 1.456 4.075 1.793 ;
      RECT 4.055 1.448 4.065 1.775 ;
      RECT 4.05 1.442 4.055 1.763 ;
      RECT 4.04 1.437 4.05 1.75 ;
      RECT 4.02 1.427 4.04 1.723 ;
      RECT 3.98 1.406 4.02 1.675 ;
      RECT 3.965 1.387 3.98 1.633 ;
      RECT 3.94 1.373 3.965 1.603 ;
      RECT 3.93 1.361 3.94 1.57 ;
      RECT 3.925 1.356 3.93 1.56 ;
      RECT 3.895 1.342 3.925 1.54 ;
      RECT 3.885 1.326 3.895 1.513 ;
      RECT 3.88 1.321 3.885 1.503 ;
      RECT 3.855 1.312 3.88 1.483 ;
      RECT 3.845 1.3 3.855 1.463 ;
      RECT 3.775 1.268 3.845 1.438 ;
      RECT 3.77 1.237 3.775 1.415 ;
      RECT 3.721 0.98 3.77 1.398 ;
      RECT 3.635 0.98 3.721 1.357 ;
      RECT 3.58 0.98 3.635 1.285 ;
      RECT 3.67 1.765 3.83 2.025 ;
      RECT 3.195 0.38 3.245 1.065 ;
      RECT 2.985 0.805 3.02 1.065 ;
      RECT 3.3 0.38 3.305 0.84 ;
      RECT 3.39 0.38 3.415 0.66 ;
      RECT 3.665 1.762 3.67 2.025 ;
      RECT 3.63 1.75 3.665 2.025 ;
      RECT 3.57 1.723 3.63 2.025 ;
      RECT 3.565 1.706 3.57 1.879 ;
      RECT 3.56 1.703 3.565 1.866 ;
      RECT 3.54 1.696 3.56 1.853 ;
      RECT 3.505 1.679 3.54 1.835 ;
      RECT 3.465 1.658 3.505 1.815 ;
      RECT 3.46 1.646 3.465 1.803 ;
      RECT 3.42 1.632 3.46 1.789 ;
      RECT 3.4 1.615 3.42 1.771 ;
      RECT 3.39 1.607 3.4 1.763 ;
      RECT 3.375 0.38 3.39 0.678 ;
      RECT 3.36 1.597 3.39 1.75 ;
      RECT 3.345 0.38 3.375 0.723 ;
      RECT 3.35 1.587 3.36 1.737 ;
      RECT 3.32 1.572 3.35 1.724 ;
      RECT 3.305 0.38 3.345 0.79 ;
      RECT 3.305 1.54 3.32 1.71 ;
      RECT 3.3 1.512 3.305 1.704 ;
      RECT 3.295 0.38 3.3 0.845 ;
      RECT 3.285 1.482 3.3 1.698 ;
      RECT 3.29 0.38 3.295 0.858 ;
      RECT 3.28 0.38 3.29 0.878 ;
      RECT 3.245 1.395 3.285 1.683 ;
      RECT 3.245 0.38 3.28 0.918 ;
      RECT 3.24 1.327 3.245 1.671 ;
      RECT 3.225 1.282 3.24 1.666 ;
      RECT 3.22 1.22 3.225 1.661 ;
      RECT 3.195 1.127 3.22 1.654 ;
      RECT 3.19 0.38 3.195 1.646 ;
      RECT 3.175 0.38 3.19 1.633 ;
      RECT 3.155 0.38 3.175 1.59 ;
      RECT 3.145 0.38 3.155 1.54 ;
      RECT 3.14 0.38 3.145 1.513 ;
      RECT 3.135 0.38 3.14 1.491 ;
      RECT 3.13 0.606 3.135 1.474 ;
      RECT 3.125 0.628 3.13 1.452 ;
      RECT 3.12 0.67 3.125 1.435 ;
      RECT 3.09 0.72 3.12 1.379 ;
      RECT 3.085 0.747 3.09 1.321 ;
      RECT 3.07 0.765 3.085 1.285 ;
      RECT 3.065 0.783 3.07 1.249 ;
      RECT 3.059 0.79 3.065 1.23 ;
      RECT 3.055 0.797 3.059 1.213 ;
      RECT 3.05 0.802 3.055 1.182 ;
      RECT 3.04 0.805 3.05 1.157 ;
      RECT 3.03 0.805 3.04 1.123 ;
      RECT 3.025 0.805 3.03 1.1 ;
      RECT 3.02 0.805 3.025 1.08 ;
      RECT 1.935 0.94 2.215 1.22 ;
      RECT 1.935 0.94 2.235 1.115 ;
      RECT 2.025 0.83 2.285 1.09 ;
      RECT 1.99 0.925 2.285 1.09 ;
      RECT 1.64 1.97 1.9 2.23 ;
      RECT 1.66 1.897 1.84 2.23 ;
      RECT 1.66 1.64 1.835 2.23 ;
      RECT 1.66 1.432 1.825 2.23 ;
      RECT 1.665 1.35 1.825 2.23 ;
      RECT 1.665 1.115 1.815 2.23 ;
      RECT 1.665 0.962 1.81 2.23 ;
      RECT 1.67 0.947 1.81 2.23 ;
      RECT 1.72 0.662 1.81 2.23 ;
      RECT 1.675 0.897 1.81 2.23 ;
      RECT 1.705 0.715 1.81 2.23 ;
      RECT 1.69 0.827 1.81 2.23 ;
      RECT 1.695 0.785 1.81 2.23 ;
      RECT 1.69 0.827 1.825 0.89 ;
      RECT 1.725 0.415 1.83 0.835 ;
      RECT 1.725 0.415 1.845 0.818 ;
      RECT 1.725 0.415 1.88 0.78 ;
      RECT 1.72 0.662 1.93 0.713 ;
      RECT 1.725 0.415 1.985 0.675 ;
      RECT 0.985 1.12 1.245 1.38 ;
      RECT 0.985 1.12 1.255 1.338 ;
      RECT 0.985 1.12 1.341 1.309 ;
      RECT 0.985 1.12 1.41 1.261 ;
      RECT 0.985 1.12 1.445 1.23 ;
      RECT 1.215 0.94 1.495 1.22 ;
      RECT 1.05 1.105 1.495 1.22 ;
      RECT 1.14 0.982 1.245 1.38 ;
      RECT 1.07 1.045 1.495 1.22 ;
    LAYER via1 ;
      RECT 7.505 0.85 7.655 1 ;
      RECT 6.485 1.555 6.635 1.705 ;
      RECT 6.255 0.975 6.405 1.125 ;
      RECT 5.91 1.575 6.06 1.725 ;
      RECT 5.67 0.595 5.82 0.745 ;
      RECT 5.36 1.925 5.51 2.075 ;
      RECT 5.22 0.53 5.37 0.68 ;
      RECT 4.585 0.615 4.735 0.765 ;
      RECT 4.475 1.255 4.625 1.405 ;
      RECT 4.15 1.815 4.3 1.965 ;
      RECT 3.98 0.805 4.13 0.955 ;
      RECT 3.625 1.82 3.775 1.97 ;
      RECT 3.565 1.035 3.715 1.185 ;
      RECT 3.2 2.025 3.35 2.175 ;
      RECT 3.04 0.86 3.19 1.01 ;
      RECT 2.475 0.935 2.625 1.085 ;
      RECT 2.08 0.885 2.23 1.035 ;
      RECT 1.78 0.47 1.93 0.62 ;
      RECT 1.695 2.025 1.845 2.175 ;
      RECT 1.04 1.175 1.19 1.325 ;
    LAYER met1 ;
      RECT 6.47 1.485 6.62 1.76 ;
      RECT 7.01 0.565 7.015 0.785 ;
      RECT 8.16 0.765 8.175 0.963 ;
      RECT 8.125 0.757 8.16 0.97 ;
      RECT 8.095 0.75 8.125 0.97 ;
      RECT 8.04 0.715 8.095 0.97 ;
      RECT 7.975 0.652 8.04 0.97 ;
      RECT 7.97 0.617 7.975 0.968 ;
      RECT 7.965 0.612 7.97 0.96 ;
      RECT 7.96 0.607 7.965 0.946 ;
      RECT 7.955 0.604 7.96 0.939 ;
      RECT 7.91 0.594 7.955 0.89 ;
      RECT 7.89 0.581 7.91 0.825 ;
      RECT 7.885 0.576 7.89 0.798 ;
      RECT 7.88 0.575 7.885 0.791 ;
      RECT 7.875 0.574 7.88 0.784 ;
      RECT 7.79 0.559 7.875 0.73 ;
      RECT 7.76 0.54 7.79 0.68 ;
      RECT 7.68 0.523 7.76 0.665 ;
      RECT 7.645 0.51 7.68 0.65 ;
      RECT 7.637 0.51 7.645 0.645 ;
      RECT 7.551 0.511 7.637 0.645 ;
      RECT 7.465 0.513 7.551 0.645 ;
      RECT 7.44 0.514 7.465 0.649 ;
      RECT 7.365 0.52 7.44 0.664 ;
      RECT 7.282 0.532 7.365 0.688 ;
      RECT 7.196 0.545 7.282 0.714 ;
      RECT 7.11 0.558 7.196 0.74 ;
      RECT 7.075 0.567 7.11 0.759 ;
      RECT 7.025 0.567 7.075 0.772 ;
      RECT 7.015 0.565 7.025 0.783 ;
      RECT 7 0.562 7.01 0.785 ;
      RECT 6.985 0.554 7 0.793 ;
      RECT 6.97 0.546 6.985 0.813 ;
      RECT 6.965 0.541 6.97 0.87 ;
      RECT 6.95 0.536 6.965 0.943 ;
      RECT 6.945 0.531 6.95 0.985 ;
      RECT 6.94 0.529 6.945 1.013 ;
      RECT 6.935 0.527 6.94 1.035 ;
      RECT 6.925 0.523 6.935 1.078 ;
      RECT 6.92 0.52 6.925 1.103 ;
      RECT 6.915 0.518 6.92 1.123 ;
      RECT 6.91 0.516 6.915 1.147 ;
      RECT 6.905 0.512 6.91 1.17 ;
      RECT 6.9 0.508 6.905 1.193 ;
      RECT 6.865 0.498 6.9 1.3 ;
      RECT 6.86 0.488 6.865 1.398 ;
      RECT 6.855 0.486 6.86 1.425 ;
      RECT 6.85 0.485 6.855 1.445 ;
      RECT 6.845 0.477 6.85 1.465 ;
      RECT 6.84 0.472 6.845 1.5 ;
      RECT 6.835 0.47 6.84 1.518 ;
      RECT 6.83 0.47 6.835 1.543 ;
      RECT 6.825 0.47 6.83 1.565 ;
      RECT 6.79 0.47 6.825 1.608 ;
      RECT 6.765 0.47 6.79 1.637 ;
      RECT 6.755 0.47 6.765 0.823 ;
      RECT 6.758 0.88 6.765 1.647 ;
      RECT 6.755 0.937 6.758 1.65 ;
      RECT 6.75 0.47 6.755 0.795 ;
      RECT 6.75 0.987 6.755 1.653 ;
      RECT 6.74 0.47 6.75 0.785 ;
      RECT 6.745 1.04 6.75 1.656 ;
      RECT 6.74 1.125 6.745 1.66 ;
      RECT 6.73 0.47 6.74 0.773 ;
      RECT 6.735 1.172 6.74 1.664 ;
      RECT 6.73 1.247 6.735 1.668 ;
      RECT 6.695 0.47 6.73 0.748 ;
      RECT 6.72 1.33 6.73 1.673 ;
      RECT 6.71 1.397 6.72 1.68 ;
      RECT 6.705 1.425 6.71 1.685 ;
      RECT 6.695 1.438 6.705 1.691 ;
      RECT 6.65 0.47 6.695 0.705 ;
      RECT 6.69 1.443 6.695 1.698 ;
      RECT 6.65 1.46 6.69 1.76 ;
      RECT 6.645 0.472 6.65 0.678 ;
      RECT 6.62 1.48 6.65 1.76 ;
      RECT 6.64 0.477 6.645 0.65 ;
      RECT 6.43 1.489 6.47 1.76 ;
      RECT 6.405 1.497 6.43 1.73 ;
      RECT 6.36 1.505 6.405 1.73 ;
      RECT 6.345 1.51 6.36 1.725 ;
      RECT 6.335 1.51 6.345 1.719 ;
      RECT 6.325 1.517 6.335 1.716 ;
      RECT 6.32 1.555 6.325 1.705 ;
      RECT 6.315 1.617 6.32 1.683 ;
      RECT 7.585 1.492 7.77 1.715 ;
      RECT 7.575 1.492 7.77 1.71 ;
      RECT 7.575 1.51 7.78 1.708 ;
      RECT 7.57 1.515 7.78 1.703 ;
      RECT 7.57 1.407 7.74 1.498 ;
      RECT 7.565 1.407 7.74 1.48 ;
      RECT 7.555 1.215 7.69 1.455 ;
      RECT 7.55 1.215 7.69 1.4 ;
      RECT 7.51 0.795 7.68 1.3 ;
      RECT 7.495 0.795 7.68 1.17 ;
      RECT 7.49 0.795 7.68 1.123 ;
      RECT 7.485 0.795 7.68 1.103 ;
      RECT 7.48 0.795 7.68 1.078 ;
      RECT 7.45 0.795 7.71 1.055 ;
      RECT 7.46 0.792 7.67 1.055 ;
      RECT 7.585 0.787 7.67 1.715 ;
      RECT 7.47 0.78 7.66 1.055 ;
      RECT 7.465 0.785 7.66 1.055 ;
      RECT 6.295 0.997 6.48 1.21 ;
      RECT 6.295 1.005 6.49 1.203 ;
      RECT 6.275 1.005 6.49 1.2 ;
      RECT 6.27 1.005 6.49 1.185 ;
      RECT 6.2 0.92 6.46 1.18 ;
      RECT 6.2 1.065 6.495 1.093 ;
      RECT 5.855 1.52 6.115 1.78 ;
      RECT 5.88 1.465 6.075 1.78 ;
      RECT 5.875 1.214 6.055 1.508 ;
      RECT 5.875 1.22 6.065 1.508 ;
      RECT 5.855 1.222 6.065 1.453 ;
      RECT 5.85 1.232 6.065 1.32 ;
      RECT 5.88 1.212 6.055 1.78 ;
      RECT 5.966 1.21 6.055 1.78 ;
      RECT 5.825 0.43 5.86 0.8 ;
      RECT 5.615 0.54 5.62 0.8 ;
      RECT 5.86 0.437 5.875 0.8 ;
      RECT 5.75 0.43 5.825 0.878 ;
      RECT 5.74 0.43 5.75 0.963 ;
      RECT 5.715 0.43 5.74 0.998 ;
      RECT 5.675 0.43 5.715 1.066 ;
      RECT 5.665 0.437 5.675 1.118 ;
      RECT 5.635 0.54 5.665 1.159 ;
      RECT 5.63 0.54 5.635 1.198 ;
      RECT 5.62 0.54 5.63 1.218 ;
      RECT 5.615 0.835 5.62 1.255 ;
      RECT 5.61 0.852 5.615 1.275 ;
      RECT 5.595 0.915 5.61 1.315 ;
      RECT 5.59 0.958 5.595 1.35 ;
      RECT 5.585 0.966 5.59 1.363 ;
      RECT 5.575 0.98 5.585 1.385 ;
      RECT 5.55 1.015 5.575 1.45 ;
      RECT 5.54 1.05 5.55 1.513 ;
      RECT 5.52 1.08 5.54 1.574 ;
      RECT 5.505 1.116 5.52 1.641 ;
      RECT 5.495 1.144 5.505 1.68 ;
      RECT 5.485 1.166 5.495 1.7 ;
      RECT 5.48 1.176 5.485 1.711 ;
      RECT 5.475 1.185 5.48 1.714 ;
      RECT 5.465 1.203 5.475 1.718 ;
      RECT 5.455 1.221 5.465 1.719 ;
      RECT 5.43 1.26 5.455 1.716 ;
      RECT 5.41 1.302 5.43 1.713 ;
      RECT 5.395 1.34 5.41 1.712 ;
      RECT 5.36 1.375 5.395 1.709 ;
      RECT 5.355 1.397 5.36 1.707 ;
      RECT 5.29 1.437 5.355 1.704 ;
      RECT 5.285 1.477 5.29 1.7 ;
      RECT 5.27 1.487 5.285 1.691 ;
      RECT 5.26 1.607 5.27 1.676 ;
      RECT 5.74 2.02 5.75 2.28 ;
      RECT 5.74 2.023 5.76 2.279 ;
      RECT 5.73 2.013 5.74 2.278 ;
      RECT 5.72 2.028 5.8 2.274 ;
      RECT 5.705 2.007 5.72 2.272 ;
      RECT 5.68 2.032 5.805 2.268 ;
      RECT 5.665 1.992 5.68 2.263 ;
      RECT 5.665 2.034 5.815 2.262 ;
      RECT 5.665 2.042 5.83 2.255 ;
      RECT 5.605 1.979 5.665 2.245 ;
      RECT 5.595 1.966 5.605 2.227 ;
      RECT 5.57 1.956 5.595 2.217 ;
      RECT 5.565 1.946 5.57 2.209 ;
      RECT 5.5 2.042 5.83 2.191 ;
      RECT 5.415 2.042 5.83 2.153 ;
      RECT 5.305 1.87 5.565 2.13 ;
      RECT 5.68 2 5.705 2.268 ;
      RECT 5.72 2.01 5.73 2.274 ;
      RECT 5.305 2.018 5.745 2.13 ;
      RECT 4.52 1.775 4.55 2.075 ;
      RECT 4.295 1.76 4.3 2.035 ;
      RECT 4.095 1.76 4.25 2.02 ;
      RECT 5.395 0.475 5.425 0.735 ;
      RECT 5.385 0.475 5.395 0.843 ;
      RECT 5.365 0.475 5.385 0.853 ;
      RECT 5.35 0.475 5.365 0.865 ;
      RECT 5.295 0.475 5.35 0.915 ;
      RECT 5.28 0.475 5.295 0.963 ;
      RECT 5.25 0.475 5.28 0.998 ;
      RECT 5.195 0.475 5.25 1.06 ;
      RECT 5.175 0.475 5.195 1.128 ;
      RECT 5.17 0.475 5.175 1.158 ;
      RECT 5.165 0.475 5.17 1.17 ;
      RECT 5.16 0.592 5.165 1.188 ;
      RECT 5.14 0.61 5.16 1.213 ;
      RECT 5.12 0.637 5.14 1.263 ;
      RECT 5.115 0.657 5.12 1.294 ;
      RECT 5.11 0.665 5.115 1.311 ;
      RECT 5.095 0.691 5.11 1.34 ;
      RECT 5.08 0.733 5.095 1.375 ;
      RECT 5.075 0.762 5.08 1.398 ;
      RECT 5.07 0.777 5.075 1.411 ;
      RECT 5.065 0.8 5.07 1.422 ;
      RECT 5.055 0.82 5.065 1.44 ;
      RECT 5.045 0.85 5.055 1.463 ;
      RECT 5.04 0.872 5.045 1.483 ;
      RECT 5.035 0.887 5.04 1.498 ;
      RECT 5.02 0.917 5.035 1.525 ;
      RECT 5.015 0.947 5.02 1.551 ;
      RECT 5.01 0.965 5.015 1.563 ;
      RECT 5 0.995 5.01 1.582 ;
      RECT 4.99 1.02 5 1.607 ;
      RECT 4.985 1.04 4.99 1.626 ;
      RECT 4.98 1.057 4.985 1.639 ;
      RECT 4.97 1.083 4.98 1.658 ;
      RECT 4.96 1.121 4.97 1.685 ;
      RECT 4.955 1.147 4.96 1.705 ;
      RECT 4.95 1.157 4.955 1.715 ;
      RECT 4.945 1.17 4.95 1.73 ;
      RECT 4.94 1.185 4.945 1.74 ;
      RECT 4.935 1.207 4.94 1.755 ;
      RECT 4.93 1.225 4.935 1.766 ;
      RECT 4.925 1.235 4.93 1.777 ;
      RECT 4.92 1.243 4.925 1.789 ;
      RECT 4.915 1.251 4.92 1.8 ;
      RECT 4.91 1.277 4.915 1.813 ;
      RECT 4.9 1.305 4.91 1.826 ;
      RECT 4.895 1.335 4.9 1.835 ;
      RECT 4.89 1.35 4.895 1.842 ;
      RECT 4.875 1.375 4.89 1.849 ;
      RECT 4.87 1.397 4.875 1.855 ;
      RECT 4.865 1.422 4.87 1.858 ;
      RECT 4.856 1.45 4.865 1.862 ;
      RECT 4.85 1.467 4.856 1.867 ;
      RECT 4.845 1.485 4.85 1.871 ;
      RECT 4.84 1.497 4.845 1.874 ;
      RECT 4.835 1.518 4.84 1.878 ;
      RECT 4.83 1.536 4.835 1.881 ;
      RECT 4.825 1.55 4.83 1.884 ;
      RECT 4.82 1.567 4.825 1.887 ;
      RECT 4.815 1.58 4.82 1.89 ;
      RECT 4.79 1.617 4.815 1.898 ;
      RECT 4.785 1.662 4.79 1.907 ;
      RECT 4.78 1.69 4.785 1.91 ;
      RECT 4.77 1.71 4.78 1.914 ;
      RECT 4.765 1.73 4.77 1.919 ;
      RECT 4.76 1.745 4.765 1.922 ;
      RECT 4.74 1.755 4.76 1.929 ;
      RECT 4.675 1.762 4.74 1.955 ;
      RECT 4.64 1.765 4.675 1.983 ;
      RECT 4.625 1.768 4.64 1.998 ;
      RECT 4.615 1.769 4.625 2.013 ;
      RECT 4.605 1.77 4.615 2.03 ;
      RECT 4.6 1.77 4.605 2.045 ;
      RECT 4.595 1.77 4.6 2.053 ;
      RECT 4.58 1.771 4.595 2.068 ;
      RECT 4.55 1.773 4.58 2.075 ;
      RECT 4.44 1.78 4.52 2.075 ;
      RECT 4.395 1.785 4.44 2.075 ;
      RECT 4.385 1.786 4.395 2.065 ;
      RECT 4.375 1.787 4.385 2.058 ;
      RECT 4.355 1.789 4.375 2.053 ;
      RECT 4.345 1.76 4.355 2.048 ;
      RECT 4.3 1.76 4.345 2.04 ;
      RECT 4.27 1.76 4.295 2.03 ;
      RECT 4.25 1.76 4.27 2.023 ;
      RECT 4.53 0.56 4.79 0.82 ;
      RECT 4.41 0.575 4.42 0.74 ;
      RECT 4.395 0.575 4.4 0.735 ;
      RECT 1.76 0.415 1.945 0.705 ;
      RECT 3.575 0.54 3.59 0.695 ;
      RECT 1.725 0.415 1.75 0.675 ;
      RECT 4.14 0.465 4.145 0.607 ;
      RECT 4.055 0.46 4.08 0.6 ;
      RECT 4.455 0.577 4.53 0.77 ;
      RECT 4.44 0.575 4.455 0.753 ;
      RECT 4.42 0.575 4.44 0.745 ;
      RECT 4.4 0.575 4.41 0.738 ;
      RECT 4.355 0.57 4.395 0.728 ;
      RECT 4.315 0.545 4.355 0.713 ;
      RECT 4.3 0.52 4.315 0.703 ;
      RECT 4.295 0.514 4.3 0.701 ;
      RECT 4.26 0.506 4.295 0.684 ;
      RECT 4.255 0.499 4.26 0.672 ;
      RECT 4.235 0.494 4.255 0.66 ;
      RECT 4.225 0.488 4.235 0.645 ;
      RECT 4.205 0.483 4.225 0.63 ;
      RECT 4.195 0.478 4.205 0.623 ;
      RECT 4.19 0.476 4.195 0.618 ;
      RECT 4.185 0.475 4.19 0.615 ;
      RECT 4.145 0.47 4.185 0.611 ;
      RECT 4.125 0.464 4.14 0.606 ;
      RECT 4.09 0.461 4.125 0.603 ;
      RECT 4.08 0.46 4.09 0.601 ;
      RECT 4.02 0.46 4.055 0.598 ;
      RECT 3.975 0.46 4.02 0.598 ;
      RECT 3.925 0.46 3.975 0.601 ;
      RECT 3.91 0.462 3.925 0.603 ;
      RECT 3.895 0.465 3.91 0.604 ;
      RECT 3.885 0.47 3.895 0.605 ;
      RECT 3.855 0.475 3.885 0.61 ;
      RECT 3.845 0.481 3.855 0.618 ;
      RECT 3.835 0.483 3.845 0.622 ;
      RECT 3.825 0.487 3.835 0.626 ;
      RECT 3.8 0.493 3.825 0.634 ;
      RECT 3.79 0.498 3.8 0.642 ;
      RECT 3.775 0.502 3.79 0.646 ;
      RECT 3.74 0.508 3.775 0.654 ;
      RECT 3.72 0.513 3.74 0.664 ;
      RECT 3.69 0.52 3.72 0.673 ;
      RECT 3.645 0.529 3.69 0.687 ;
      RECT 3.64 0.534 3.645 0.698 ;
      RECT 3.62 0.537 3.64 0.699 ;
      RECT 3.59 0.54 3.62 0.697 ;
      RECT 3.555 0.54 3.575 0.693 ;
      RECT 3.485 0.54 3.555 0.684 ;
      RECT 3.47 0.537 3.485 0.676 ;
      RECT 3.43 0.53 3.47 0.671 ;
      RECT 3.405 0.52 3.43 0.664 ;
      RECT 3.4 0.514 3.405 0.661 ;
      RECT 3.36 0.508 3.4 0.658 ;
      RECT 3.345 0.501 3.36 0.653 ;
      RECT 3.325 0.497 3.345 0.648 ;
      RECT 3.31 0.492 3.325 0.644 ;
      RECT 3.295 0.487 3.31 0.642 ;
      RECT 3.28 0.483 3.295 0.641 ;
      RECT 3.265 0.481 3.28 0.637 ;
      RECT 3.255 0.479 3.265 0.632 ;
      RECT 3.24 0.476 3.255 0.628 ;
      RECT 3.23 0.474 3.24 0.623 ;
      RECT 3.21 0.471 3.23 0.619 ;
      RECT 3.165 0.47 3.21 0.617 ;
      RECT 3.105 0.472 3.165 0.618 ;
      RECT 3.085 0.474 3.105 0.62 ;
      RECT 3.055 0.477 3.085 0.621 ;
      RECT 3.005 0.482 3.055 0.623 ;
      RECT 3 0.485 3.005 0.625 ;
      RECT 2.99 0.487 3 0.628 ;
      RECT 2.985 0.489 2.99 0.631 ;
      RECT 2.935 0.492 2.985 0.638 ;
      RECT 2.915 0.496 2.935 0.65 ;
      RECT 2.905 0.499 2.915 0.656 ;
      RECT 2.895 0.5 2.905 0.659 ;
      RECT 2.856 0.503 2.895 0.661 ;
      RECT 2.77 0.51 2.856 0.664 ;
      RECT 2.696 0.52 2.77 0.668 ;
      RECT 2.61 0.531 2.696 0.673 ;
      RECT 2.595 0.538 2.61 0.675 ;
      RECT 2.54 0.542 2.595 0.676 ;
      RECT 2.526 0.545 2.54 0.678 ;
      RECT 2.44 0.545 2.526 0.68 ;
      RECT 2.4 0.542 2.44 0.683 ;
      RECT 2.376 0.538 2.4 0.685 ;
      RECT 2.29 0.528 2.376 0.688 ;
      RECT 2.26 0.517 2.29 0.689 ;
      RECT 2.241 0.513 2.26 0.688 ;
      RECT 2.155 0.506 2.241 0.685 ;
      RECT 2.095 0.495 2.155 0.682 ;
      RECT 2.075 0.487 2.095 0.68 ;
      RECT 2.04 0.482 2.075 0.679 ;
      RECT 2.015 0.477 2.04 0.678 ;
      RECT 1.985 0.472 2.015 0.677 ;
      RECT 1.96 0.415 1.985 0.676 ;
      RECT 1.945 0.415 1.96 0.7 ;
      RECT 1.75 0.415 1.76 0.7 ;
      RECT 3.525 1.435 3.53 1.575 ;
      RECT 3.185 1.435 3.22 1.573 ;
      RECT 2.76 1.42 2.775 1.565 ;
      RECT 4.59 1.2 4.68 1.46 ;
      RECT 4.42 1.065 4.52 1.46 ;
      RECT 1.455 1.04 1.535 1.25 ;
      RECT 4.545 1.177 4.59 1.46 ;
      RECT 4.535 1.147 4.545 1.46 ;
      RECT 4.52 1.07 4.535 1.46 ;
      RECT 4.335 1.065 4.42 1.425 ;
      RECT 4.33 1.067 4.335 1.42 ;
      RECT 4.325 1.072 4.33 1.42 ;
      RECT 4.29 1.172 4.325 1.42 ;
      RECT 4.28 1.2 4.29 1.42 ;
      RECT 4.27 1.215 4.28 1.42 ;
      RECT 4.26 1.227 4.27 1.42 ;
      RECT 4.255 1.237 4.26 1.42 ;
      RECT 4.24 1.247 4.255 1.422 ;
      RECT 4.235 1.262 4.24 1.424 ;
      RECT 4.22 1.275 4.235 1.426 ;
      RECT 4.215 1.29 4.22 1.429 ;
      RECT 4.195 1.3 4.215 1.433 ;
      RECT 4.18 1.31 4.195 1.436 ;
      RECT 4.145 1.317 4.18 1.441 ;
      RECT 4.101 1.324 4.145 1.449 ;
      RECT 4.015 1.336 4.101 1.462 ;
      RECT 3.99 1.347 4.015 1.473 ;
      RECT 3.96 1.352 3.99 1.478 ;
      RECT 3.925 1.357 3.96 1.486 ;
      RECT 3.895 1.362 3.925 1.493 ;
      RECT 3.87 1.367 3.895 1.498 ;
      RECT 3.805 1.374 3.87 1.507 ;
      RECT 3.735 1.387 3.805 1.523 ;
      RECT 3.705 1.397 3.735 1.535 ;
      RECT 3.68 1.402 3.705 1.542 ;
      RECT 3.625 1.409 3.68 1.55 ;
      RECT 3.62 1.416 3.625 1.555 ;
      RECT 3.615 1.418 3.62 1.556 ;
      RECT 3.6 1.42 3.615 1.558 ;
      RECT 3.595 1.42 3.6 1.561 ;
      RECT 3.53 1.427 3.595 1.568 ;
      RECT 3.495 1.437 3.525 1.578 ;
      RECT 3.478 1.44 3.495 1.58 ;
      RECT 3.392 1.439 3.478 1.579 ;
      RECT 3.306 1.437 3.392 1.576 ;
      RECT 3.22 1.436 3.306 1.574 ;
      RECT 3.119 1.434 3.185 1.573 ;
      RECT 3.033 1.431 3.119 1.571 ;
      RECT 2.947 1.427 3.033 1.569 ;
      RECT 2.861 1.424 2.947 1.568 ;
      RECT 2.775 1.421 2.861 1.566 ;
      RECT 2.675 1.42 2.76 1.563 ;
      RECT 2.625 1.418 2.675 1.561 ;
      RECT 2.605 1.415 2.625 1.559 ;
      RECT 2.585 1.413 2.605 1.556 ;
      RECT 2.56 1.409 2.585 1.553 ;
      RECT 2.515 1.403 2.56 1.548 ;
      RECT 2.475 1.397 2.515 1.54 ;
      RECT 2.45 1.392 2.475 1.533 ;
      RECT 2.395 1.385 2.45 1.525 ;
      RECT 2.371 1.378 2.395 1.518 ;
      RECT 2.285 1.369 2.371 1.508 ;
      RECT 2.255 1.361 2.285 1.498 ;
      RECT 2.225 1.357 2.255 1.493 ;
      RECT 2.22 1.354 2.225 1.49 ;
      RECT 2.215 1.353 2.22 1.49 ;
      RECT 2.14 1.346 2.215 1.483 ;
      RECT 2.101 1.337 2.14 1.472 ;
      RECT 2.015 1.327 2.101 1.46 ;
      RECT 1.975 1.317 2.015 1.448 ;
      RECT 1.936 1.312 1.975 1.441 ;
      RECT 1.85 1.302 1.936 1.43 ;
      RECT 1.81 1.29 1.85 1.419 ;
      RECT 1.775 1.275 1.81 1.412 ;
      RECT 1.765 1.265 1.775 1.409 ;
      RECT 1.745 1.25 1.765 1.407 ;
      RECT 1.715 1.22 1.745 1.403 ;
      RECT 1.705 1.2 1.715 1.398 ;
      RECT 1.7 1.192 1.705 1.395 ;
      RECT 1.695 1.185 1.7 1.393 ;
      RECT 1.68 1.172 1.695 1.386 ;
      RECT 1.675 1.162 1.68 1.378 ;
      RECT 1.67 1.155 1.675 1.373 ;
      RECT 1.665 1.15 1.67 1.369 ;
      RECT 1.65 1.137 1.665 1.361 ;
      RECT 1.645 1.047 1.65 1.35 ;
      RECT 1.64 1.042 1.645 1.343 ;
      RECT 1.565 1.04 1.64 1.303 ;
      RECT 1.535 1.04 1.565 1.258 ;
      RECT 1.44 1.045 1.455 1.245 ;
      RECT 3.925 0.75 4.185 1.01 ;
      RECT 3.91 0.738 4.09 0.975 ;
      RECT 3.905 0.739 4.09 0.973 ;
      RECT 3.89 0.743 4.1 0.963 ;
      RECT 3.885 0.748 4.105 0.933 ;
      RECT 3.89 0.745 4.105 0.963 ;
      RECT 3.905 0.74 4.1 0.973 ;
      RECT 3.925 0.737 4.09 1.01 ;
      RECT 3.925 0.736 4.08 1.01 ;
      RECT 3.95 0.735 4.08 1.01 ;
      RECT 3.51 0.98 3.77 1.24 ;
      RECT 3.385 1.025 3.77 1.235 ;
      RECT 3.375 1.03 3.77 1.23 ;
      RECT 3.39 1.97 3.405 2.28 ;
      RECT 1.985 1.74 1.995 1.87 ;
      RECT 1.765 1.735 1.87 1.87 ;
      RECT 1.68 1.74 1.73 1.87 ;
      RECT 0.23 0.475 0.235 1.58 ;
      RECT 3.485 2.062 3.49 2.198 ;
      RECT 3.48 2.057 3.485 2.258 ;
      RECT 3.475 2.055 3.48 2.271 ;
      RECT 3.46 2.052 3.475 2.273 ;
      RECT 3.455 2.047 3.46 2.275 ;
      RECT 3.45 2.043 3.455 2.278 ;
      RECT 3.435 2.038 3.45 2.28 ;
      RECT 3.405 2.03 3.435 2.28 ;
      RECT 3.366 1.97 3.39 2.28 ;
      RECT 3.28 1.97 3.366 2.277 ;
      RECT 3.25 1.97 3.28 2.27 ;
      RECT 3.225 1.97 3.25 2.263 ;
      RECT 3.2 1.97 3.225 2.255 ;
      RECT 3.185 1.97 3.2 2.248 ;
      RECT 3.16 1.97 3.185 2.24 ;
      RECT 3.145 1.97 3.16 2.233 ;
      RECT 3.105 1.98 3.145 2.222 ;
      RECT 3.095 1.975 3.105 2.212 ;
      RECT 3.091 1.974 3.095 2.209 ;
      RECT 3.005 1.966 3.091 2.192 ;
      RECT 2.972 1.955 3.005 2.169 ;
      RECT 2.886 1.944 2.972 2.147 ;
      RECT 2.8 1.928 2.886 2.116 ;
      RECT 2.73 1.913 2.8 2.088 ;
      RECT 2.72 1.906 2.73 2.075 ;
      RECT 2.69 1.903 2.72 2.065 ;
      RECT 2.665 1.899 2.69 2.058 ;
      RECT 2.65 1.896 2.665 2.053 ;
      RECT 2.645 1.895 2.65 2.048 ;
      RECT 2.615 1.89 2.645 2.041 ;
      RECT 2.61 1.885 2.615 2.036 ;
      RECT 2.595 1.882 2.61 2.031 ;
      RECT 2.59 1.877 2.595 2.026 ;
      RECT 2.57 1.872 2.59 2.023 ;
      RECT 2.555 1.867 2.57 2.015 ;
      RECT 2.54 1.861 2.555 2.01 ;
      RECT 2.51 1.852 2.54 2.003 ;
      RECT 2.505 1.845 2.51 1.995 ;
      RECT 2.5 1.843 2.505 1.993 ;
      RECT 2.495 1.842 2.5 1.99 ;
      RECT 2.455 1.835 2.495 1.983 ;
      RECT 2.441 1.825 2.455 1.973 ;
      RECT 2.39 1.814 2.441 1.961 ;
      RECT 2.365 1.8 2.39 1.947 ;
      RECT 2.34 1.789 2.365 1.939 ;
      RECT 2.32 1.778 2.34 1.933 ;
      RECT 2.31 1.772 2.32 1.928 ;
      RECT 2.305 1.77 2.31 1.924 ;
      RECT 2.285 1.765 2.305 1.919 ;
      RECT 2.255 1.755 2.285 1.909 ;
      RECT 2.25 1.747 2.255 1.902 ;
      RECT 2.235 1.745 2.25 1.898 ;
      RECT 2.215 1.745 2.235 1.893 ;
      RECT 2.21 1.744 2.215 1.891 ;
      RECT 2.205 1.744 2.21 1.888 ;
      RECT 2.165 1.743 2.205 1.883 ;
      RECT 2.14 1.742 2.165 1.878 ;
      RECT 2.08 1.741 2.14 1.875 ;
      RECT 1.995 1.74 2.08 1.873 ;
      RECT 1.956 1.739 1.985 1.87 ;
      RECT 1.87 1.737 1.956 1.87 ;
      RECT 1.73 1.737 1.765 1.87 ;
      RECT 1.64 1.741 1.68 1.873 ;
      RECT 1.625 1.744 1.64 1.88 ;
      RECT 1.615 1.745 1.625 1.887 ;
      RECT 1.59 1.748 1.615 1.892 ;
      RECT 1.585 1.75 1.59 1.895 ;
      RECT 1.535 1.752 1.585 1.896 ;
      RECT 1.496 1.756 1.535 1.898 ;
      RECT 1.41 1.758 1.496 1.901 ;
      RECT 1.392 1.76 1.41 1.903 ;
      RECT 1.306 1.763 1.392 1.905 ;
      RECT 1.22 1.767 1.306 1.908 ;
      RECT 1.183 1.771 1.22 1.911 ;
      RECT 1.097 1.774 1.183 1.914 ;
      RECT 1.011 1.778 1.097 1.917 ;
      RECT 0.925 1.783 1.011 1.921 ;
      RECT 0.905 1.785 0.925 1.924 ;
      RECT 0.885 1.784 0.905 1.925 ;
      RECT 0.836 1.781 0.885 1.926 ;
      RECT 0.75 1.776 0.836 1.929 ;
      RECT 0.7 1.771 0.75 1.931 ;
      RECT 0.676 1.769 0.7 1.932 ;
      RECT 0.59 1.764 0.676 1.934 ;
      RECT 0.565 1.76 0.59 1.933 ;
      RECT 0.555 1.757 0.565 1.931 ;
      RECT 0.545 1.75 0.555 1.928 ;
      RECT 0.54 1.73 0.545 1.923 ;
      RECT 0.53 1.7 0.54 1.918 ;
      RECT 0.515 1.57 0.53 1.909 ;
      RECT 0.51 1.562 0.515 1.902 ;
      RECT 0.49 1.555 0.51 1.894 ;
      RECT 0.485 1.537 0.49 1.886 ;
      RECT 0.475 1.517 0.485 1.881 ;
      RECT 0.47 1.49 0.475 1.877 ;
      RECT 0.465 1.467 0.47 1.874 ;
      RECT 0.445 1.425 0.465 1.866 ;
      RECT 0.41 1.34 0.445 1.85 ;
      RECT 0.405 1.272 0.41 1.838 ;
      RECT 0.39 1.242 0.405 1.832 ;
      RECT 0.385 0.487 0.39 0.733 ;
      RECT 0.375 1.212 0.39 1.823 ;
      RECT 0.38 0.482 0.385 0.765 ;
      RECT 0.375 0.477 0.38 0.808 ;
      RECT 0.37 0.475 0.375 0.843 ;
      RECT 0.355 1.175 0.375 1.813 ;
      RECT 0.365 0.475 0.37 0.88 ;
      RECT 0.35 0.475 0.365 0.978 ;
      RECT 0.35 1.148 0.355 1.806 ;
      RECT 0.345 0.475 0.35 1.053 ;
      RECT 0.345 1.136 0.35 1.803 ;
      RECT 0.34 0.475 0.345 1.085 ;
      RECT 0.34 1.115 0.345 1.8 ;
      RECT 0.335 0.475 0.34 1.797 ;
      RECT 0.3 0.475 0.335 1.783 ;
      RECT 0.285 0.475 0.3 1.765 ;
      RECT 0.265 0.475 0.285 1.755 ;
      RECT 0.24 0.475 0.265 1.738 ;
      RECT 0.235 0.475 0.24 1.688 ;
      RECT 0.225 0.475 0.23 1.518 ;
      RECT 0.22 0.475 0.225 1.425 ;
      RECT 0.215 0.475 0.22 1.338 ;
      RECT 0.21 0.475 0.215 1.27 ;
      RECT 0.205 0.475 0.21 1.213 ;
      RECT 0.195 0.475 0.205 1.108 ;
      RECT 0.19 0.475 0.195 0.98 ;
      RECT 0.185 0.475 0.19 0.898 ;
      RECT 0.18 0.477 0.185 0.815 ;
      RECT 0.175 0.482 0.18 0.748 ;
      RECT 0.17 0.487 0.175 0.675 ;
      RECT 2.985 0.805 3.245 1.065 ;
      RECT 3.005 0.772 3.215 1.065 ;
      RECT 3.005 0.77 3.205 1.065 ;
      RECT 3.015 0.757 3.205 1.065 ;
      RECT 3.015 0.755 3.13 1.065 ;
      RECT 2.49 0.88 2.665 1.16 ;
      RECT 2.485 0.88 2.665 1.158 ;
      RECT 2.485 0.88 2.68 1.155 ;
      RECT 2.475 0.88 2.68 1.153 ;
      RECT 2.42 0.88 2.68 1.14 ;
      RECT 2.42 0.955 2.685 1.118 ;
      RECT 1.965 0.892 1.985 1.135 ;
      RECT 1.965 0.892 2.025 1.134 ;
      RECT 1.96 0.894 2.025 1.133 ;
      RECT 1.96 0.894 2.111 1.132 ;
      RECT 1.96 0.894 2.18 1.131 ;
      RECT 1.96 0.894 2.2 1.123 ;
      RECT 1.94 0.897 2.2 1.121 ;
      RECT 1.925 0.907 2.2 1.106 ;
      RECT 1.925 0.907 2.215 1.105 ;
      RECT 1.92 0.916 2.215 1.097 ;
      RECT 1.92 0.916 2.22 1.093 ;
      RECT 2.025 0.83 2.285 1.09 ;
      RECT 1.915 0.918 2.285 0.975 ;
      RECT 1.985 0.885 2.285 1.09 ;
      RECT 1.95 2.078 1.955 2.285 ;
      RECT 1.9 2.072 1.95 2.284 ;
      RECT 1.867 2.086 1.96 2.283 ;
      RECT 1.781 2.086 1.96 2.282 ;
      RECT 1.695 2.086 1.96 2.281 ;
      RECT 1.695 2.185 1.965 2.278 ;
      RECT 1.69 2.185 1.965 2.273 ;
      RECT 1.685 2.185 1.965 2.255 ;
      RECT 1.68 2.185 1.965 2.238 ;
      RECT 1.64 1.97 1.9 2.23 ;
      RECT 1.1 1.12 1.186 1.534 ;
      RECT 1.1 1.12 1.225 1.531 ;
      RECT 1.1 1.12 1.245 1.521 ;
      RECT 1.055 1.12 1.245 1.518 ;
      RECT 1.055 1.272 1.255 1.508 ;
      RECT 1.055 1.293 1.26 1.502 ;
      RECT 1.055 1.311 1.265 1.498 ;
      RECT 1.055 1.331 1.275 1.493 ;
      RECT 1.03 1.331 1.275 1.49 ;
      RECT 1.02 1.331 1.275 1.468 ;
      RECT 1.02 1.347 1.28 1.438 ;
      RECT 0.985 1.12 1.245 1.425 ;
      RECT 0.985 1.359 1.285 1.38 ;
      RECT 0 -0.24 8.74 0.24 ;
      RECT 0 2.48 8.74 2.96 ;
      RECT 3.57 1.765 3.83 2.025 ;
    LAYER mcon ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 8.425 2.635 8.595 2.805 ;
      RECT 7.985 0.78 8.155 0.95 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.965 2.635 8.135 2.805 ;
      RECT 7.59 1.525 7.76 1.695 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.505 2.635 7.675 2.805 ;
      RECT 7.48 0.8 7.65 0.97 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 7.045 2.635 7.215 2.805 ;
      RECT 6.66 0.49 6.83 0.66 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.585 2.635 6.755 2.805 ;
      RECT 6.345 1.53 6.515 1.7 ;
      RECT 6.3 1.02 6.47 1.19 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 6.125 2.635 6.295 2.805 ;
      RECT 5.875 1.23 6.045 1.4 ;
      RECT 5.685 0.45 5.855 0.62 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.665 2.635 5.835 2.805 ;
      RECT 5.635 2.06 5.805 2.23 ;
      RECT 5.3 1.5 5.47 1.67 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 5.205 0.66 5.375 0.83 ;
      RECT 5.205 2.635 5.375 2.805 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.745 2.635 4.915 2.805 ;
      RECT 4.405 1.885 4.575 2.055 ;
      RECT 4.345 1.085 4.515 1.255 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 4.285 2.635 4.455 2.805 ;
      RECT 3.905 0.755 4.075 0.925 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.825 2.635 3.995 2.805 ;
      RECT 3.64 1.805 3.81 1.975 ;
      RECT 3.395 1.045 3.565 1.215 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 3.365 2.635 3.535 2.805 ;
      RECT 3.3 2.075 3.47 2.245 ;
      RECT 3.025 0.77 3.195 0.94 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.905 2.635 3.075 2.805 ;
      RECT 2.495 0.97 2.665 1.14 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 2.445 2.635 2.615 2.805 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.985 2.635 2.155 2.805 ;
      RECT 1.975 0.915 2.145 1.085 ;
      RECT 1.77 0.515 1.94 0.685 ;
      RECT 1.77 2.095 1.94 2.265 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.525 2.635 1.695 2.805 ;
      RECT 1.46 1.06 1.63 1.23 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 1.065 2.635 1.235 2.805 ;
      RECT 1.05 1.285 1.22 1.455 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.34 1.585 0.51 1.755 ;
      RECT 0.195 0.495 0.365 0.665 ;
      RECT 0.145 -0.085 0.315 0.085 ;
      RECT 0.145 2.635 0.315 2.805 ;
    LAYER li ;
      RECT 7.97 -0.085 8.14 0.585 ;
      RECT 7.03 -0.085 7.2 0.585 ;
      RECT 6.07 -0.085 6.24 0.585 ;
      RECT 4.15 -0.085 4.32 0.585 ;
      RECT 3.19 -0.085 3.36 0.585 ;
      RECT 1.27 -0.085 1.44 0.585 ;
      RECT 0 -0.085 8.74 0.085 ;
      RECT 0 2.635 8.74 2.805 ;
      RECT 7.03 2.135 7.2 2.805 ;
      RECT 5.11 2.135 5.28 2.805 ;
      RECT 4.17 2.135 4.34 2.805 ;
      RECT 2.71 2.135 2.88 2.805 ;
      RECT 0.79 2.135 0.96 2.805 ;
      RECT 8.16 1.626 8.165 1.798 ;
      RECT 8.155 1.619 8.16 1.888 ;
      RECT 8.15 1.613 8.155 1.907 ;
      RECT 8.13 1.607 8.15 1.917 ;
      RECT 8.115 1.602 8.13 1.925 ;
      RECT 8.078 1.596 8.115 1.923 ;
      RECT 7.992 1.582 8.078 1.919 ;
      RECT 7.906 1.564 7.992 1.914 ;
      RECT 7.82 1.545 7.906 1.908 ;
      RECT 7.79 1.533 7.82 1.904 ;
      RECT 7.77 1.527 7.79 1.903 ;
      RECT 7.705 1.525 7.77 1.901 ;
      RECT 7.69 1.525 7.705 1.893 ;
      RECT 7.675 1.525 7.69 1.88 ;
      RECT 7.67 1.525 7.675 1.87 ;
      RECT 7.655 1.525 7.67 1.848 ;
      RECT 7.64 1.525 7.655 1.815 ;
      RECT 7.635 1.525 7.64 1.793 ;
      RECT 7.625 1.525 7.635 1.775 ;
      RECT 7.61 1.525 7.625 1.753 ;
      RECT 7.59 1.525 7.61 1.715 ;
      RECT 7.94 0.81 7.975 1.249 ;
      RECT 7.94 0.81 7.98 1.248 ;
      RECT 7.885 0.87 7.98 1.247 ;
      RECT 7.75 1.042 7.98 1.246 ;
      RECT 7.86 0.92 7.98 1.246 ;
      RECT 7.75 1.042 8.005 1.236 ;
      RECT 7.805 0.987 8.085 1.153 ;
      RECT 7.98 0.781 7.985 1.244 ;
      RECT 7.835 0.957 8.125 1.03 ;
      RECT 7.85 0.94 7.98 1.246 ;
      RECT 7.985 0.78 8.155 0.968 ;
      RECT 7.975 0.783 8.155 0.968 ;
      RECT 7.48 0.66 7.65 0.97 ;
      RECT 7.48 0.66 7.655 0.943 ;
      RECT 7.48 0.66 7.66 0.92 ;
      RECT 7.48 0.66 7.67 0.87 ;
      RECT 7.475 0.765 7.67 0.84 ;
      RECT 7.51 0.335 7.68 0.813 ;
      RECT 7.51 0.335 7.695 0.734 ;
      RECT 7.5 0.545 7.695 0.734 ;
      RECT 7.51 0.345 7.705 0.649 ;
      RECT 7.44 1.087 7.445 1.29 ;
      RECT 7.43 1.075 7.44 1.4 ;
      RECT 7.405 1.075 7.43 1.44 ;
      RECT 7.325 1.075 7.405 1.525 ;
      RECT 7.315 1.075 7.325 1.595 ;
      RECT 7.29 1.075 7.315 1.618 ;
      RECT 7.27 1.075 7.29 1.653 ;
      RECT 7.225 1.085 7.27 1.696 ;
      RECT 7.215 1.097 7.225 1.733 ;
      RECT 7.195 1.111 7.215 1.753 ;
      RECT 7.185 1.129 7.195 1.769 ;
      RECT 7.17 1.155 7.185 1.779 ;
      RECT 7.155 1.196 7.17 1.793 ;
      RECT 7.145 1.231 7.155 1.803 ;
      RECT 7.14 1.247 7.145 1.808 ;
      RECT 7.13 1.262 7.14 1.813 ;
      RECT 7.11 1.305 7.13 1.823 ;
      RECT 7.09 1.342 7.11 1.836 ;
      RECT 7.055 1.365 7.09 1.854 ;
      RECT 7.045 1.379 7.055 1.87 ;
      RECT 7.025 1.389 7.045 1.88 ;
      RECT 7.02 1.398 7.025 1.888 ;
      RECT 7.01 1.405 7.02 1.895 ;
      RECT 7 1.412 7.01 1.903 ;
      RECT 6.985 1.422 7 1.911 ;
      RECT 6.975 1.436 6.985 1.921 ;
      RECT 6.965 1.448 6.975 1.933 ;
      RECT 6.95 1.47 6.965 1.946 ;
      RECT 6.94 1.492 6.95 1.957 ;
      RECT 6.93 1.512 6.94 1.966 ;
      RECT 6.925 1.527 6.93 1.973 ;
      RECT 6.895 1.56 6.925 1.987 ;
      RECT 6.885 1.595 6.895 2.002 ;
      RECT 6.88 1.602 6.885 2.008 ;
      RECT 6.86 1.617 6.88 2.015 ;
      RECT 6.855 1.632 6.86 2.023 ;
      RECT 6.85 1.641 6.855 2.028 ;
      RECT 6.835 1.647 6.85 2.035 ;
      RECT 6.83 1.653 6.835 2.043 ;
      RECT 6.825 1.657 6.83 2.05 ;
      RECT 6.82 1.661 6.825 2.06 ;
      RECT 6.81 1.666 6.82 2.07 ;
      RECT 6.79 1.677 6.81 2.098 ;
      RECT 6.775 1.689 6.79 2.125 ;
      RECT 6.755 1.702 6.775 2.15 ;
      RECT 6.735 1.717 6.755 2.174 ;
      RECT 6.72 1.732 6.735 2.189 ;
      RECT 6.715 1.743 6.72 2.198 ;
      RECT 6.65 1.788 6.715 2.208 ;
      RECT 6.615 1.847 6.65 2.221 ;
      RECT 6.61 1.87 6.615 2.227 ;
      RECT 6.605 1.877 6.61 2.229 ;
      RECT 6.59 1.887 6.605 2.232 ;
      RECT 6.56 1.912 6.59 2.236 ;
      RECT 6.555 1.93 6.56 2.24 ;
      RECT 6.55 1.937 6.555 2.241 ;
      RECT 6.53 1.945 6.55 2.245 ;
      RECT 6.52 1.952 6.53 2.249 ;
      RECT 6.476 1.963 6.52 2.256 ;
      RECT 6.39 1.991 6.476 2.272 ;
      RECT 6.33 2.015 6.39 2.29 ;
      RECT 6.285 2.025 6.33 2.304 ;
      RECT 6.226 2.033 6.285 2.318 ;
      RECT 6.14 2.04 6.226 2.337 ;
      RECT 6.115 2.045 6.14 2.352 ;
      RECT 6.035 2.048 6.115 2.355 ;
      RECT 5.955 2.052 6.035 2.342 ;
      RECT 5.946 2.055 5.955 2.327 ;
      RECT 5.86 2.055 5.946 2.312 ;
      RECT 5.8 2.057 5.86 2.289 ;
      RECT 5.796 2.06 5.8 2.279 ;
      RECT 5.71 2.06 5.796 2.264 ;
      RECT 5.635 2.06 5.71 2.24 ;
      RECT 6.95 1.069 6.96 1.245 ;
      RECT 6.905 1.036 6.95 1.245 ;
      RECT 6.86 0.987 6.905 1.245 ;
      RECT 6.83 0.957 6.86 1.246 ;
      RECT 6.825 0.94 6.83 1.247 ;
      RECT 6.8 0.92 6.825 1.248 ;
      RECT 6.785 0.895 6.8 1.249 ;
      RECT 6.78 0.882 6.785 1.25 ;
      RECT 6.775 0.876 6.78 1.248 ;
      RECT 6.77 0.868 6.775 1.242 ;
      RECT 6.745 0.86 6.77 1.222 ;
      RECT 6.725 0.849 6.745 1.193 ;
      RECT 6.695 0.834 6.725 1.164 ;
      RECT 6.675 0.82 6.695 1.136 ;
      RECT 6.665 0.814 6.675 1.115 ;
      RECT 6.66 0.811 6.665 1.098 ;
      RECT 6.655 0.808 6.66 1.083 ;
      RECT 6.64 0.803 6.655 1.048 ;
      RECT 6.635 0.799 6.64 1.015 ;
      RECT 6.615 0.794 6.635 0.991 ;
      RECT 6.585 0.786 6.615 0.956 ;
      RECT 6.57 0.78 6.585 0.933 ;
      RECT 6.53 0.773 6.57 0.918 ;
      RECT 6.505 0.765 6.53 0.898 ;
      RECT 6.485 0.76 6.505 0.888 ;
      RECT 6.45 0.754 6.485 0.883 ;
      RECT 6.405 0.745 6.45 0.882 ;
      RECT 6.375 0.741 6.405 0.884 ;
      RECT 6.29 0.749 6.375 0.888 ;
      RECT 6.22 0.76 6.29 0.91 ;
      RECT 6.207 0.766 6.22 0.933 ;
      RECT 6.121 0.773 6.207 0.955 ;
      RECT 6.035 0.785 6.121 0.992 ;
      RECT 6.035 1.162 6.045 1.4 ;
      RECT 6.03 0.791 6.035 1.015 ;
      RECT 6.025 1.047 6.035 1.4 ;
      RECT 6.025 0.792 6.03 1.02 ;
      RECT 6.02 0.793 6.025 1.4 ;
      RECT 5.996 0.795 6.02 1.401 ;
      RECT 5.91 0.803 5.996 1.403 ;
      RECT 5.89 0.817 5.91 1.406 ;
      RECT 5.885 0.845 5.89 1.407 ;
      RECT 5.88 0.857 5.885 1.408 ;
      RECT 5.875 0.872 5.88 1.409 ;
      RECT 5.865 0.902 5.875 1.41 ;
      RECT 5.86 0.94 5.865 1.408 ;
      RECT 5.855 0.96 5.86 1.403 ;
      RECT 5.84 0.995 5.855 1.388 ;
      RECT 5.83 1.047 5.84 1.368 ;
      RECT 5.825 1.077 5.83 1.356 ;
      RECT 5.81 1.09 5.825 1.339 ;
      RECT 5.785 1.094 5.81 1.306 ;
      RECT 5.77 1.092 5.785 1.283 ;
      RECT 5.755 1.091 5.77 1.28 ;
      RECT 5.695 1.089 5.755 1.278 ;
      RECT 5.685 1.087 5.695 1.273 ;
      RECT 5.645 1.086 5.685 1.27 ;
      RECT 5.575 1.083 5.645 1.268 ;
      RECT 5.52 1.081 5.575 1.263 ;
      RECT 5.45 1.075 5.52 1.258 ;
      RECT 5.441 1.075 5.45 1.255 ;
      RECT 5.355 1.075 5.441 1.25 ;
      RECT 5.35 1.075 5.355 1.245 ;
      RECT 6.655 0.31 6.83 0.66 ;
      RECT 6.655 0.325 6.84 0.658 ;
      RECT 6.63 0.275 6.775 0.655 ;
      RECT 6.61 0.276 6.775 0.648 ;
      RECT 6.6 0.277 6.785 0.643 ;
      RECT 6.57 0.278 6.785 0.63 ;
      RECT 6.52 0.279 6.785 0.606 ;
      RECT 6.515 0.281 6.785 0.591 ;
      RECT 6.515 0.347 6.845 0.585 ;
      RECT 6.495 0.288 6.8 0.565 ;
      RECT 6.485 0.297 6.81 0.42 ;
      RECT 6.495 0.292 6.81 0.565 ;
      RECT 6.515 0.282 6.8 0.591 ;
      RECT 6.1 1.607 6.27 1.895 ;
      RECT 6.095 1.625 6.28 1.89 ;
      RECT 6.06 1.633 6.345 1.81 ;
      RECT 6.06 1.633 6.431 1.8 ;
      RECT 6.06 1.633 6.485 1.746 ;
      RECT 6.345 1.53 6.515 1.714 ;
      RECT 6.06 1.685 6.52 1.702 ;
      RECT 6.045 1.655 6.515 1.698 ;
      RECT 6.305 1.537 6.345 1.849 ;
      RECT 6.185 1.574 6.515 1.714 ;
      RECT 6.28 1.549 6.305 1.875 ;
      RECT 6.27 1.556 6.515 1.714 ;
      RECT 6.401 1.02 6.47 1.279 ;
      RECT 6.401 1.075 6.475 1.278 ;
      RECT 6.315 1.075 6.475 1.277 ;
      RECT 6.31 1.075 6.48 1.27 ;
      RECT 6.3 1.02 6.47 1.265 ;
      RECT 5.68 0.319 5.855 0.62 ;
      RECT 5.665 0.307 5.68 0.605 ;
      RECT 5.635 0.306 5.665 0.558 ;
      RECT 5.635 0.324 5.86 0.553 ;
      RECT 5.62 0.308 5.68 0.518 ;
      RECT 5.615 0.33 5.87 0.418 ;
      RECT 5.615 0.313 5.766 0.418 ;
      RECT 5.615 0.315 5.77 0.418 ;
      RECT 5.62 0.311 5.766 0.518 ;
      RECT 5.725 1.547 5.73 1.895 ;
      RECT 5.715 1.537 5.725 1.901 ;
      RECT 5.68 1.527 5.715 1.903 ;
      RECT 5.642 1.522 5.68 1.907 ;
      RECT 5.556 1.515 5.642 1.914 ;
      RECT 5.47 1.505 5.556 1.924 ;
      RECT 5.425 1.5 5.47 1.932 ;
      RECT 5.421 1.5 5.425 1.936 ;
      RECT 5.335 1.5 5.421 1.943 ;
      RECT 5.32 1.5 5.335 1.943 ;
      RECT 5.31 1.498 5.32 1.915 ;
      RECT 5.3 1.494 5.31 1.858 ;
      RECT 5.28 1.488 5.3 1.79 ;
      RECT 5.275 1.484 5.28 1.738 ;
      RECT 5.265 1.483 5.275 1.705 ;
      RECT 5.215 1.481 5.265 1.69 ;
      RECT 5.19 1.479 5.215 1.685 ;
      RECT 5.147 1.477 5.19 1.681 ;
      RECT 5.061 1.473 5.147 1.669 ;
      RECT 4.975 1.468 5.061 1.653 ;
      RECT 4.945 1.465 4.975 1.64 ;
      RECT 4.92 1.464 4.945 1.628 ;
      RECT 4.915 1.464 4.92 1.618 ;
      RECT 4.875 1.463 4.915 1.61 ;
      RECT 4.86 1.462 4.875 1.603 ;
      RECT 4.81 1.461 4.86 1.595 ;
      RECT 4.808 1.46 4.81 1.59 ;
      RECT 4.722 1.458 4.808 1.59 ;
      RECT 4.636 1.453 4.722 1.59 ;
      RECT 4.55 1.449 4.636 1.59 ;
      RECT 4.501 1.445 4.55 1.588 ;
      RECT 4.415 1.442 4.501 1.583 ;
      RECT 4.392 1.439 4.415 1.579 ;
      RECT 4.306 1.436 4.392 1.574 ;
      RECT 4.22 1.432 4.306 1.565 ;
      RECT 4.195 1.425 4.22 1.56 ;
      RECT 4.135 1.39 4.195 1.557 ;
      RECT 4.115 1.315 4.135 1.554 ;
      RECT 4.11 1.257 4.115 1.553 ;
      RECT 4.085 1.197 4.11 1.552 ;
      RECT 4.01 1.075 4.085 1.548 ;
      RECT 4 1.075 4.01 1.54 ;
      RECT 3.985 1.075 4 1.53 ;
      RECT 3.97 1.075 3.985 1.5 ;
      RECT 3.955 1.075 3.97 1.445 ;
      RECT 3.94 1.075 3.955 1.383 ;
      RECT 3.915 1.075 3.94 1.308 ;
      RECT 3.91 1.075 3.915 1.258 ;
      RECT 5.255 0.62 5.275 0.929 ;
      RECT 5.241 0.622 5.29 0.926 ;
      RECT 5.241 0.627 5.31 0.917 ;
      RECT 5.155 0.625 5.29 0.911 ;
      RECT 5.155 0.633 5.345 0.894 ;
      RECT 5.12 0.635 5.345 0.893 ;
      RECT 5.09 0.643 5.345 0.884 ;
      RECT 5.08 0.648 5.365 0.87 ;
      RECT 5.12 0.638 5.365 0.87 ;
      RECT 5.12 0.641 5.375 0.858 ;
      RECT 5.09 0.643 5.385 0.845 ;
      RECT 5.09 0.647 5.395 0.788 ;
      RECT 5.08 0.652 5.4 0.703 ;
      RECT 5.241 0.62 5.275 0.926 ;
      RECT 4.68 0.723 4.685 0.935 ;
      RECT 4.555 0.72 4.57 0.935 ;
      RECT 4.02 0.75 4.09 0.935 ;
      RECT 3.905 0.75 3.94 0.93 ;
      RECT 5.026 1.052 5.045 1.246 ;
      RECT 4.94 1.007 5.026 1.247 ;
      RECT 4.93 0.96 4.94 1.249 ;
      RECT 4.925 0.94 4.93 1.25 ;
      RECT 4.905 0.905 4.925 1.251 ;
      RECT 4.89 0.855 4.905 1.252 ;
      RECT 4.87 0.792 4.89 1.253 ;
      RECT 4.86 0.755 4.87 1.254 ;
      RECT 4.845 0.744 4.86 1.255 ;
      RECT 4.84 0.736 4.845 1.253 ;
      RECT 4.83 0.735 4.84 1.245 ;
      RECT 4.8 0.732 4.83 1.224 ;
      RECT 4.725 0.727 4.8 1.169 ;
      RECT 4.71 0.723 4.725 1.115 ;
      RECT 4.7 0.723 4.71 1.01 ;
      RECT 4.685 0.723 4.7 0.943 ;
      RECT 4.67 0.723 4.68 0.933 ;
      RECT 4.615 0.722 4.67 0.93 ;
      RECT 4.57 0.72 4.615 0.933 ;
      RECT 4.542 0.72 4.555 0.936 ;
      RECT 4.456 0.724 4.542 0.938 ;
      RECT 4.37 0.73 4.456 0.943 ;
      RECT 4.35 0.734 4.37 0.945 ;
      RECT 4.348 0.735 4.35 0.944 ;
      RECT 4.262 0.737 4.348 0.943 ;
      RECT 4.176 0.742 4.262 0.94 ;
      RECT 4.09 0.747 4.176 0.937 ;
      RECT 3.94 0.75 4.02 0.933 ;
      RECT 4.716 1.725 4.765 2.059 ;
      RECT 4.716 1.725 4.77 2.058 ;
      RECT 4.63 1.725 4.77 2.057 ;
      RECT 4.405 1.833 4.775 2.055 ;
      RECT 4.63 1.725 4.8 2.048 ;
      RECT 4.6 1.737 4.805 2.039 ;
      RECT 4.585 1.755 4.81 2.036 ;
      RECT 4.4 1.839 4.81 1.963 ;
      RECT 4.395 1.846 4.81 1.923 ;
      RECT 4.41 1.812 4.81 2.036 ;
      RECT 4.571 1.758 4.775 2.055 ;
      RECT 4.485 1.778 4.81 2.036 ;
      RECT 4.585 1.752 4.805 2.039 ;
      RECT 4.355 1.076 4.545 1.27 ;
      RECT 4.35 1.078 4.545 1.269 ;
      RECT 4.345 1.082 4.56 1.266 ;
      RECT 4.36 1.075 4.56 1.266 ;
      RECT 4.345 1.185 4.565 1.261 ;
      RECT 3.64 1.685 3.731 1.983 ;
      RECT 3.635 1.687 3.81 1.978 ;
      RECT 3.64 1.685 3.81 1.978 ;
      RECT 3.635 1.691 3.83 1.976 ;
      RECT 3.635 1.746 3.87 1.975 ;
      RECT 3.635 1.781 3.885 1.969 ;
      RECT 3.635 1.815 3.895 1.959 ;
      RECT 3.625 1.695 3.83 1.81 ;
      RECT 3.625 1.715 3.845 1.81 ;
      RECT 3.625 1.698 3.835 1.81 ;
      RECT 3.85 0.466 3.855 0.528 ;
      RECT 3.845 0.388 3.85 0.551 ;
      RECT 3.84 0.345 3.845 0.562 ;
      RECT 3.835 0.335 3.84 0.574 ;
      RECT 3.83 0.335 3.835 0.583 ;
      RECT 3.805 0.335 3.83 0.615 ;
      RECT 3.8 0.335 3.805 0.648 ;
      RECT 3.785 0.335 3.8 0.673 ;
      RECT 3.775 0.335 3.785 0.7 ;
      RECT 3.77 0.335 3.775 0.713 ;
      RECT 3.765 0.335 3.77 0.728 ;
      RECT 3.755 0.335 3.765 0.743 ;
      RECT 3.75 0.335 3.755 0.763 ;
      RECT 3.725 0.335 3.75 0.798 ;
      RECT 3.68 0.335 3.725 0.843 ;
      RECT 3.67 0.335 3.68 0.856 ;
      RECT 3.585 0.42 3.67 0.863 ;
      RECT 3.55 0.542 3.585 0.872 ;
      RECT 3.545 0.582 3.55 0.876 ;
      RECT 3.525 0.605 3.545 0.878 ;
      RECT 3.52 0.635 3.525 0.881 ;
      RECT 3.51 0.647 3.52 0.882 ;
      RECT 3.465 0.67 3.51 0.887 ;
      RECT 3.425 0.7 3.465 0.895 ;
      RECT 3.39 0.712 3.425 0.901 ;
      RECT 3.385 0.717 3.39 0.905 ;
      RECT 3.315 0.727 3.385 0.912 ;
      RECT 3.275 0.737 3.315 0.922 ;
      RECT 3.255 0.742 3.275 0.928 ;
      RECT 3.245 0.746 3.255 0.933 ;
      RECT 3.24 0.749 3.245 0.936 ;
      RECT 3.23 0.75 3.24 0.937 ;
      RECT 3.205 0.752 3.23 0.941 ;
      RECT 3.195 0.757 3.205 0.944 ;
      RECT 3.15 0.765 3.195 0.945 ;
      RECT 3.025 0.77 3.15 0.945 ;
      RECT 3.58 1.067 3.6 1.249 ;
      RECT 3.531 1.052 3.58 1.248 ;
      RECT 3.445 1.067 3.6 1.246 ;
      RECT 3.43 1.067 3.6 1.245 ;
      RECT 3.395 1.045 3.565 1.23 ;
      RECT 3.465 2.065 3.48 2.274 ;
      RECT 3.465 2.073 3.485 2.273 ;
      RECT 3.41 2.073 3.485 2.272 ;
      RECT 3.39 2.077 3.49 2.27 ;
      RECT 3.37 2.027 3.41 2.269 ;
      RECT 3.315 2.085 3.495 2.267 ;
      RECT 3.28 2.042 3.41 2.265 ;
      RECT 3.276 2.045 3.465 2.264 ;
      RECT 3.19 2.053 3.465 2.262 ;
      RECT 3.19 2.097 3.5 2.255 ;
      RECT 3.18 2.19 3.5 2.253 ;
      RECT 3.19 2.109 3.505 2.238 ;
      RECT 3.19 2.13 3.52 2.208 ;
      RECT 3.19 2.157 3.525 2.178 ;
      RECT 3.315 2.035 3.41 2.267 ;
      RECT 2.945 1.08 2.95 1.618 ;
      RECT 2.75 1.41 2.755 1.605 ;
      RECT 1.05 1.075 1.065 1.455 ;
      RECT 3.115 1.075 3.12 1.245 ;
      RECT 3.11 1.075 3.115 1.255 ;
      RECT 3.105 1.075 3.11 1.268 ;
      RECT 3.08 1.075 3.105 1.31 ;
      RECT 3.055 1.075 3.08 1.383 ;
      RECT 3.04 1.075 3.055 1.435 ;
      RECT 3.035 1.075 3.04 1.465 ;
      RECT 3.01 1.075 3.035 1.505 ;
      RECT 2.995 1.075 3.01 1.56 ;
      RECT 2.99 1.075 2.995 1.593 ;
      RECT 2.965 1.075 2.99 1.613 ;
      RECT 2.95 1.075 2.965 1.619 ;
      RECT 2.88 1.11 2.945 1.615 ;
      RECT 2.83 1.165 2.88 1.61 ;
      RECT 2.82 1.197 2.83 1.608 ;
      RECT 2.815 1.222 2.82 1.608 ;
      RECT 2.795 1.295 2.815 1.608 ;
      RECT 2.785 1.375 2.795 1.607 ;
      RECT 2.77 1.405 2.785 1.607 ;
      RECT 2.755 1.41 2.77 1.606 ;
      RECT 2.695 1.412 2.75 1.603 ;
      RECT 2.665 1.417 2.695 1.599 ;
      RECT 2.663 1.42 2.665 1.598 ;
      RECT 2.577 1.422 2.663 1.595 ;
      RECT 2.491 1.428 2.577 1.589 ;
      RECT 2.405 1.433 2.491 1.583 ;
      RECT 2.332 1.438 2.405 1.584 ;
      RECT 2.246 1.444 2.332 1.592 ;
      RECT 2.16 1.45 2.246 1.601 ;
      RECT 2.14 1.454 2.16 1.606 ;
      RECT 2.093 1.456 2.14 1.609 ;
      RECT 2.007 1.461 2.093 1.615 ;
      RECT 1.921 1.466 2.007 1.624 ;
      RECT 1.835 1.472 1.921 1.632 ;
      RECT 1.75 1.47 1.835 1.641 ;
      RECT 1.746 1.465 1.75 1.645 ;
      RECT 1.66 1.46 1.746 1.637 ;
      RECT 1.596 1.451 1.66 1.625 ;
      RECT 1.51 1.442 1.596 1.612 ;
      RECT 1.486 1.435 1.51 1.603 ;
      RECT 1.4 1.429 1.486 1.59 ;
      RECT 1.36 1.422 1.4 1.576 ;
      RECT 1.355 1.412 1.36 1.572 ;
      RECT 1.345 1.4 1.355 1.571 ;
      RECT 1.325 1.37 1.345 1.568 ;
      RECT 1.27 1.29 1.325 1.562 ;
      RECT 1.25 1.209 1.27 1.557 ;
      RECT 1.23 1.167 1.25 1.553 ;
      RECT 1.205 1.12 1.23 1.547 ;
      RECT 1.2 1.095 1.205 1.544 ;
      RECT 1.165 1.075 1.2 1.539 ;
      RECT 1.156 1.075 1.165 1.532 ;
      RECT 1.07 1.075 1.156 1.502 ;
      RECT 1.065 1.075 1.07 1.465 ;
      RECT 1.03 1.075 1.05 1.387 ;
      RECT 1.025 1.117 1.03 1.352 ;
      RECT 1.02 1.192 1.025 1.308 ;
      RECT 2.47 0.997 2.645 1.245 ;
      RECT 2.47 0.997 2.65 1.243 ;
      RECT 2.465 1.029 2.65 1.203 ;
      RECT 2.495 0.97 2.665 1.19 ;
      RECT 2.46 1.047 2.665 1.123 ;
      RECT 1.77 0.51 1.94 0.685 ;
      RECT 1.77 0.51 2.112 0.677 ;
      RECT 1.77 0.51 2.195 0.671 ;
      RECT 1.77 0.51 2.23 0.667 ;
      RECT 1.77 0.51 2.25 0.666 ;
      RECT 1.77 0.51 2.336 0.662 ;
      RECT 2.23 0.335 2.4 0.657 ;
      RECT 1.805 0.442 2.43 0.655 ;
      RECT 1.795 0.497 2.435 0.653 ;
      RECT 1.77 0.533 2.445 0.648 ;
      RECT 1.77 0.56 2.45 0.578 ;
      RECT 1.835 0.385 2.41 0.655 ;
      RECT 2.026 0.37 2.41 0.655 ;
      RECT 1.86 0.373 2.41 0.655 ;
      RECT 1.94 0.371 2.026 0.682 ;
      RECT 2.026 0.368 2.405 0.655 ;
      RECT 2.21 0.345 2.405 0.655 ;
      RECT 2.112 0.366 2.405 0.655 ;
      RECT 2.195 0.36 2.21 0.668 ;
      RECT 2.345 1.725 2.35 1.925 ;
      RECT 1.81 1.79 1.855 1.925 ;
      RECT 2.38 1.725 2.4 1.898 ;
      RECT 2.35 1.725 2.38 1.913 ;
      RECT 2.285 1.725 2.345 1.95 ;
      RECT 2.27 1.725 2.285 1.98 ;
      RECT 2.255 1.725 2.27 1.993 ;
      RECT 2.235 1.725 2.255 2.008 ;
      RECT 2.23 1.725 2.235 2.017 ;
      RECT 2.22 1.729 2.23 2.022 ;
      RECT 2.205 1.739 2.22 2.033 ;
      RECT 2.18 1.755 2.205 2.043 ;
      RECT 2.17 1.769 2.18 2.045 ;
      RECT 2.15 1.781 2.17 2.042 ;
      RECT 2.12 1.802 2.15 2.036 ;
      RECT 2.11 1.814 2.12 2.031 ;
      RECT 2.1 1.812 2.11 2.028 ;
      RECT 2.085 1.811 2.1 2.023 ;
      RECT 2.08 1.81 2.085 2.018 ;
      RECT 2.045 1.808 2.08 2.008 ;
      RECT 2.025 1.805 2.045 1.99 ;
      RECT 2.015 1.803 2.025 1.985 ;
      RECT 2.005 1.802 2.015 1.98 ;
      RECT 1.97 1.8 2.005 1.968 ;
      RECT 1.915 1.796 1.97 1.948 ;
      RECT 1.905 1.794 1.915 1.933 ;
      RECT 1.9 1.794 1.905 1.928 ;
      RECT 1.855 1.792 1.9 1.925 ;
      RECT 1.76 1.79 1.81 1.929 ;
      RECT 1.75 1.791 1.76 1.934 ;
      RECT 1.69 1.798 1.75 1.948 ;
      RECT 1.665 1.806 1.69 1.968 ;
      RECT 1.655 1.81 1.665 1.98 ;
      RECT 1.65 1.811 1.655 1.985 ;
      RECT 1.635 1.813 1.65 1.988 ;
      RECT 1.62 1.815 1.635 1.993 ;
      RECT 1.615 1.815 1.62 1.996 ;
      RECT 1.57 1.82 1.615 2.007 ;
      RECT 1.565 1.824 1.57 2.019 ;
      RECT 1.54 1.82 1.565 2.023 ;
      RECT 1.53 1.816 1.54 2.027 ;
      RECT 1.52 1.815 1.53 2.031 ;
      RECT 1.505 1.805 1.52 2.037 ;
      RECT 1.5 1.793 1.505 2.041 ;
      RECT 1.495 1.79 1.5 2.042 ;
      RECT 1.49 1.787 1.495 2.044 ;
      RECT 1.475 1.775 1.49 2.043 ;
      RECT 1.46 1.757 1.475 2.04 ;
      RECT 1.44 1.736 1.46 2.033 ;
      RECT 1.375 1.725 1.44 2.005 ;
      RECT 1.371 1.725 1.375 1.984 ;
      RECT 1.285 1.725 1.371 1.954 ;
      RECT 1.27 1.725 1.285 1.91 ;
      RECT 1.845 0.825 1.85 1.06 ;
      RECT 0.975 0.741 0.98 0.945 ;
      RECT 1.555 0.77 1.56 0.925 ;
      RECT 1.475 0.75 1.48 0.925 ;
      RECT 2.145 0.892 2.16 1.245 ;
      RECT 2.071 0.877 2.145 1.245 ;
      RECT 1.985 0.86 2.071 1.245 ;
      RECT 1.975 0.85 1.985 1.243 ;
      RECT 1.97 0.848 1.975 1.238 ;
      RECT 1.955 0.846 1.97 1.224 ;
      RECT 1.885 0.838 1.955 1.164 ;
      RECT 1.865 0.829 1.885 1.098 ;
      RECT 1.86 0.826 1.865 1.078 ;
      RECT 1.85 0.825 1.86 1.068 ;
      RECT 1.84 0.825 1.845 1.052 ;
      RECT 1.83 0.824 1.84 1.042 ;
      RECT 1.82 0.822 1.83 1.03 ;
      RECT 1.805 0.819 1.82 1.01 ;
      RECT 1.795 0.817 1.805 0.995 ;
      RECT 1.775 0.814 1.795 0.983 ;
      RECT 1.77 0.812 1.775 0.973 ;
      RECT 1.745 0.81 1.77 0.96 ;
      RECT 1.715 0.805 1.745 0.945 ;
      RECT 1.635 0.796 1.715 0.936 ;
      RECT 1.59 0.785 1.635 0.929 ;
      RECT 1.57 0.776 1.59 0.926 ;
      RECT 1.56 0.771 1.57 0.925 ;
      RECT 1.515 0.765 1.555 0.925 ;
      RECT 1.5 0.757 1.515 0.925 ;
      RECT 1.48 0.752 1.5 0.925 ;
      RECT 1.46 0.749 1.475 0.925 ;
      RECT 1.377 0.748 1.46 0.924 ;
      RECT 1.291 0.747 1.377 0.92 ;
      RECT 1.205 0.745 1.291 0.917 ;
      RECT 1.152 0.744 1.205 0.919 ;
      RECT 1.066 0.743 1.152 0.928 ;
      RECT 0.98 0.742 1.066 0.94 ;
      RECT 0.96 0.741 0.975 0.948 ;
      RECT 0.88 0.74 0.96 0.96 ;
      RECT 0.855 0.74 0.88 0.973 ;
      RECT 0.83 0.74 0.855 0.988 ;
      RECT 0.825 0.74 0.83 1.01 ;
      RECT 0.82 0.74 0.825 1.028 ;
      RECT 0.815 0.74 0.82 1.045 ;
      RECT 0.81 0.74 0.815 1.058 ;
      RECT 0.805 0.74 0.81 1.068 ;
      RECT 0.765 0.74 0.805 1.153 ;
      RECT 0.75 0.74 0.765 1.238 ;
      RECT 0.74 0.741 0.75 1.25 ;
      RECT 0.705 0.746 0.74 1.255 ;
      RECT 0.665 0.755 0.705 1.255 ;
      RECT 0.65 0.765 0.665 1.255 ;
      RECT 0.645 0.775 0.65 1.255 ;
      RECT 0.625 0.802 0.645 1.255 ;
      RECT 0.575 0.885 0.625 1.255 ;
      RECT 0.57 0.947 0.575 1.255 ;
      RECT 0.56 0.96 0.57 1.255 ;
      RECT 0.55 0.982 0.56 1.255 ;
      RECT 0.54 1.007 0.55 1.25 ;
      RECT 0.535 1.045 0.54 1.243 ;
      RECT 0.525 1.155 0.535 1.238 ;
      RECT 1.92 2.076 1.935 2.335 ;
      RECT 1.92 2.091 1.94 2.334 ;
      RECT 1.836 2.091 1.94 2.332 ;
      RECT 1.836 2.105 1.945 2.331 ;
      RECT 1.75 2.147 1.95 2.328 ;
      RECT 1.745 2.09 1.935 2.323 ;
      RECT 1.745 2.161 1.955 2.32 ;
      RECT 1.74 2.192 1.955 2.318 ;
      RECT 1.745 2.189 1.97 2.308 ;
      RECT 1.74 2.235 1.985 2.293 ;
      RECT 1.74 2.263 1.99 2.278 ;
      RECT 1.75 2.065 1.92 2.328 ;
      RECT 1.51 1.075 1.68 1.245 ;
      RECT 1.475 1.075 1.68 1.24 ;
      RECT 1.465 1.075 1.68 1.233 ;
      RECT 1.46 1.06 1.63 1.23 ;
      RECT 0.29 1.597 0.555 2.04 ;
      RECT 0.285 1.568 0.5 2.038 ;
      RECT 0.28 1.722 0.56 2.033 ;
      RECT 0.285 1.617 0.56 2.033 ;
      RECT 0.285 1.628 0.57 2.02 ;
      RECT 0.285 1.575 0.53 2.038 ;
      RECT 0.29 1.562 0.5 2.04 ;
      RECT 0.29 1.56 0.45 2.04 ;
      RECT 0.391 1.552 0.45 2.04 ;
      RECT 0.305 1.553 0.45 2.04 ;
      RECT 0.391 1.551 0.44 2.04 ;
      RECT 0.195 0.366 0.37 0.665 ;
      RECT 0.245 0.328 0.37 0.665 ;
      RECT 0.23 0.33 0.456 0.657 ;
      RECT 0.23 0.333 0.495 0.644 ;
      RECT 0.23 0.334 0.505 0.63 ;
      RECT 0.185 0.385 0.505 0.62 ;
      RECT 0.23 0.335 0.51 0.615 ;
      RECT 0.185 0.545 0.515 0.605 ;
      RECT 0.17 0.405 0.51 0.545 ;
      RECT 0.165 0.421 0.51 0.485 ;
      RECT 0.21 0.345 0.51 0.615 ;
      RECT 0.245 0.326 0.331 0.665 ;
  END
END scs130hd_mpr2ya_8

MACRO sky130_osu_ring_oscillator_mpr2aa_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2aa_8 0 0 ;
  SIZE 79.25 BY 8.88 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT 72.065 1.85 72.395 2.58 ;
      RECT 72.025 1.735 72.205 2.385 ;
      RECT 68.525 3.535 68.855 3.865 ;
      RECT 67.32 3.55 68.855 3.85 ;
      RECT 67.32 2.43 67.62 3.85 ;
      RECT 67.065 2.415 67.395 2.745 ;
      RECT 56.215 1.85 56.545 2.58 ;
      RECT 56.175 1.735 56.355 2.385 ;
      RECT 52.675 3.535 53.005 3.865 ;
      RECT 51.47 3.55 53.005 3.85 ;
      RECT 51.47 2.43 51.77 3.85 ;
      RECT 51.215 2.415 51.545 2.745 ;
      RECT 40.365 1.85 40.695 2.58 ;
      RECT 40.325 1.735 40.505 2.385 ;
      RECT 36.825 3.535 37.155 3.865 ;
      RECT 35.62 3.55 37.155 3.85 ;
      RECT 35.62 2.43 35.92 3.85 ;
      RECT 35.365 2.415 35.695 2.745 ;
      RECT 24.515 1.85 24.845 2.58 ;
      RECT 24.475 1.735 24.655 2.385 ;
      RECT 20.975 3.535 21.305 3.865 ;
      RECT 19.77 3.55 21.305 3.85 ;
      RECT 19.77 2.43 20.07 3.85 ;
      RECT 19.515 2.415 19.845 2.745 ;
      RECT 8.665 1.85 8.995 2.58 ;
      RECT 8.625 1.735 8.805 2.385 ;
      RECT 5.125 3.535 5.455 3.865 ;
      RECT 3.92 3.55 5.455 3.85 ;
      RECT 3.92 2.43 4.22 3.85 ;
      RECT 3.665 2.415 3.995 2.745 ;
      RECT 72.545 2.975 72.875 3.705 ;
      RECT 70.465 2.575 70.795 3.305 ;
      RECT 68.905 2.015 69.235 2.745 ;
      RECT 68.025 2.015 68.355 2.745 ;
      RECT 66.345 2.415 66.675 3.145 ;
      RECT 65.345 1.855 65.675 2.585 ;
      RECT 63.905 2.575 64.235 3.305 ;
      RECT 56.695 2.975 57.025 3.705 ;
      RECT 54.615 2.575 54.945 3.305 ;
      RECT 53.055 2.015 53.385 2.745 ;
      RECT 52.175 2.015 52.505 2.745 ;
      RECT 50.495 2.415 50.825 3.145 ;
      RECT 49.495 1.855 49.825 2.585 ;
      RECT 48.055 2.575 48.385 3.305 ;
      RECT 40.845 2.975 41.175 3.705 ;
      RECT 38.765 2.575 39.095 3.305 ;
      RECT 37.205 2.015 37.535 2.745 ;
      RECT 36.325 2.015 36.655 2.745 ;
      RECT 34.645 2.415 34.975 3.145 ;
      RECT 33.645 1.855 33.975 2.585 ;
      RECT 32.205 2.575 32.535 3.305 ;
      RECT 24.995 2.975 25.325 3.705 ;
      RECT 22.915 2.575 23.245 3.305 ;
      RECT 21.355 2.015 21.685 2.745 ;
      RECT 20.475 2.015 20.805 2.745 ;
      RECT 18.795 2.415 19.125 3.145 ;
      RECT 17.795 1.855 18.125 2.585 ;
      RECT 16.355 2.575 16.685 3.305 ;
      RECT 9.145 2.975 9.475 3.705 ;
      RECT 7.065 2.575 7.395 3.305 ;
      RECT 5.505 2.015 5.835 2.745 ;
      RECT 4.625 2.015 4.955 2.745 ;
      RECT 2.945 2.415 3.275 3.145 ;
      RECT 1.945 1.855 2.275 2.585 ;
      RECT 0.505 2.575 0.835 3.305 ;
    LAYER via2 ;
      RECT 72.61 3.04 72.81 3.24 ;
      RECT 72.13 2.315 72.33 2.515 ;
      RECT 70.53 3.04 70.73 3.24 ;
      RECT 68.97 2.48 69.17 2.68 ;
      RECT 68.59 3.6 68.79 3.8 ;
      RECT 68.09 2.48 68.29 2.68 ;
      RECT 67.13 2.48 67.33 2.68 ;
      RECT 66.41 2.48 66.61 2.68 ;
      RECT 65.41 1.92 65.61 2.12 ;
      RECT 63.97 3.04 64.17 3.24 ;
      RECT 56.76 3.04 56.96 3.24 ;
      RECT 56.28 2.315 56.48 2.515 ;
      RECT 54.68 3.04 54.88 3.24 ;
      RECT 53.12 2.48 53.32 2.68 ;
      RECT 52.74 3.6 52.94 3.8 ;
      RECT 52.24 2.48 52.44 2.68 ;
      RECT 51.28 2.48 51.48 2.68 ;
      RECT 50.56 2.48 50.76 2.68 ;
      RECT 49.56 1.92 49.76 2.12 ;
      RECT 48.12 3.04 48.32 3.24 ;
      RECT 40.91 3.04 41.11 3.24 ;
      RECT 40.43 2.315 40.63 2.515 ;
      RECT 38.83 3.04 39.03 3.24 ;
      RECT 37.27 2.48 37.47 2.68 ;
      RECT 36.89 3.6 37.09 3.8 ;
      RECT 36.39 2.48 36.59 2.68 ;
      RECT 35.43 2.48 35.63 2.68 ;
      RECT 34.71 2.48 34.91 2.68 ;
      RECT 33.71 1.92 33.91 2.12 ;
      RECT 32.27 3.04 32.47 3.24 ;
      RECT 25.06 3.04 25.26 3.24 ;
      RECT 24.58 2.315 24.78 2.515 ;
      RECT 22.98 3.04 23.18 3.24 ;
      RECT 21.42 2.48 21.62 2.68 ;
      RECT 21.04 3.6 21.24 3.8 ;
      RECT 20.54 2.48 20.74 2.68 ;
      RECT 19.58 2.48 19.78 2.68 ;
      RECT 18.86 2.48 19.06 2.68 ;
      RECT 17.86 1.92 18.06 2.12 ;
      RECT 16.42 3.04 16.62 3.24 ;
      RECT 9.21 3.04 9.41 3.24 ;
      RECT 8.73 2.315 8.93 2.515 ;
      RECT 7.13 3.04 7.33 3.24 ;
      RECT 5.57 2.48 5.77 2.68 ;
      RECT 5.19 3.6 5.39 3.8 ;
      RECT 4.69 2.48 4.89 2.68 ;
      RECT 3.73 2.48 3.93 2.68 ;
      RECT 3.01 2.48 3.21 2.68 ;
      RECT 2.01 1.92 2.21 2.12 ;
      RECT 0.57 3.04 0.77 3.24 ;
    LAYER met2 ;
      RECT 12.12 6.28 12.44 6.605 ;
      RECT 12.15 5.695 12.32 6.605 ;
      RECT 12.15 5.695 12.325 6.045 ;
      RECT 12.15 5.695 13.125 5.87 ;
      RECT 12.95 1.965 13.125 5.87 ;
      RECT 9.17 2.84 9.45 3.28 ;
      RECT 9.17 2.84 9.455 3.238 ;
      RECT 9.17 2.84 9.46 3.135 ;
      RECT 9.17 2.84 9.462 3.015 ;
      RECT 9.17 2.84 10.095 3.01 ;
      RECT 9.925 2.025 10.095 3.01 ;
      RECT 9.17 2.805 9.43 3.28 ;
      RECT 78.71 0.305 78.885 2.525 ;
      RECT 78.655 2.165 79.005 2.515 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 9.925 2.025 13.245 2.195 ;
      RECT 78.705 0.305 78.89 2.515 ;
      RECT 10.95 0.305 11.11 2.195 ;
      RECT 10.95 0.305 78.89 0.465 ;
      RECT 75.52 6.28 75.84 6.605 ;
      RECT 75.55 5.695 75.72 6.605 ;
      RECT 75.55 5.695 75.725 6.045 ;
      RECT 75.55 5.695 76.525 5.87 ;
      RECT 76.35 1.965 76.525 5.87 ;
      RECT 72.57 2.84 72.85 3.28 ;
      RECT 72.57 2.84 72.855 3.238 ;
      RECT 72.57 2.84 72.86 3.135 ;
      RECT 72.57 2.84 72.862 3.015 ;
      RECT 72.57 2.84 73.495 3.01 ;
      RECT 73.325 2.025 73.495 3.01 ;
      RECT 72.57 2.805 72.83 3.28 ;
      RECT 76.295 1.965 76.645 2.315 ;
      RECT 73.325 2.025 76.645 2.195 ;
      RECT 74.555 0.915 74.725 2.195 ;
      RECT 62.83 0.885 63.18 1.235 ;
      RECT 62.83 0.915 74.725 1.085 ;
      RECT 76.32 6.655 76.645 6.98 ;
      RECT 75.205 6.745 76.645 6.915 ;
      RECT 75.205 2.395 75.365 6.915 ;
      RECT 75.52 2.365 75.84 2.685 ;
      RECT 75.205 2.395 75.84 2.565 ;
      RECT 74.47 5.855 74.82 6.205 ;
      RECT 74.54 2.705 74.715 6.205 ;
      RECT 74.465 2.705 74.815 3.055 ;
      RECT 63.93 3 64.21 3.28 ;
      RECT 63.9 3 64.21 3.265 ;
      RECT 63.895 2.963 64.155 3.263 ;
      RECT 63.89 2.964 64.155 3.257 ;
      RECT 63.885 2.967 64.155 3.25 ;
      RECT 63.88 3 64.21 3.243 ;
      RECT 63.85 2.97 64.155 3.23 ;
      RECT 63.85 2.997 64.175 3.23 ;
      RECT 63.85 2.987 64.17 3.23 ;
      RECT 63.85 2.972 64.165 3.23 ;
      RECT 63.95 2.962 64.155 3.28 ;
      RECT 63.95 2.957 64.145 3.28 ;
      RECT 63.95 2.955 64.13 3.28 ;
      RECT 63.95 1.42 64.125 3.28 ;
      RECT 73.86 1.34 74.21 1.69 ;
      RECT 63.95 1.42 74.21 1.595 ;
      RECT 69.64 2.455 69.875 2.715 ;
      RECT 72.785 2.235 72.95 2.495 ;
      RECT 72.69 2.225 72.705 2.495 ;
      RECT 71.29 1.795 71.33 1.935 ;
      RECT 72.705 2.23 72.785 2.495 ;
      RECT 72.65 2.225 72.69 2.461 ;
      RECT 72.636 2.225 72.65 2.461 ;
      RECT 72.55 2.23 72.636 2.463 ;
      RECT 72.505 2.237 72.55 2.465 ;
      RECT 72.475 2.237 72.505 2.467 ;
      RECT 72.45 2.232 72.475 2.469 ;
      RECT 72.42 2.228 72.45 2.478 ;
      RECT 72.41 2.225 72.42 2.49 ;
      RECT 72.405 2.225 72.41 2.498 ;
      RECT 72.4 2.225 72.405 2.503 ;
      RECT 72.39 2.224 72.4 2.513 ;
      RECT 72.385 2.223 72.39 2.523 ;
      RECT 72.37 2.222 72.385 2.528 ;
      RECT 72.342 2.219 72.37 2.555 ;
      RECT 72.256 2.211 72.342 2.555 ;
      RECT 72.17 2.2 72.256 2.555 ;
      RECT 72.13 2.185 72.17 2.555 ;
      RECT 72.09 2.159 72.13 2.555 ;
      RECT 72.085 2.141 72.09 2.367 ;
      RECT 72.075 2.137 72.085 2.357 ;
      RECT 72.06 2.127 72.075 2.344 ;
      RECT 72.04 2.111 72.06 2.329 ;
      RECT 72.025 2.096 72.04 2.314 ;
      RECT 72.015 2.085 72.025 2.304 ;
      RECT 71.99 2.069 72.015 2.293 ;
      RECT 71.985 2.056 71.99 2.283 ;
      RECT 71.98 2.052 71.985 2.278 ;
      RECT 71.925 2.038 71.98 2.256 ;
      RECT 71.886 2.019 71.925 2.22 ;
      RECT 71.8 1.993 71.886 2.173 ;
      RECT 71.796 1.975 71.8 2.139 ;
      RECT 71.71 1.956 71.796 2.117 ;
      RECT 71.705 1.938 71.71 2.095 ;
      RECT 71.7 1.936 71.705 2.093 ;
      RECT 71.69 1.935 71.7 2.088 ;
      RECT 71.63 1.922 71.69 2.074 ;
      RECT 71.585 1.9 71.63 2.053 ;
      RECT 71.525 1.877 71.585 2.032 ;
      RECT 71.461 1.852 71.525 2.007 ;
      RECT 71.375 1.822 71.461 1.976 ;
      RECT 71.36 1.802 71.375 1.955 ;
      RECT 71.33 1.797 71.36 1.946 ;
      RECT 71.277 1.795 71.29 1.935 ;
      RECT 71.191 1.795 71.277 1.937 ;
      RECT 71.105 1.795 71.191 1.939 ;
      RECT 71.085 1.795 71.105 1.943 ;
      RECT 71.04 1.797 71.085 1.954 ;
      RECT 71 1.807 71.04 1.97 ;
      RECT 70.996 1.816 71 1.978 ;
      RECT 70.91 1.836 70.996 1.994 ;
      RECT 70.9 1.855 70.91 2.012 ;
      RECT 70.895 1.857 70.9 2.015 ;
      RECT 70.885 1.861 70.895 2.018 ;
      RECT 70.865 1.866 70.885 2.028 ;
      RECT 70.835 1.876 70.865 2.048 ;
      RECT 70.83 1.883 70.835 2.062 ;
      RECT 70.82 1.887 70.83 2.069 ;
      RECT 70.805 1.895 70.82 2.08 ;
      RECT 70.795 1.905 70.805 2.091 ;
      RECT 70.785 1.912 70.795 2.099 ;
      RECT 70.76 1.925 70.785 2.114 ;
      RECT 70.696 1.961 70.76 2.153 ;
      RECT 70.61 2.024 70.696 2.217 ;
      RECT 70.575 2.075 70.61 2.27 ;
      RECT 70.57 2.092 70.575 2.287 ;
      RECT 70.555 2.101 70.57 2.294 ;
      RECT 70.535 2.116 70.555 2.308 ;
      RECT 70.53 2.127 70.535 2.318 ;
      RECT 70.51 2.14 70.53 2.328 ;
      RECT 70.505 2.15 70.51 2.338 ;
      RECT 70.49 2.155 70.505 2.347 ;
      RECT 70.48 2.165 70.49 2.358 ;
      RECT 70.45 2.182 70.48 2.375 ;
      RECT 70.44 2.2 70.45 2.393 ;
      RECT 70.425 2.211 70.44 2.404 ;
      RECT 70.385 2.235 70.425 2.42 ;
      RECT 70.35 2.269 70.385 2.437 ;
      RECT 70.32 2.292 70.35 2.449 ;
      RECT 70.305 2.302 70.32 2.458 ;
      RECT 70.265 2.312 70.305 2.469 ;
      RECT 70.245 2.323 70.265 2.481 ;
      RECT 70.24 2.327 70.245 2.488 ;
      RECT 70.225 2.331 70.24 2.493 ;
      RECT 70.215 2.336 70.225 2.498 ;
      RECT 70.21 2.339 70.215 2.501 ;
      RECT 70.18 2.345 70.21 2.508 ;
      RECT 70.145 2.355 70.18 2.522 ;
      RECT 70.085 2.37 70.145 2.542 ;
      RECT 70.03 2.39 70.085 2.566 ;
      RECT 70.001 2.405 70.03 2.584 ;
      RECT 69.915 2.425 70.001 2.609 ;
      RECT 69.91 2.44 69.915 2.629 ;
      RECT 69.9 2.443 69.91 2.63 ;
      RECT 69.875 2.45 69.9 2.715 ;
      RECT 70.29 3.685 70.3 3.875 ;
      RECT 68.55 3.56 68.83 3.84 ;
      RECT 71.595 2.5 71.6 2.985 ;
      RECT 71.49 2.5 71.55 2.76 ;
      RECT 71.815 3.47 71.82 3.545 ;
      RECT 71.805 3.337 71.815 3.58 ;
      RECT 71.795 3.172 71.805 3.601 ;
      RECT 71.79 3.042 71.795 3.617 ;
      RECT 71.78 2.932 71.79 3.633 ;
      RECT 71.775 2.831 71.78 3.65 ;
      RECT 71.77 2.813 71.775 3.66 ;
      RECT 71.765 2.795 71.77 3.67 ;
      RECT 71.755 2.77 71.765 3.685 ;
      RECT 71.75 2.75 71.755 3.7 ;
      RECT 71.73 2.5 71.75 3.725 ;
      RECT 71.715 2.5 71.73 3.758 ;
      RECT 71.685 2.5 71.715 3.78 ;
      RECT 71.665 2.5 71.685 3.794 ;
      RECT 71.645 2.5 71.665 3.31 ;
      RECT 71.66 3.377 71.665 3.799 ;
      RECT 71.655 3.407 71.66 3.801 ;
      RECT 71.65 3.42 71.655 3.804 ;
      RECT 71.645 3.43 71.65 3.808 ;
      RECT 71.64 2.5 71.645 3.228 ;
      RECT 71.64 3.44 71.645 3.81 ;
      RECT 71.635 2.5 71.64 3.205 ;
      RECT 71.625 3.462 71.64 3.81 ;
      RECT 71.62 2.5 71.635 3.15 ;
      RECT 71.615 3.487 71.625 3.81 ;
      RECT 71.615 2.5 71.62 3.095 ;
      RECT 71.605 2.5 71.615 3.043 ;
      RECT 71.61 3.5 71.615 3.811 ;
      RECT 71.605 3.512 71.61 3.812 ;
      RECT 71.6 2.5 71.605 3.003 ;
      RECT 71.6 3.525 71.605 3.813 ;
      RECT 71.585 3.54 71.6 3.814 ;
      RECT 71.59 2.5 71.595 2.965 ;
      RECT 71.585 2.5 71.59 2.93 ;
      RECT 71.58 2.5 71.585 2.905 ;
      RECT 71.575 3.567 71.585 3.816 ;
      RECT 71.57 2.5 71.58 2.863 ;
      RECT 71.57 3.585 71.575 3.817 ;
      RECT 71.565 2.5 71.57 2.823 ;
      RECT 71.565 3.592 71.57 3.818 ;
      RECT 71.56 2.5 71.565 2.795 ;
      RECT 71.555 3.61 71.565 3.819 ;
      RECT 71.55 2.5 71.56 2.775 ;
      RECT 71.545 3.63 71.555 3.821 ;
      RECT 71.535 3.647 71.545 3.822 ;
      RECT 71.5 3.67 71.535 3.825 ;
      RECT 71.445 3.688 71.5 3.831 ;
      RECT 71.359 3.696 71.445 3.84 ;
      RECT 71.273 3.707 71.359 3.851 ;
      RECT 71.187 3.717 71.273 3.862 ;
      RECT 71.101 3.727 71.187 3.874 ;
      RECT 71.015 3.737 71.101 3.885 ;
      RECT 70.995 3.743 71.015 3.891 ;
      RECT 70.915 3.745 70.995 3.895 ;
      RECT 70.91 3.744 70.915 3.9 ;
      RECT 70.902 3.743 70.91 3.9 ;
      RECT 70.816 3.739 70.902 3.898 ;
      RECT 70.73 3.731 70.816 3.895 ;
      RECT 70.644 3.722 70.73 3.891 ;
      RECT 70.558 3.714 70.644 3.888 ;
      RECT 70.472 3.706 70.558 3.884 ;
      RECT 70.386 3.697 70.472 3.881 ;
      RECT 70.3 3.689 70.386 3.877 ;
      RECT 70.245 3.682 70.29 3.875 ;
      RECT 70.16 3.675 70.245 3.873 ;
      RECT 70.086 3.667 70.16 3.869 ;
      RECT 70 3.659 70.086 3.866 ;
      RECT 69.997 3.655 70 3.864 ;
      RECT 69.911 3.651 69.997 3.863 ;
      RECT 69.825 3.643 69.911 3.86 ;
      RECT 69.74 3.638 69.825 3.857 ;
      RECT 69.654 3.635 69.74 3.854 ;
      RECT 69.568 3.633 69.654 3.851 ;
      RECT 69.482 3.63 69.568 3.848 ;
      RECT 69.396 3.627 69.482 3.845 ;
      RECT 69.31 3.624 69.396 3.842 ;
      RECT 69.234 3.622 69.31 3.839 ;
      RECT 69.148 3.619 69.234 3.836 ;
      RECT 69.062 3.616 69.148 3.834 ;
      RECT 68.976 3.614 69.062 3.831 ;
      RECT 68.89 3.611 68.976 3.828 ;
      RECT 68.83 3.602 68.89 3.826 ;
      RECT 71.34 3.22 71.415 3.48 ;
      RECT 71.32 3.2 71.325 3.48 ;
      RECT 70.64 2.985 70.745 3.28 ;
      RECT 65.085 2.96 65.155 3.22 ;
      RECT 70.98 2.835 70.985 3.206 ;
      RECT 70.97 2.89 70.975 3.206 ;
      RECT 71.275 2.06 71.335 2.32 ;
      RECT 71.33 3.215 71.34 3.48 ;
      RECT 71.325 3.205 71.33 3.48 ;
      RECT 71.245 3.152 71.32 3.48 ;
      RECT 71.27 2.06 71.275 2.34 ;
      RECT 71.26 2.06 71.27 2.36 ;
      RECT 71.245 2.06 71.26 2.39 ;
      RECT 71.23 2.06 71.245 2.433 ;
      RECT 71.225 3.095 71.245 3.48 ;
      RECT 71.215 2.06 71.23 2.47 ;
      RECT 71.21 3.075 71.225 3.48 ;
      RECT 71.21 2.06 71.215 2.493 ;
      RECT 71.2 2.06 71.21 2.518 ;
      RECT 71.17 3.042 71.21 3.48 ;
      RECT 71.175 2.06 71.2 2.568 ;
      RECT 71.17 2.06 71.175 2.623 ;
      RECT 71.165 2.06 71.17 2.665 ;
      RECT 71.155 3.005 71.17 3.48 ;
      RECT 71.16 2.06 71.165 2.708 ;
      RECT 71.155 2.06 71.16 2.773 ;
      RECT 71.15 2.06 71.155 2.795 ;
      RECT 71.15 2.993 71.155 3.345 ;
      RECT 71.145 2.06 71.15 2.863 ;
      RECT 71.145 2.985 71.15 3.328 ;
      RECT 71.14 2.06 71.145 2.908 ;
      RECT 71.135 2.967 71.145 3.305 ;
      RECT 71.135 2.06 71.14 2.945 ;
      RECT 71.125 2.06 71.135 3.285 ;
      RECT 71.12 2.06 71.125 3.268 ;
      RECT 71.115 2.06 71.12 3.253 ;
      RECT 71.11 2.06 71.115 3.238 ;
      RECT 71.09 2.06 71.11 3.228 ;
      RECT 71.085 2.06 71.09 3.218 ;
      RECT 71.075 2.06 71.085 3.214 ;
      RECT 71.07 2.337 71.075 3.213 ;
      RECT 71.065 2.36 71.07 3.212 ;
      RECT 71.06 2.39 71.065 3.211 ;
      RECT 71.055 2.417 71.06 3.21 ;
      RECT 71.05 2.445 71.055 3.21 ;
      RECT 71.045 2.472 71.05 3.21 ;
      RECT 71.04 2.492 71.045 3.21 ;
      RECT 71.035 2.52 71.04 3.21 ;
      RECT 71.025 2.562 71.035 3.21 ;
      RECT 71.015 2.607 71.025 3.209 ;
      RECT 71.01 2.66 71.015 3.208 ;
      RECT 71.005 2.692 71.01 3.207 ;
      RECT 71 2.712 71.005 3.206 ;
      RECT 70.995 2.75 71 3.206 ;
      RECT 70.99 2.772 70.995 3.206 ;
      RECT 70.985 2.797 70.99 3.206 ;
      RECT 70.975 2.862 70.98 3.206 ;
      RECT 70.96 2.922 70.97 3.206 ;
      RECT 70.945 2.932 70.96 3.206 ;
      RECT 70.925 2.942 70.945 3.206 ;
      RECT 70.895 2.947 70.925 3.203 ;
      RECT 70.835 2.957 70.895 3.2 ;
      RECT 70.815 2.966 70.835 3.205 ;
      RECT 70.79 2.972 70.815 3.218 ;
      RECT 70.77 2.977 70.79 3.233 ;
      RECT 70.745 2.982 70.77 3.28 ;
      RECT 70.616 2.984 70.64 3.28 ;
      RECT 70.53 2.979 70.616 3.28 ;
      RECT 70.49 2.976 70.53 3.28 ;
      RECT 70.44 2.978 70.49 3.26 ;
      RECT 70.41 2.982 70.44 3.26 ;
      RECT 70.331 2.992 70.41 3.26 ;
      RECT 70.245 3.007 70.331 3.261 ;
      RECT 70.195 3.017 70.245 3.262 ;
      RECT 70.187 3.02 70.195 3.262 ;
      RECT 70.101 3.022 70.187 3.263 ;
      RECT 70.015 3.026 70.101 3.263 ;
      RECT 69.929 3.03 70.015 3.264 ;
      RECT 69.843 3.033 69.929 3.265 ;
      RECT 69.757 3.037 69.843 3.265 ;
      RECT 69.671 3.041 69.757 3.266 ;
      RECT 69.585 3.044 69.671 3.267 ;
      RECT 69.499 3.048 69.585 3.267 ;
      RECT 69.413 3.052 69.499 3.268 ;
      RECT 69.327 3.056 69.413 3.269 ;
      RECT 69.241 3.059 69.327 3.269 ;
      RECT 69.155 3.063 69.241 3.27 ;
      RECT 69.125 3.065 69.155 3.27 ;
      RECT 69.039 3.068 69.125 3.271 ;
      RECT 68.953 3.072 69.039 3.272 ;
      RECT 68.867 3.076 68.953 3.273 ;
      RECT 68.781 3.079 68.867 3.273 ;
      RECT 68.695 3.083 68.781 3.274 ;
      RECT 68.66 3.088 68.695 3.275 ;
      RECT 68.605 3.098 68.66 3.282 ;
      RECT 68.58 3.11 68.605 3.292 ;
      RECT 68.545 3.123 68.58 3.3 ;
      RECT 68.505 3.14 68.545 3.323 ;
      RECT 68.485 3.153 68.505 3.35 ;
      RECT 68.455 3.165 68.485 3.378 ;
      RECT 68.45 3.173 68.455 3.398 ;
      RECT 68.445 3.176 68.45 3.408 ;
      RECT 68.395 3.188 68.445 3.442 ;
      RECT 68.385 3.203 68.395 3.475 ;
      RECT 68.375 3.209 68.385 3.488 ;
      RECT 68.365 3.216 68.375 3.5 ;
      RECT 68.34 3.229 68.365 3.518 ;
      RECT 68.325 3.244 68.34 3.54 ;
      RECT 68.315 3.252 68.325 3.556 ;
      RECT 68.3 3.261 68.315 3.571 ;
      RECT 68.29 3.271 68.3 3.585 ;
      RECT 68.271 3.284 68.29 3.602 ;
      RECT 68.185 3.329 68.271 3.667 ;
      RECT 68.17 3.374 68.185 3.725 ;
      RECT 68.165 3.383 68.17 3.738 ;
      RECT 68.155 3.39 68.165 3.743 ;
      RECT 68.15 3.395 68.155 3.747 ;
      RECT 68.13 3.405 68.15 3.754 ;
      RECT 68.105 3.425 68.13 3.768 ;
      RECT 68.07 3.45 68.105 3.788 ;
      RECT 68.055 3.473 68.07 3.803 ;
      RECT 68.045 3.483 68.055 3.808 ;
      RECT 68.035 3.491 68.045 3.815 ;
      RECT 68.025 3.5 68.035 3.821 ;
      RECT 68.005 3.512 68.025 3.823 ;
      RECT 67.995 3.525 68.005 3.825 ;
      RECT 67.97 3.54 67.995 3.828 ;
      RECT 67.95 3.557 67.97 3.832 ;
      RECT 67.91 3.585 67.95 3.838 ;
      RECT 67.845 3.632 67.91 3.847 ;
      RECT 67.83 3.665 67.845 3.855 ;
      RECT 67.825 3.672 67.83 3.857 ;
      RECT 67.775 3.697 67.825 3.862 ;
      RECT 67.76 3.721 67.775 3.869 ;
      RECT 67.71 3.726 67.76 3.87 ;
      RECT 67.624 3.73 67.71 3.87 ;
      RECT 67.538 3.73 67.624 3.87 ;
      RECT 67.452 3.73 67.538 3.871 ;
      RECT 67.366 3.73 67.452 3.871 ;
      RECT 67.28 3.73 67.366 3.871 ;
      RECT 67.214 3.73 67.28 3.871 ;
      RECT 67.128 3.73 67.214 3.872 ;
      RECT 67.042 3.73 67.128 3.872 ;
      RECT 66.956 3.731 67.042 3.873 ;
      RECT 66.87 3.731 66.956 3.873 ;
      RECT 66.784 3.731 66.87 3.873 ;
      RECT 66.698 3.731 66.784 3.874 ;
      RECT 66.612 3.731 66.698 3.874 ;
      RECT 66.526 3.732 66.612 3.875 ;
      RECT 66.44 3.732 66.526 3.875 ;
      RECT 66.42 3.732 66.44 3.875 ;
      RECT 66.334 3.732 66.42 3.875 ;
      RECT 66.248 3.732 66.334 3.875 ;
      RECT 66.162 3.733 66.248 3.875 ;
      RECT 66.076 3.733 66.162 3.875 ;
      RECT 65.99 3.733 66.076 3.875 ;
      RECT 65.904 3.734 65.99 3.875 ;
      RECT 65.818 3.734 65.904 3.875 ;
      RECT 65.732 3.734 65.818 3.875 ;
      RECT 65.646 3.734 65.732 3.875 ;
      RECT 65.56 3.735 65.646 3.875 ;
      RECT 65.51 3.732 65.56 3.875 ;
      RECT 65.5 3.73 65.51 3.874 ;
      RECT 65.496 3.73 65.5 3.873 ;
      RECT 65.41 3.725 65.496 3.868 ;
      RECT 65.388 3.718 65.41 3.862 ;
      RECT 65.302 3.709 65.388 3.856 ;
      RECT 65.216 3.696 65.302 3.847 ;
      RECT 65.13 3.682 65.216 3.837 ;
      RECT 65.085 3.672 65.13 3.83 ;
      RECT 65.065 2.96 65.085 3.238 ;
      RECT 65.065 3.665 65.085 3.826 ;
      RECT 65.035 2.96 65.065 3.26 ;
      RECT 65.025 3.632 65.065 3.823 ;
      RECT 65.02 2.96 65.035 3.28 ;
      RECT 65.02 3.597 65.025 3.821 ;
      RECT 65.015 2.96 65.02 3.405 ;
      RECT 65.015 3.557 65.02 3.821 ;
      RECT 65.005 2.96 65.015 3.821 ;
      RECT 64.93 2.96 65.005 3.815 ;
      RECT 64.9 2.96 64.93 3.805 ;
      RECT 64.895 2.96 64.9 3.797 ;
      RECT 64.89 3.002 64.895 3.79 ;
      RECT 64.88 3.071 64.89 3.781 ;
      RECT 64.875 3.141 64.88 3.733 ;
      RECT 64.87 3.205 64.875 3.63 ;
      RECT 64.865 3.24 64.87 3.585 ;
      RECT 64.863 3.277 64.865 3.477 ;
      RECT 64.86 3.285 64.863 3.47 ;
      RECT 64.855 3.35 64.86 3.413 ;
      RECT 68.93 2.44 69.21 2.72 ;
      RECT 68.92 2.44 69.21 2.583 ;
      RECT 68.875 2.305 69.135 2.565 ;
      RECT 68.875 2.42 69.19 2.565 ;
      RECT 68.875 2.39 69.185 2.565 ;
      RECT 68.875 2.377 69.175 2.565 ;
      RECT 68.875 2.367 69.17 2.565 ;
      RECT 64.85 2.35 65.11 2.61 ;
      RECT 68.62 1.9 68.88 2.16 ;
      RECT 68.61 1.925 68.88 2.12 ;
      RECT 68.605 1.925 68.61 2.119 ;
      RECT 68.535 1.92 68.605 2.111 ;
      RECT 68.45 1.907 68.535 2.094 ;
      RECT 68.446 1.899 68.45 2.084 ;
      RECT 68.36 1.892 68.446 2.074 ;
      RECT 68.351 1.884 68.36 2.064 ;
      RECT 68.265 1.877 68.351 2.052 ;
      RECT 68.245 1.868 68.265 2.038 ;
      RECT 68.19 1.863 68.245 2.03 ;
      RECT 68.18 1.857 68.19 2.024 ;
      RECT 68.16 1.855 68.18 2.02 ;
      RECT 68.152 1.854 68.16 2.016 ;
      RECT 68.066 1.846 68.152 2.005 ;
      RECT 67.98 1.832 68.066 1.985 ;
      RECT 67.92 1.82 67.98 1.97 ;
      RECT 67.91 1.815 67.92 1.965 ;
      RECT 67.86 1.815 67.91 1.967 ;
      RECT 67.813 1.817 67.86 1.971 ;
      RECT 67.727 1.824 67.813 1.976 ;
      RECT 67.641 1.832 67.727 1.982 ;
      RECT 67.555 1.841 67.641 1.988 ;
      RECT 67.496 1.847 67.555 1.993 ;
      RECT 67.41 1.852 67.496 1.999 ;
      RECT 67.335 1.857 67.41 2.005 ;
      RECT 67.296 1.859 67.335 2.01 ;
      RECT 67.21 1.856 67.296 2.015 ;
      RECT 67.125 1.854 67.21 2.022 ;
      RECT 67.093 1.853 67.125 2.025 ;
      RECT 67.007 1.852 67.093 2.026 ;
      RECT 66.921 1.851 67.007 2.027 ;
      RECT 66.835 1.85 66.921 2.027 ;
      RECT 66.749 1.849 66.835 2.028 ;
      RECT 66.663 1.848 66.749 2.029 ;
      RECT 66.577 1.847 66.663 2.03 ;
      RECT 66.491 1.846 66.577 2.03 ;
      RECT 66.405 1.845 66.491 2.031 ;
      RECT 66.355 1.845 66.405 2.032 ;
      RECT 66.341 1.846 66.355 2.032 ;
      RECT 66.255 1.853 66.341 2.033 ;
      RECT 66.181 1.864 66.255 2.034 ;
      RECT 66.095 1.873 66.181 2.035 ;
      RECT 66.06 1.88 66.095 2.05 ;
      RECT 66.035 1.883 66.06 2.08 ;
      RECT 66.01 1.892 66.035 2.109 ;
      RECT 66 1.903 66.01 2.129 ;
      RECT 65.99 1.911 66 2.143 ;
      RECT 65.985 1.917 65.99 2.153 ;
      RECT 65.96 1.934 65.985 2.17 ;
      RECT 65.945 1.956 65.96 2.198 ;
      RECT 65.915 1.982 65.945 2.228 ;
      RECT 65.895 2.011 65.915 2.258 ;
      RECT 65.89 2.026 65.895 2.275 ;
      RECT 65.87 2.041 65.89 2.29 ;
      RECT 65.86 2.059 65.87 2.308 ;
      RECT 65.85 2.07 65.86 2.323 ;
      RECT 65.8 2.102 65.85 2.349 ;
      RECT 65.795 2.132 65.8 2.369 ;
      RECT 65.785 2.145 65.795 2.375 ;
      RECT 65.776 2.155 65.785 2.383 ;
      RECT 65.765 2.166 65.776 2.391 ;
      RECT 65.76 2.176 65.765 2.397 ;
      RECT 65.745 2.197 65.76 2.404 ;
      RECT 65.73 2.227 65.745 2.412 ;
      RECT 65.695 2.257 65.73 2.418 ;
      RECT 65.67 2.275 65.695 2.425 ;
      RECT 65.62 2.283 65.67 2.434 ;
      RECT 65.595 2.288 65.62 2.443 ;
      RECT 65.54 2.294 65.595 2.453 ;
      RECT 65.535 2.299 65.54 2.461 ;
      RECT 65.521 2.302 65.535 2.463 ;
      RECT 65.435 2.314 65.521 2.475 ;
      RECT 65.425 2.326 65.435 2.488 ;
      RECT 65.34 2.339 65.425 2.5 ;
      RECT 65.296 2.356 65.34 2.514 ;
      RECT 65.21 2.373 65.296 2.53 ;
      RECT 65.18 2.387 65.21 2.544 ;
      RECT 65.17 2.392 65.18 2.549 ;
      RECT 65.11 2.395 65.17 2.558 ;
      RECT 68 2.665 68.26 2.925 ;
      RECT 68 2.665 68.28 2.778 ;
      RECT 68 2.665 68.305 2.745 ;
      RECT 68 2.665 68.31 2.725 ;
      RECT 68.05 2.44 68.33 2.72 ;
      RECT 67.605 3.175 67.865 3.435 ;
      RECT 67.595 3.032 67.79 3.373 ;
      RECT 67.59 3.14 67.805 3.365 ;
      RECT 67.585 3.19 67.865 3.355 ;
      RECT 67.575 3.267 67.865 3.34 ;
      RECT 67.595 3.115 67.805 3.373 ;
      RECT 67.605 2.99 67.79 3.435 ;
      RECT 67.605 2.885 67.77 3.435 ;
      RECT 67.615 2.872 67.77 3.435 ;
      RECT 67.615 2.83 67.76 3.435 ;
      RECT 67.62 2.755 67.76 3.435 ;
      RECT 67.65 2.405 67.76 3.435 ;
      RECT 67.655 2.135 67.78 2.758 ;
      RECT 67.625 2.71 67.78 2.758 ;
      RECT 67.64 2.512 67.76 3.435 ;
      RECT 67.63 2.622 67.78 2.758 ;
      RECT 67.655 2.135 67.795 2.615 ;
      RECT 67.655 2.135 67.815 2.49 ;
      RECT 67.62 2.135 67.88 2.395 ;
      RECT 67.09 2.44 67.37 2.72 ;
      RECT 67.075 2.44 67.37 2.7 ;
      RECT 65.13 3.305 65.39 3.565 ;
      RECT 66.915 3.16 67.175 3.42 ;
      RECT 66.895 3.18 67.175 3.395 ;
      RECT 66.852 3.18 66.895 3.394 ;
      RECT 66.766 3.181 66.852 3.391 ;
      RECT 66.68 3.182 66.766 3.387 ;
      RECT 66.605 3.184 66.68 3.384 ;
      RECT 66.582 3.185 66.605 3.382 ;
      RECT 66.496 3.186 66.582 3.38 ;
      RECT 66.41 3.187 66.496 3.377 ;
      RECT 66.386 3.188 66.41 3.375 ;
      RECT 66.3 3.19 66.386 3.372 ;
      RECT 66.215 3.192 66.3 3.373 ;
      RECT 66.158 3.193 66.215 3.379 ;
      RECT 66.072 3.195 66.158 3.389 ;
      RECT 65.986 3.198 66.072 3.402 ;
      RECT 65.9 3.2 65.986 3.414 ;
      RECT 65.886 3.201 65.9 3.421 ;
      RECT 65.8 3.202 65.886 3.429 ;
      RECT 65.76 3.204 65.8 3.438 ;
      RECT 65.751 3.205 65.76 3.441 ;
      RECT 65.665 3.213 65.751 3.447 ;
      RECT 65.645 3.222 65.665 3.455 ;
      RECT 65.56 3.237 65.645 3.463 ;
      RECT 65.5 3.26 65.56 3.474 ;
      RECT 65.49 3.272 65.5 3.479 ;
      RECT 65.45 3.282 65.49 3.483 ;
      RECT 65.395 3.299 65.45 3.491 ;
      RECT 65.39 3.309 65.395 3.495 ;
      RECT 66.456 2.44 66.515 2.837 ;
      RECT 66.37 2.44 66.575 2.828 ;
      RECT 66.365 2.47 66.575 2.823 ;
      RECT 66.331 2.47 66.575 2.821 ;
      RECT 66.245 2.47 66.575 2.815 ;
      RECT 66.2 2.47 66.595 2.793 ;
      RECT 66.2 2.47 66.615 2.748 ;
      RECT 66.16 2.47 66.615 2.738 ;
      RECT 66.37 2.44 66.65 2.72 ;
      RECT 66.105 2.44 66.365 2.7 ;
      RECT 65.29 1.92 65.55 2.18 ;
      RECT 65.345 1.88 65.65 2.16 ;
      RECT 65.345 1.855 65.52 2.18 ;
      RECT 59.67 6.28 59.99 6.605 ;
      RECT 59.7 5.695 59.87 6.605 ;
      RECT 59.7 5.695 59.875 6.045 ;
      RECT 59.7 5.695 60.675 5.87 ;
      RECT 60.5 1.965 60.675 5.87 ;
      RECT 56.72 2.84 57 3.28 ;
      RECT 56.72 2.84 57.005 3.238 ;
      RECT 56.72 2.84 57.01 3.135 ;
      RECT 56.72 2.84 57.012 3.015 ;
      RECT 56.72 2.84 57.645 3.01 ;
      RECT 57.475 2.025 57.645 3.01 ;
      RECT 56.72 2.805 56.98 3.28 ;
      RECT 60.445 1.965 60.795 2.315 ;
      RECT 57.475 2.025 60.795 2.195 ;
      RECT 59.365 0.915 59.535 2.195 ;
      RECT 46.98 0.885 47.33 1.235 ;
      RECT 46.98 0.915 59.535 1.085 ;
      RECT 60.47 6.655 60.795 6.98 ;
      RECT 59.355 6.745 60.795 6.915 ;
      RECT 59.355 2.395 59.515 6.915 ;
      RECT 59.67 2.365 59.99 2.685 ;
      RECT 59.355 2.395 59.99 2.565 ;
      RECT 58.62 5.855 58.97 6.205 ;
      RECT 58.69 2.705 58.865 6.205 ;
      RECT 58.615 2.705 58.965 3.055 ;
      RECT 48.08 3 48.36 3.28 ;
      RECT 48.05 3 48.36 3.265 ;
      RECT 48.045 2.963 48.305 3.263 ;
      RECT 48.04 2.964 48.305 3.257 ;
      RECT 48.035 2.967 48.305 3.25 ;
      RECT 48.03 3 48.36 3.243 ;
      RECT 48 2.97 48.305 3.23 ;
      RECT 48 2.997 48.325 3.23 ;
      RECT 48 2.987 48.32 3.23 ;
      RECT 48 2.972 48.315 3.23 ;
      RECT 48.1 2.962 48.305 3.28 ;
      RECT 48.1 2.957 48.295 3.28 ;
      RECT 48.1 2.955 48.28 3.28 ;
      RECT 48.1 1.42 48.275 3.28 ;
      RECT 58.01 1.34 58.36 1.69 ;
      RECT 48.1 1.42 58.36 1.595 ;
      RECT 53.79 2.455 54.025 2.715 ;
      RECT 56.935 2.235 57.1 2.495 ;
      RECT 56.84 2.225 56.855 2.495 ;
      RECT 55.44 1.795 55.48 1.935 ;
      RECT 56.855 2.23 56.935 2.495 ;
      RECT 56.8 2.225 56.84 2.461 ;
      RECT 56.786 2.225 56.8 2.461 ;
      RECT 56.7 2.23 56.786 2.463 ;
      RECT 56.655 2.237 56.7 2.465 ;
      RECT 56.625 2.237 56.655 2.467 ;
      RECT 56.6 2.232 56.625 2.469 ;
      RECT 56.57 2.228 56.6 2.478 ;
      RECT 56.56 2.225 56.57 2.49 ;
      RECT 56.555 2.225 56.56 2.498 ;
      RECT 56.55 2.225 56.555 2.503 ;
      RECT 56.54 2.224 56.55 2.513 ;
      RECT 56.535 2.223 56.54 2.523 ;
      RECT 56.52 2.222 56.535 2.528 ;
      RECT 56.492 2.219 56.52 2.555 ;
      RECT 56.406 2.211 56.492 2.555 ;
      RECT 56.32 2.2 56.406 2.555 ;
      RECT 56.28 2.185 56.32 2.555 ;
      RECT 56.24 2.159 56.28 2.555 ;
      RECT 56.235 2.141 56.24 2.367 ;
      RECT 56.225 2.137 56.235 2.357 ;
      RECT 56.21 2.127 56.225 2.344 ;
      RECT 56.19 2.111 56.21 2.329 ;
      RECT 56.175 2.096 56.19 2.314 ;
      RECT 56.165 2.085 56.175 2.304 ;
      RECT 56.14 2.069 56.165 2.293 ;
      RECT 56.135 2.056 56.14 2.283 ;
      RECT 56.13 2.052 56.135 2.278 ;
      RECT 56.075 2.038 56.13 2.256 ;
      RECT 56.036 2.019 56.075 2.22 ;
      RECT 55.95 1.993 56.036 2.173 ;
      RECT 55.946 1.975 55.95 2.139 ;
      RECT 55.86 1.956 55.946 2.117 ;
      RECT 55.855 1.938 55.86 2.095 ;
      RECT 55.85 1.936 55.855 2.093 ;
      RECT 55.84 1.935 55.85 2.088 ;
      RECT 55.78 1.922 55.84 2.074 ;
      RECT 55.735 1.9 55.78 2.053 ;
      RECT 55.675 1.877 55.735 2.032 ;
      RECT 55.611 1.852 55.675 2.007 ;
      RECT 55.525 1.822 55.611 1.976 ;
      RECT 55.51 1.802 55.525 1.955 ;
      RECT 55.48 1.797 55.51 1.946 ;
      RECT 55.427 1.795 55.44 1.935 ;
      RECT 55.341 1.795 55.427 1.937 ;
      RECT 55.255 1.795 55.341 1.939 ;
      RECT 55.235 1.795 55.255 1.943 ;
      RECT 55.19 1.797 55.235 1.954 ;
      RECT 55.15 1.807 55.19 1.97 ;
      RECT 55.146 1.816 55.15 1.978 ;
      RECT 55.06 1.836 55.146 1.994 ;
      RECT 55.05 1.855 55.06 2.012 ;
      RECT 55.045 1.857 55.05 2.015 ;
      RECT 55.035 1.861 55.045 2.018 ;
      RECT 55.015 1.866 55.035 2.028 ;
      RECT 54.985 1.876 55.015 2.048 ;
      RECT 54.98 1.883 54.985 2.062 ;
      RECT 54.97 1.887 54.98 2.069 ;
      RECT 54.955 1.895 54.97 2.08 ;
      RECT 54.945 1.905 54.955 2.091 ;
      RECT 54.935 1.912 54.945 2.099 ;
      RECT 54.91 1.925 54.935 2.114 ;
      RECT 54.846 1.961 54.91 2.153 ;
      RECT 54.76 2.024 54.846 2.217 ;
      RECT 54.725 2.075 54.76 2.27 ;
      RECT 54.72 2.092 54.725 2.287 ;
      RECT 54.705 2.101 54.72 2.294 ;
      RECT 54.685 2.116 54.705 2.308 ;
      RECT 54.68 2.127 54.685 2.318 ;
      RECT 54.66 2.14 54.68 2.328 ;
      RECT 54.655 2.15 54.66 2.338 ;
      RECT 54.64 2.155 54.655 2.347 ;
      RECT 54.63 2.165 54.64 2.358 ;
      RECT 54.6 2.182 54.63 2.375 ;
      RECT 54.59 2.2 54.6 2.393 ;
      RECT 54.575 2.211 54.59 2.404 ;
      RECT 54.535 2.235 54.575 2.42 ;
      RECT 54.5 2.269 54.535 2.437 ;
      RECT 54.47 2.292 54.5 2.449 ;
      RECT 54.455 2.302 54.47 2.458 ;
      RECT 54.415 2.312 54.455 2.469 ;
      RECT 54.395 2.323 54.415 2.481 ;
      RECT 54.39 2.327 54.395 2.488 ;
      RECT 54.375 2.331 54.39 2.493 ;
      RECT 54.365 2.336 54.375 2.498 ;
      RECT 54.36 2.339 54.365 2.501 ;
      RECT 54.33 2.345 54.36 2.508 ;
      RECT 54.295 2.355 54.33 2.522 ;
      RECT 54.235 2.37 54.295 2.542 ;
      RECT 54.18 2.39 54.235 2.566 ;
      RECT 54.151 2.405 54.18 2.584 ;
      RECT 54.065 2.425 54.151 2.609 ;
      RECT 54.06 2.44 54.065 2.629 ;
      RECT 54.05 2.443 54.06 2.63 ;
      RECT 54.025 2.45 54.05 2.715 ;
      RECT 54.44 3.685 54.45 3.875 ;
      RECT 52.7 3.56 52.98 3.84 ;
      RECT 55.745 2.5 55.75 2.985 ;
      RECT 55.64 2.5 55.7 2.76 ;
      RECT 55.965 3.47 55.97 3.545 ;
      RECT 55.955 3.337 55.965 3.58 ;
      RECT 55.945 3.172 55.955 3.601 ;
      RECT 55.94 3.042 55.945 3.617 ;
      RECT 55.93 2.932 55.94 3.633 ;
      RECT 55.925 2.831 55.93 3.65 ;
      RECT 55.92 2.813 55.925 3.66 ;
      RECT 55.915 2.795 55.92 3.67 ;
      RECT 55.905 2.77 55.915 3.685 ;
      RECT 55.9 2.75 55.905 3.7 ;
      RECT 55.88 2.5 55.9 3.725 ;
      RECT 55.865 2.5 55.88 3.758 ;
      RECT 55.835 2.5 55.865 3.78 ;
      RECT 55.815 2.5 55.835 3.794 ;
      RECT 55.795 2.5 55.815 3.31 ;
      RECT 55.81 3.377 55.815 3.799 ;
      RECT 55.805 3.407 55.81 3.801 ;
      RECT 55.8 3.42 55.805 3.804 ;
      RECT 55.795 3.43 55.8 3.808 ;
      RECT 55.79 2.5 55.795 3.228 ;
      RECT 55.79 3.44 55.795 3.81 ;
      RECT 55.785 2.5 55.79 3.205 ;
      RECT 55.775 3.462 55.79 3.81 ;
      RECT 55.77 2.5 55.785 3.15 ;
      RECT 55.765 3.487 55.775 3.81 ;
      RECT 55.765 2.5 55.77 3.095 ;
      RECT 55.755 2.5 55.765 3.043 ;
      RECT 55.76 3.5 55.765 3.811 ;
      RECT 55.755 3.512 55.76 3.812 ;
      RECT 55.75 2.5 55.755 3.003 ;
      RECT 55.75 3.525 55.755 3.813 ;
      RECT 55.735 3.54 55.75 3.814 ;
      RECT 55.74 2.5 55.745 2.965 ;
      RECT 55.735 2.5 55.74 2.93 ;
      RECT 55.73 2.5 55.735 2.905 ;
      RECT 55.725 3.567 55.735 3.816 ;
      RECT 55.72 2.5 55.73 2.863 ;
      RECT 55.72 3.585 55.725 3.817 ;
      RECT 55.715 2.5 55.72 2.823 ;
      RECT 55.715 3.592 55.72 3.818 ;
      RECT 55.71 2.5 55.715 2.795 ;
      RECT 55.705 3.61 55.715 3.819 ;
      RECT 55.7 2.5 55.71 2.775 ;
      RECT 55.695 3.63 55.705 3.821 ;
      RECT 55.685 3.647 55.695 3.822 ;
      RECT 55.65 3.67 55.685 3.825 ;
      RECT 55.595 3.688 55.65 3.831 ;
      RECT 55.509 3.696 55.595 3.84 ;
      RECT 55.423 3.707 55.509 3.851 ;
      RECT 55.337 3.717 55.423 3.862 ;
      RECT 55.251 3.727 55.337 3.874 ;
      RECT 55.165 3.737 55.251 3.885 ;
      RECT 55.145 3.743 55.165 3.891 ;
      RECT 55.065 3.745 55.145 3.895 ;
      RECT 55.06 3.744 55.065 3.9 ;
      RECT 55.052 3.743 55.06 3.9 ;
      RECT 54.966 3.739 55.052 3.898 ;
      RECT 54.88 3.731 54.966 3.895 ;
      RECT 54.794 3.722 54.88 3.891 ;
      RECT 54.708 3.714 54.794 3.888 ;
      RECT 54.622 3.706 54.708 3.884 ;
      RECT 54.536 3.697 54.622 3.881 ;
      RECT 54.45 3.689 54.536 3.877 ;
      RECT 54.395 3.682 54.44 3.875 ;
      RECT 54.31 3.675 54.395 3.873 ;
      RECT 54.236 3.667 54.31 3.869 ;
      RECT 54.15 3.659 54.236 3.866 ;
      RECT 54.147 3.655 54.15 3.864 ;
      RECT 54.061 3.651 54.147 3.863 ;
      RECT 53.975 3.643 54.061 3.86 ;
      RECT 53.89 3.638 53.975 3.857 ;
      RECT 53.804 3.635 53.89 3.854 ;
      RECT 53.718 3.633 53.804 3.851 ;
      RECT 53.632 3.63 53.718 3.848 ;
      RECT 53.546 3.627 53.632 3.845 ;
      RECT 53.46 3.624 53.546 3.842 ;
      RECT 53.384 3.622 53.46 3.839 ;
      RECT 53.298 3.619 53.384 3.836 ;
      RECT 53.212 3.616 53.298 3.834 ;
      RECT 53.126 3.614 53.212 3.831 ;
      RECT 53.04 3.611 53.126 3.828 ;
      RECT 52.98 3.602 53.04 3.826 ;
      RECT 55.49 3.22 55.565 3.48 ;
      RECT 55.47 3.2 55.475 3.48 ;
      RECT 54.79 2.985 54.895 3.28 ;
      RECT 49.235 2.96 49.305 3.22 ;
      RECT 55.13 2.835 55.135 3.206 ;
      RECT 55.12 2.89 55.125 3.206 ;
      RECT 55.425 2.06 55.485 2.32 ;
      RECT 55.48 3.215 55.49 3.48 ;
      RECT 55.475 3.205 55.48 3.48 ;
      RECT 55.395 3.152 55.47 3.48 ;
      RECT 55.42 2.06 55.425 2.34 ;
      RECT 55.41 2.06 55.42 2.36 ;
      RECT 55.395 2.06 55.41 2.39 ;
      RECT 55.38 2.06 55.395 2.433 ;
      RECT 55.375 3.095 55.395 3.48 ;
      RECT 55.365 2.06 55.38 2.47 ;
      RECT 55.36 3.075 55.375 3.48 ;
      RECT 55.36 2.06 55.365 2.493 ;
      RECT 55.35 2.06 55.36 2.518 ;
      RECT 55.32 3.042 55.36 3.48 ;
      RECT 55.325 2.06 55.35 2.568 ;
      RECT 55.32 2.06 55.325 2.623 ;
      RECT 55.315 2.06 55.32 2.665 ;
      RECT 55.305 3.005 55.32 3.48 ;
      RECT 55.31 2.06 55.315 2.708 ;
      RECT 55.305 2.06 55.31 2.773 ;
      RECT 55.3 2.06 55.305 2.795 ;
      RECT 55.3 2.993 55.305 3.345 ;
      RECT 55.295 2.06 55.3 2.863 ;
      RECT 55.295 2.985 55.3 3.328 ;
      RECT 55.29 2.06 55.295 2.908 ;
      RECT 55.285 2.967 55.295 3.305 ;
      RECT 55.285 2.06 55.29 2.945 ;
      RECT 55.275 2.06 55.285 3.285 ;
      RECT 55.27 2.06 55.275 3.268 ;
      RECT 55.265 2.06 55.27 3.253 ;
      RECT 55.26 2.06 55.265 3.238 ;
      RECT 55.24 2.06 55.26 3.228 ;
      RECT 55.235 2.06 55.24 3.218 ;
      RECT 55.225 2.06 55.235 3.214 ;
      RECT 55.22 2.337 55.225 3.213 ;
      RECT 55.215 2.36 55.22 3.212 ;
      RECT 55.21 2.39 55.215 3.211 ;
      RECT 55.205 2.417 55.21 3.21 ;
      RECT 55.2 2.445 55.205 3.21 ;
      RECT 55.195 2.472 55.2 3.21 ;
      RECT 55.19 2.492 55.195 3.21 ;
      RECT 55.185 2.52 55.19 3.21 ;
      RECT 55.175 2.562 55.185 3.21 ;
      RECT 55.165 2.607 55.175 3.209 ;
      RECT 55.16 2.66 55.165 3.208 ;
      RECT 55.155 2.692 55.16 3.207 ;
      RECT 55.15 2.712 55.155 3.206 ;
      RECT 55.145 2.75 55.15 3.206 ;
      RECT 55.14 2.772 55.145 3.206 ;
      RECT 55.135 2.797 55.14 3.206 ;
      RECT 55.125 2.862 55.13 3.206 ;
      RECT 55.11 2.922 55.12 3.206 ;
      RECT 55.095 2.932 55.11 3.206 ;
      RECT 55.075 2.942 55.095 3.206 ;
      RECT 55.045 2.947 55.075 3.203 ;
      RECT 54.985 2.957 55.045 3.2 ;
      RECT 54.965 2.966 54.985 3.205 ;
      RECT 54.94 2.972 54.965 3.218 ;
      RECT 54.92 2.977 54.94 3.233 ;
      RECT 54.895 2.982 54.92 3.28 ;
      RECT 54.766 2.984 54.79 3.28 ;
      RECT 54.68 2.979 54.766 3.28 ;
      RECT 54.64 2.976 54.68 3.28 ;
      RECT 54.59 2.978 54.64 3.26 ;
      RECT 54.56 2.982 54.59 3.26 ;
      RECT 54.481 2.992 54.56 3.26 ;
      RECT 54.395 3.007 54.481 3.261 ;
      RECT 54.345 3.017 54.395 3.262 ;
      RECT 54.337 3.02 54.345 3.262 ;
      RECT 54.251 3.022 54.337 3.263 ;
      RECT 54.165 3.026 54.251 3.263 ;
      RECT 54.079 3.03 54.165 3.264 ;
      RECT 53.993 3.033 54.079 3.265 ;
      RECT 53.907 3.037 53.993 3.265 ;
      RECT 53.821 3.041 53.907 3.266 ;
      RECT 53.735 3.044 53.821 3.267 ;
      RECT 53.649 3.048 53.735 3.267 ;
      RECT 53.563 3.052 53.649 3.268 ;
      RECT 53.477 3.056 53.563 3.269 ;
      RECT 53.391 3.059 53.477 3.269 ;
      RECT 53.305 3.063 53.391 3.27 ;
      RECT 53.275 3.065 53.305 3.27 ;
      RECT 53.189 3.068 53.275 3.271 ;
      RECT 53.103 3.072 53.189 3.272 ;
      RECT 53.017 3.076 53.103 3.273 ;
      RECT 52.931 3.079 53.017 3.273 ;
      RECT 52.845 3.083 52.931 3.274 ;
      RECT 52.81 3.088 52.845 3.275 ;
      RECT 52.755 3.098 52.81 3.282 ;
      RECT 52.73 3.11 52.755 3.292 ;
      RECT 52.695 3.123 52.73 3.3 ;
      RECT 52.655 3.14 52.695 3.323 ;
      RECT 52.635 3.153 52.655 3.35 ;
      RECT 52.605 3.165 52.635 3.378 ;
      RECT 52.6 3.173 52.605 3.398 ;
      RECT 52.595 3.176 52.6 3.408 ;
      RECT 52.545 3.188 52.595 3.442 ;
      RECT 52.535 3.203 52.545 3.475 ;
      RECT 52.525 3.209 52.535 3.488 ;
      RECT 52.515 3.216 52.525 3.5 ;
      RECT 52.49 3.229 52.515 3.518 ;
      RECT 52.475 3.244 52.49 3.54 ;
      RECT 52.465 3.252 52.475 3.556 ;
      RECT 52.45 3.261 52.465 3.571 ;
      RECT 52.44 3.271 52.45 3.585 ;
      RECT 52.421 3.284 52.44 3.602 ;
      RECT 52.335 3.329 52.421 3.667 ;
      RECT 52.32 3.374 52.335 3.725 ;
      RECT 52.315 3.383 52.32 3.738 ;
      RECT 52.305 3.39 52.315 3.743 ;
      RECT 52.3 3.395 52.305 3.747 ;
      RECT 52.28 3.405 52.3 3.754 ;
      RECT 52.255 3.425 52.28 3.768 ;
      RECT 52.22 3.45 52.255 3.788 ;
      RECT 52.205 3.473 52.22 3.803 ;
      RECT 52.195 3.483 52.205 3.808 ;
      RECT 52.185 3.491 52.195 3.815 ;
      RECT 52.175 3.5 52.185 3.821 ;
      RECT 52.155 3.512 52.175 3.823 ;
      RECT 52.145 3.525 52.155 3.825 ;
      RECT 52.12 3.54 52.145 3.828 ;
      RECT 52.1 3.557 52.12 3.832 ;
      RECT 52.06 3.585 52.1 3.838 ;
      RECT 51.995 3.632 52.06 3.847 ;
      RECT 51.98 3.665 51.995 3.855 ;
      RECT 51.975 3.672 51.98 3.857 ;
      RECT 51.925 3.697 51.975 3.862 ;
      RECT 51.91 3.721 51.925 3.869 ;
      RECT 51.86 3.726 51.91 3.87 ;
      RECT 51.774 3.73 51.86 3.87 ;
      RECT 51.688 3.73 51.774 3.87 ;
      RECT 51.602 3.73 51.688 3.871 ;
      RECT 51.516 3.73 51.602 3.871 ;
      RECT 51.43 3.73 51.516 3.871 ;
      RECT 51.364 3.73 51.43 3.871 ;
      RECT 51.278 3.73 51.364 3.872 ;
      RECT 51.192 3.73 51.278 3.872 ;
      RECT 51.106 3.731 51.192 3.873 ;
      RECT 51.02 3.731 51.106 3.873 ;
      RECT 50.934 3.731 51.02 3.873 ;
      RECT 50.848 3.731 50.934 3.874 ;
      RECT 50.762 3.731 50.848 3.874 ;
      RECT 50.676 3.732 50.762 3.875 ;
      RECT 50.59 3.732 50.676 3.875 ;
      RECT 50.57 3.732 50.59 3.875 ;
      RECT 50.484 3.732 50.57 3.875 ;
      RECT 50.398 3.732 50.484 3.875 ;
      RECT 50.312 3.733 50.398 3.875 ;
      RECT 50.226 3.733 50.312 3.875 ;
      RECT 50.14 3.733 50.226 3.875 ;
      RECT 50.054 3.734 50.14 3.875 ;
      RECT 49.968 3.734 50.054 3.875 ;
      RECT 49.882 3.734 49.968 3.875 ;
      RECT 49.796 3.734 49.882 3.875 ;
      RECT 49.71 3.735 49.796 3.875 ;
      RECT 49.66 3.732 49.71 3.875 ;
      RECT 49.65 3.73 49.66 3.874 ;
      RECT 49.646 3.73 49.65 3.873 ;
      RECT 49.56 3.725 49.646 3.868 ;
      RECT 49.538 3.718 49.56 3.862 ;
      RECT 49.452 3.709 49.538 3.856 ;
      RECT 49.366 3.696 49.452 3.847 ;
      RECT 49.28 3.682 49.366 3.837 ;
      RECT 49.235 3.672 49.28 3.83 ;
      RECT 49.215 2.96 49.235 3.238 ;
      RECT 49.215 3.665 49.235 3.826 ;
      RECT 49.185 2.96 49.215 3.26 ;
      RECT 49.175 3.632 49.215 3.823 ;
      RECT 49.17 2.96 49.185 3.28 ;
      RECT 49.17 3.597 49.175 3.821 ;
      RECT 49.165 2.96 49.17 3.405 ;
      RECT 49.165 3.557 49.17 3.821 ;
      RECT 49.155 2.96 49.165 3.821 ;
      RECT 49.08 2.96 49.155 3.815 ;
      RECT 49.05 2.96 49.08 3.805 ;
      RECT 49.045 2.96 49.05 3.797 ;
      RECT 49.04 3.002 49.045 3.79 ;
      RECT 49.03 3.071 49.04 3.781 ;
      RECT 49.025 3.141 49.03 3.733 ;
      RECT 49.02 3.205 49.025 3.63 ;
      RECT 49.015 3.24 49.02 3.585 ;
      RECT 49.013 3.277 49.015 3.477 ;
      RECT 49.01 3.285 49.013 3.47 ;
      RECT 49.005 3.35 49.01 3.413 ;
      RECT 53.08 2.44 53.36 2.72 ;
      RECT 53.07 2.44 53.36 2.583 ;
      RECT 53.025 2.305 53.285 2.565 ;
      RECT 53.025 2.42 53.34 2.565 ;
      RECT 53.025 2.39 53.335 2.565 ;
      RECT 53.025 2.377 53.325 2.565 ;
      RECT 53.025 2.367 53.32 2.565 ;
      RECT 49 2.35 49.26 2.61 ;
      RECT 52.77 1.9 53.03 2.16 ;
      RECT 52.76 1.925 53.03 2.12 ;
      RECT 52.755 1.925 52.76 2.119 ;
      RECT 52.685 1.92 52.755 2.111 ;
      RECT 52.6 1.907 52.685 2.094 ;
      RECT 52.596 1.899 52.6 2.084 ;
      RECT 52.51 1.892 52.596 2.074 ;
      RECT 52.501 1.884 52.51 2.064 ;
      RECT 52.415 1.877 52.501 2.052 ;
      RECT 52.395 1.868 52.415 2.038 ;
      RECT 52.34 1.863 52.395 2.03 ;
      RECT 52.33 1.857 52.34 2.024 ;
      RECT 52.31 1.855 52.33 2.02 ;
      RECT 52.302 1.854 52.31 2.016 ;
      RECT 52.216 1.846 52.302 2.005 ;
      RECT 52.13 1.832 52.216 1.985 ;
      RECT 52.07 1.82 52.13 1.97 ;
      RECT 52.06 1.815 52.07 1.965 ;
      RECT 52.01 1.815 52.06 1.967 ;
      RECT 51.963 1.817 52.01 1.971 ;
      RECT 51.877 1.824 51.963 1.976 ;
      RECT 51.791 1.832 51.877 1.982 ;
      RECT 51.705 1.841 51.791 1.988 ;
      RECT 51.646 1.847 51.705 1.993 ;
      RECT 51.56 1.852 51.646 1.999 ;
      RECT 51.485 1.857 51.56 2.005 ;
      RECT 51.446 1.859 51.485 2.01 ;
      RECT 51.36 1.856 51.446 2.015 ;
      RECT 51.275 1.854 51.36 2.022 ;
      RECT 51.243 1.853 51.275 2.025 ;
      RECT 51.157 1.852 51.243 2.026 ;
      RECT 51.071 1.851 51.157 2.027 ;
      RECT 50.985 1.85 51.071 2.027 ;
      RECT 50.899 1.849 50.985 2.028 ;
      RECT 50.813 1.848 50.899 2.029 ;
      RECT 50.727 1.847 50.813 2.03 ;
      RECT 50.641 1.846 50.727 2.03 ;
      RECT 50.555 1.845 50.641 2.031 ;
      RECT 50.505 1.845 50.555 2.032 ;
      RECT 50.491 1.846 50.505 2.032 ;
      RECT 50.405 1.853 50.491 2.033 ;
      RECT 50.331 1.864 50.405 2.034 ;
      RECT 50.245 1.873 50.331 2.035 ;
      RECT 50.21 1.88 50.245 2.05 ;
      RECT 50.185 1.883 50.21 2.08 ;
      RECT 50.16 1.892 50.185 2.109 ;
      RECT 50.15 1.903 50.16 2.129 ;
      RECT 50.14 1.911 50.15 2.143 ;
      RECT 50.135 1.917 50.14 2.153 ;
      RECT 50.11 1.934 50.135 2.17 ;
      RECT 50.095 1.956 50.11 2.198 ;
      RECT 50.065 1.982 50.095 2.228 ;
      RECT 50.045 2.011 50.065 2.258 ;
      RECT 50.04 2.026 50.045 2.275 ;
      RECT 50.02 2.041 50.04 2.29 ;
      RECT 50.01 2.059 50.02 2.308 ;
      RECT 50 2.07 50.01 2.323 ;
      RECT 49.95 2.102 50 2.349 ;
      RECT 49.945 2.132 49.95 2.369 ;
      RECT 49.935 2.145 49.945 2.375 ;
      RECT 49.926 2.155 49.935 2.383 ;
      RECT 49.915 2.166 49.926 2.391 ;
      RECT 49.91 2.176 49.915 2.397 ;
      RECT 49.895 2.197 49.91 2.404 ;
      RECT 49.88 2.227 49.895 2.412 ;
      RECT 49.845 2.257 49.88 2.418 ;
      RECT 49.82 2.275 49.845 2.425 ;
      RECT 49.77 2.283 49.82 2.434 ;
      RECT 49.745 2.288 49.77 2.443 ;
      RECT 49.69 2.294 49.745 2.453 ;
      RECT 49.685 2.299 49.69 2.461 ;
      RECT 49.671 2.302 49.685 2.463 ;
      RECT 49.585 2.314 49.671 2.475 ;
      RECT 49.575 2.326 49.585 2.488 ;
      RECT 49.49 2.339 49.575 2.5 ;
      RECT 49.446 2.356 49.49 2.514 ;
      RECT 49.36 2.373 49.446 2.53 ;
      RECT 49.33 2.387 49.36 2.544 ;
      RECT 49.32 2.392 49.33 2.549 ;
      RECT 49.26 2.395 49.32 2.558 ;
      RECT 52.15 2.665 52.41 2.925 ;
      RECT 52.15 2.665 52.43 2.778 ;
      RECT 52.15 2.665 52.455 2.745 ;
      RECT 52.15 2.665 52.46 2.725 ;
      RECT 52.2 2.44 52.48 2.72 ;
      RECT 51.755 3.175 52.015 3.435 ;
      RECT 51.745 3.032 51.94 3.373 ;
      RECT 51.74 3.14 51.955 3.365 ;
      RECT 51.735 3.19 52.015 3.355 ;
      RECT 51.725 3.267 52.015 3.34 ;
      RECT 51.745 3.115 51.955 3.373 ;
      RECT 51.755 2.99 51.94 3.435 ;
      RECT 51.755 2.885 51.92 3.435 ;
      RECT 51.765 2.872 51.92 3.435 ;
      RECT 51.765 2.83 51.91 3.435 ;
      RECT 51.77 2.755 51.91 3.435 ;
      RECT 51.8 2.405 51.91 3.435 ;
      RECT 51.805 2.135 51.93 2.758 ;
      RECT 51.775 2.71 51.93 2.758 ;
      RECT 51.79 2.512 51.91 3.435 ;
      RECT 51.78 2.622 51.93 2.758 ;
      RECT 51.805 2.135 51.945 2.615 ;
      RECT 51.805 2.135 51.965 2.49 ;
      RECT 51.77 2.135 52.03 2.395 ;
      RECT 51.24 2.44 51.52 2.72 ;
      RECT 51.225 2.44 51.52 2.7 ;
      RECT 49.28 3.305 49.54 3.565 ;
      RECT 51.065 3.16 51.325 3.42 ;
      RECT 51.045 3.18 51.325 3.395 ;
      RECT 51.002 3.18 51.045 3.394 ;
      RECT 50.916 3.181 51.002 3.391 ;
      RECT 50.83 3.182 50.916 3.387 ;
      RECT 50.755 3.184 50.83 3.384 ;
      RECT 50.732 3.185 50.755 3.382 ;
      RECT 50.646 3.186 50.732 3.38 ;
      RECT 50.56 3.187 50.646 3.377 ;
      RECT 50.536 3.188 50.56 3.375 ;
      RECT 50.45 3.19 50.536 3.372 ;
      RECT 50.365 3.192 50.45 3.373 ;
      RECT 50.308 3.193 50.365 3.379 ;
      RECT 50.222 3.195 50.308 3.389 ;
      RECT 50.136 3.198 50.222 3.402 ;
      RECT 50.05 3.2 50.136 3.414 ;
      RECT 50.036 3.201 50.05 3.421 ;
      RECT 49.95 3.202 50.036 3.429 ;
      RECT 49.91 3.204 49.95 3.438 ;
      RECT 49.901 3.205 49.91 3.441 ;
      RECT 49.815 3.213 49.901 3.447 ;
      RECT 49.795 3.222 49.815 3.455 ;
      RECT 49.71 3.237 49.795 3.463 ;
      RECT 49.65 3.26 49.71 3.474 ;
      RECT 49.64 3.272 49.65 3.479 ;
      RECT 49.6 3.282 49.64 3.483 ;
      RECT 49.545 3.299 49.6 3.491 ;
      RECT 49.54 3.309 49.545 3.495 ;
      RECT 50.606 2.44 50.665 2.837 ;
      RECT 50.52 2.44 50.725 2.828 ;
      RECT 50.515 2.47 50.725 2.823 ;
      RECT 50.481 2.47 50.725 2.821 ;
      RECT 50.395 2.47 50.725 2.815 ;
      RECT 50.35 2.47 50.745 2.793 ;
      RECT 50.35 2.47 50.765 2.748 ;
      RECT 50.31 2.47 50.765 2.738 ;
      RECT 50.52 2.44 50.8 2.72 ;
      RECT 50.255 2.44 50.515 2.7 ;
      RECT 49.44 1.92 49.7 2.18 ;
      RECT 49.495 1.88 49.8 2.16 ;
      RECT 49.495 1.855 49.67 2.18 ;
      RECT 43.82 6.28 44.14 6.605 ;
      RECT 43.85 5.695 44.02 6.605 ;
      RECT 43.85 5.695 44.025 6.045 ;
      RECT 43.85 5.695 44.825 5.87 ;
      RECT 44.65 1.965 44.825 5.87 ;
      RECT 40.87 2.84 41.15 3.28 ;
      RECT 40.87 2.84 41.155 3.238 ;
      RECT 40.87 2.84 41.16 3.135 ;
      RECT 40.87 2.84 41.162 3.015 ;
      RECT 40.87 2.84 41.795 3.01 ;
      RECT 41.625 2.025 41.795 3.01 ;
      RECT 40.87 2.805 41.13 3.28 ;
      RECT 44.595 1.965 44.945 2.315 ;
      RECT 43.2 0.915 43.37 2.205 ;
      RECT 41.625 2.025 44.945 2.195 ;
      RECT 31.13 0.885 31.48 1.235 ;
      RECT 31.13 0.915 43.37 1.085 ;
      RECT 44.62 6.655 44.945 6.98 ;
      RECT 43.505 6.745 44.945 6.915 ;
      RECT 43.505 2.395 43.665 6.915 ;
      RECT 43.82 2.365 44.14 2.685 ;
      RECT 43.505 2.395 44.14 2.565 ;
      RECT 42.77 5.855 43.12 6.205 ;
      RECT 42.84 2.705 43.015 6.205 ;
      RECT 42.765 2.705 43.115 3.055 ;
      RECT 32.23 3 32.51 3.28 ;
      RECT 32.2 3 32.51 3.265 ;
      RECT 32.195 2.963 32.455 3.263 ;
      RECT 32.19 2.964 32.455 3.257 ;
      RECT 32.185 2.967 32.455 3.25 ;
      RECT 32.18 3 32.51 3.243 ;
      RECT 32.15 2.97 32.455 3.23 ;
      RECT 32.15 2.997 32.475 3.23 ;
      RECT 32.15 2.987 32.47 3.23 ;
      RECT 32.15 2.972 32.465 3.23 ;
      RECT 32.25 2.962 32.455 3.28 ;
      RECT 32.25 2.957 32.445 3.28 ;
      RECT 32.25 2.955 32.43 3.28 ;
      RECT 32.25 1.42 32.425 3.28 ;
      RECT 42.16 1.34 42.51 1.69 ;
      RECT 32.25 1.42 42.51 1.595 ;
      RECT 37.94 2.455 38.175 2.715 ;
      RECT 41.085 2.235 41.25 2.495 ;
      RECT 40.99 2.225 41.005 2.495 ;
      RECT 39.59 1.795 39.63 1.935 ;
      RECT 41.005 2.23 41.085 2.495 ;
      RECT 40.95 2.225 40.99 2.461 ;
      RECT 40.936 2.225 40.95 2.461 ;
      RECT 40.85 2.23 40.936 2.463 ;
      RECT 40.805 2.237 40.85 2.465 ;
      RECT 40.775 2.237 40.805 2.467 ;
      RECT 40.75 2.232 40.775 2.469 ;
      RECT 40.72 2.228 40.75 2.478 ;
      RECT 40.71 2.225 40.72 2.49 ;
      RECT 40.705 2.225 40.71 2.498 ;
      RECT 40.7 2.225 40.705 2.503 ;
      RECT 40.69 2.224 40.7 2.513 ;
      RECT 40.685 2.223 40.69 2.523 ;
      RECT 40.67 2.222 40.685 2.528 ;
      RECT 40.642 2.219 40.67 2.555 ;
      RECT 40.556 2.211 40.642 2.555 ;
      RECT 40.47 2.2 40.556 2.555 ;
      RECT 40.43 2.185 40.47 2.555 ;
      RECT 40.39 2.159 40.43 2.555 ;
      RECT 40.385 2.141 40.39 2.367 ;
      RECT 40.375 2.137 40.385 2.357 ;
      RECT 40.36 2.127 40.375 2.344 ;
      RECT 40.34 2.111 40.36 2.329 ;
      RECT 40.325 2.096 40.34 2.314 ;
      RECT 40.315 2.085 40.325 2.304 ;
      RECT 40.29 2.069 40.315 2.293 ;
      RECT 40.285 2.056 40.29 2.283 ;
      RECT 40.28 2.052 40.285 2.278 ;
      RECT 40.225 2.038 40.28 2.256 ;
      RECT 40.186 2.019 40.225 2.22 ;
      RECT 40.1 1.993 40.186 2.173 ;
      RECT 40.096 1.975 40.1 2.139 ;
      RECT 40.01 1.956 40.096 2.117 ;
      RECT 40.005 1.938 40.01 2.095 ;
      RECT 40 1.936 40.005 2.093 ;
      RECT 39.99 1.935 40 2.088 ;
      RECT 39.93 1.922 39.99 2.074 ;
      RECT 39.885 1.9 39.93 2.053 ;
      RECT 39.825 1.877 39.885 2.032 ;
      RECT 39.761 1.852 39.825 2.007 ;
      RECT 39.675 1.822 39.761 1.976 ;
      RECT 39.66 1.802 39.675 1.955 ;
      RECT 39.63 1.797 39.66 1.946 ;
      RECT 39.577 1.795 39.59 1.935 ;
      RECT 39.491 1.795 39.577 1.937 ;
      RECT 39.405 1.795 39.491 1.939 ;
      RECT 39.385 1.795 39.405 1.943 ;
      RECT 39.34 1.797 39.385 1.954 ;
      RECT 39.3 1.807 39.34 1.97 ;
      RECT 39.296 1.816 39.3 1.978 ;
      RECT 39.21 1.836 39.296 1.994 ;
      RECT 39.2 1.855 39.21 2.012 ;
      RECT 39.195 1.857 39.2 2.015 ;
      RECT 39.185 1.861 39.195 2.018 ;
      RECT 39.165 1.866 39.185 2.028 ;
      RECT 39.135 1.876 39.165 2.048 ;
      RECT 39.13 1.883 39.135 2.062 ;
      RECT 39.12 1.887 39.13 2.069 ;
      RECT 39.105 1.895 39.12 2.08 ;
      RECT 39.095 1.905 39.105 2.091 ;
      RECT 39.085 1.912 39.095 2.099 ;
      RECT 39.06 1.925 39.085 2.114 ;
      RECT 38.996 1.961 39.06 2.153 ;
      RECT 38.91 2.024 38.996 2.217 ;
      RECT 38.875 2.075 38.91 2.27 ;
      RECT 38.87 2.092 38.875 2.287 ;
      RECT 38.855 2.101 38.87 2.294 ;
      RECT 38.835 2.116 38.855 2.308 ;
      RECT 38.83 2.127 38.835 2.318 ;
      RECT 38.81 2.14 38.83 2.328 ;
      RECT 38.805 2.15 38.81 2.338 ;
      RECT 38.79 2.155 38.805 2.347 ;
      RECT 38.78 2.165 38.79 2.358 ;
      RECT 38.75 2.182 38.78 2.375 ;
      RECT 38.74 2.2 38.75 2.393 ;
      RECT 38.725 2.211 38.74 2.404 ;
      RECT 38.685 2.235 38.725 2.42 ;
      RECT 38.65 2.269 38.685 2.437 ;
      RECT 38.62 2.292 38.65 2.449 ;
      RECT 38.605 2.302 38.62 2.458 ;
      RECT 38.565 2.312 38.605 2.469 ;
      RECT 38.545 2.323 38.565 2.481 ;
      RECT 38.54 2.327 38.545 2.488 ;
      RECT 38.525 2.331 38.54 2.493 ;
      RECT 38.515 2.336 38.525 2.498 ;
      RECT 38.51 2.339 38.515 2.501 ;
      RECT 38.48 2.345 38.51 2.508 ;
      RECT 38.445 2.355 38.48 2.522 ;
      RECT 38.385 2.37 38.445 2.542 ;
      RECT 38.33 2.39 38.385 2.566 ;
      RECT 38.301 2.405 38.33 2.584 ;
      RECT 38.215 2.425 38.301 2.609 ;
      RECT 38.21 2.44 38.215 2.629 ;
      RECT 38.2 2.443 38.21 2.63 ;
      RECT 38.175 2.45 38.2 2.715 ;
      RECT 38.59 3.685 38.6 3.875 ;
      RECT 36.85 3.56 37.13 3.84 ;
      RECT 39.895 2.5 39.9 2.985 ;
      RECT 39.79 2.5 39.85 2.76 ;
      RECT 40.115 3.47 40.12 3.545 ;
      RECT 40.105 3.337 40.115 3.58 ;
      RECT 40.095 3.172 40.105 3.601 ;
      RECT 40.09 3.042 40.095 3.617 ;
      RECT 40.08 2.932 40.09 3.633 ;
      RECT 40.075 2.831 40.08 3.65 ;
      RECT 40.07 2.813 40.075 3.66 ;
      RECT 40.065 2.795 40.07 3.67 ;
      RECT 40.055 2.77 40.065 3.685 ;
      RECT 40.05 2.75 40.055 3.7 ;
      RECT 40.03 2.5 40.05 3.725 ;
      RECT 40.015 2.5 40.03 3.758 ;
      RECT 39.985 2.5 40.015 3.78 ;
      RECT 39.965 2.5 39.985 3.794 ;
      RECT 39.945 2.5 39.965 3.31 ;
      RECT 39.96 3.377 39.965 3.799 ;
      RECT 39.955 3.407 39.96 3.801 ;
      RECT 39.95 3.42 39.955 3.804 ;
      RECT 39.945 3.43 39.95 3.808 ;
      RECT 39.94 2.5 39.945 3.228 ;
      RECT 39.94 3.44 39.945 3.81 ;
      RECT 39.935 2.5 39.94 3.205 ;
      RECT 39.925 3.462 39.94 3.81 ;
      RECT 39.92 2.5 39.935 3.15 ;
      RECT 39.915 3.487 39.925 3.81 ;
      RECT 39.915 2.5 39.92 3.095 ;
      RECT 39.905 2.5 39.915 3.043 ;
      RECT 39.91 3.5 39.915 3.811 ;
      RECT 39.905 3.512 39.91 3.812 ;
      RECT 39.9 2.5 39.905 3.003 ;
      RECT 39.9 3.525 39.905 3.813 ;
      RECT 39.885 3.54 39.9 3.814 ;
      RECT 39.89 2.5 39.895 2.965 ;
      RECT 39.885 2.5 39.89 2.93 ;
      RECT 39.88 2.5 39.885 2.905 ;
      RECT 39.875 3.567 39.885 3.816 ;
      RECT 39.87 2.5 39.88 2.863 ;
      RECT 39.87 3.585 39.875 3.817 ;
      RECT 39.865 2.5 39.87 2.823 ;
      RECT 39.865 3.592 39.87 3.818 ;
      RECT 39.86 2.5 39.865 2.795 ;
      RECT 39.855 3.61 39.865 3.819 ;
      RECT 39.85 2.5 39.86 2.775 ;
      RECT 39.845 3.63 39.855 3.821 ;
      RECT 39.835 3.647 39.845 3.822 ;
      RECT 39.8 3.67 39.835 3.825 ;
      RECT 39.745 3.688 39.8 3.831 ;
      RECT 39.659 3.696 39.745 3.84 ;
      RECT 39.573 3.707 39.659 3.851 ;
      RECT 39.487 3.717 39.573 3.862 ;
      RECT 39.401 3.727 39.487 3.874 ;
      RECT 39.315 3.737 39.401 3.885 ;
      RECT 39.295 3.743 39.315 3.891 ;
      RECT 39.215 3.745 39.295 3.895 ;
      RECT 39.21 3.744 39.215 3.9 ;
      RECT 39.202 3.743 39.21 3.9 ;
      RECT 39.116 3.739 39.202 3.898 ;
      RECT 39.03 3.731 39.116 3.895 ;
      RECT 38.944 3.722 39.03 3.891 ;
      RECT 38.858 3.714 38.944 3.888 ;
      RECT 38.772 3.706 38.858 3.884 ;
      RECT 38.686 3.697 38.772 3.881 ;
      RECT 38.6 3.689 38.686 3.877 ;
      RECT 38.545 3.682 38.59 3.875 ;
      RECT 38.46 3.675 38.545 3.873 ;
      RECT 38.386 3.667 38.46 3.869 ;
      RECT 38.3 3.659 38.386 3.866 ;
      RECT 38.297 3.655 38.3 3.864 ;
      RECT 38.211 3.651 38.297 3.863 ;
      RECT 38.125 3.643 38.211 3.86 ;
      RECT 38.04 3.638 38.125 3.857 ;
      RECT 37.954 3.635 38.04 3.854 ;
      RECT 37.868 3.633 37.954 3.851 ;
      RECT 37.782 3.63 37.868 3.848 ;
      RECT 37.696 3.627 37.782 3.845 ;
      RECT 37.61 3.624 37.696 3.842 ;
      RECT 37.534 3.622 37.61 3.839 ;
      RECT 37.448 3.619 37.534 3.836 ;
      RECT 37.362 3.616 37.448 3.834 ;
      RECT 37.276 3.614 37.362 3.831 ;
      RECT 37.19 3.611 37.276 3.828 ;
      RECT 37.13 3.602 37.19 3.826 ;
      RECT 39.64 3.22 39.715 3.48 ;
      RECT 39.62 3.2 39.625 3.48 ;
      RECT 38.94 2.985 39.045 3.28 ;
      RECT 33.385 2.96 33.455 3.22 ;
      RECT 39.28 2.835 39.285 3.206 ;
      RECT 39.27 2.89 39.275 3.206 ;
      RECT 39.575 2.06 39.635 2.32 ;
      RECT 39.63 3.215 39.64 3.48 ;
      RECT 39.625 3.205 39.63 3.48 ;
      RECT 39.545 3.152 39.62 3.48 ;
      RECT 39.57 2.06 39.575 2.34 ;
      RECT 39.56 2.06 39.57 2.36 ;
      RECT 39.545 2.06 39.56 2.39 ;
      RECT 39.53 2.06 39.545 2.433 ;
      RECT 39.525 3.095 39.545 3.48 ;
      RECT 39.515 2.06 39.53 2.47 ;
      RECT 39.51 3.075 39.525 3.48 ;
      RECT 39.51 2.06 39.515 2.493 ;
      RECT 39.5 2.06 39.51 2.518 ;
      RECT 39.47 3.042 39.51 3.48 ;
      RECT 39.475 2.06 39.5 2.568 ;
      RECT 39.47 2.06 39.475 2.623 ;
      RECT 39.465 2.06 39.47 2.665 ;
      RECT 39.455 3.005 39.47 3.48 ;
      RECT 39.46 2.06 39.465 2.708 ;
      RECT 39.455 2.06 39.46 2.773 ;
      RECT 39.45 2.06 39.455 2.795 ;
      RECT 39.45 2.993 39.455 3.345 ;
      RECT 39.445 2.06 39.45 2.863 ;
      RECT 39.445 2.985 39.45 3.328 ;
      RECT 39.44 2.06 39.445 2.908 ;
      RECT 39.435 2.967 39.445 3.305 ;
      RECT 39.435 2.06 39.44 2.945 ;
      RECT 39.425 2.06 39.435 3.285 ;
      RECT 39.42 2.06 39.425 3.268 ;
      RECT 39.415 2.06 39.42 3.253 ;
      RECT 39.41 2.06 39.415 3.238 ;
      RECT 39.39 2.06 39.41 3.228 ;
      RECT 39.385 2.06 39.39 3.218 ;
      RECT 39.375 2.06 39.385 3.214 ;
      RECT 39.37 2.337 39.375 3.213 ;
      RECT 39.365 2.36 39.37 3.212 ;
      RECT 39.36 2.39 39.365 3.211 ;
      RECT 39.355 2.417 39.36 3.21 ;
      RECT 39.35 2.445 39.355 3.21 ;
      RECT 39.345 2.472 39.35 3.21 ;
      RECT 39.34 2.492 39.345 3.21 ;
      RECT 39.335 2.52 39.34 3.21 ;
      RECT 39.325 2.562 39.335 3.21 ;
      RECT 39.315 2.607 39.325 3.209 ;
      RECT 39.31 2.66 39.315 3.208 ;
      RECT 39.305 2.692 39.31 3.207 ;
      RECT 39.3 2.712 39.305 3.206 ;
      RECT 39.295 2.75 39.3 3.206 ;
      RECT 39.29 2.772 39.295 3.206 ;
      RECT 39.285 2.797 39.29 3.206 ;
      RECT 39.275 2.862 39.28 3.206 ;
      RECT 39.26 2.922 39.27 3.206 ;
      RECT 39.245 2.932 39.26 3.206 ;
      RECT 39.225 2.942 39.245 3.206 ;
      RECT 39.195 2.947 39.225 3.203 ;
      RECT 39.135 2.957 39.195 3.2 ;
      RECT 39.115 2.966 39.135 3.205 ;
      RECT 39.09 2.972 39.115 3.218 ;
      RECT 39.07 2.977 39.09 3.233 ;
      RECT 39.045 2.982 39.07 3.28 ;
      RECT 38.916 2.984 38.94 3.28 ;
      RECT 38.83 2.979 38.916 3.28 ;
      RECT 38.79 2.976 38.83 3.28 ;
      RECT 38.74 2.978 38.79 3.26 ;
      RECT 38.71 2.982 38.74 3.26 ;
      RECT 38.631 2.992 38.71 3.26 ;
      RECT 38.545 3.007 38.631 3.261 ;
      RECT 38.495 3.017 38.545 3.262 ;
      RECT 38.487 3.02 38.495 3.262 ;
      RECT 38.401 3.022 38.487 3.263 ;
      RECT 38.315 3.026 38.401 3.263 ;
      RECT 38.229 3.03 38.315 3.264 ;
      RECT 38.143 3.033 38.229 3.265 ;
      RECT 38.057 3.037 38.143 3.265 ;
      RECT 37.971 3.041 38.057 3.266 ;
      RECT 37.885 3.044 37.971 3.267 ;
      RECT 37.799 3.048 37.885 3.267 ;
      RECT 37.713 3.052 37.799 3.268 ;
      RECT 37.627 3.056 37.713 3.269 ;
      RECT 37.541 3.059 37.627 3.269 ;
      RECT 37.455 3.063 37.541 3.27 ;
      RECT 37.425 3.065 37.455 3.27 ;
      RECT 37.339 3.068 37.425 3.271 ;
      RECT 37.253 3.072 37.339 3.272 ;
      RECT 37.167 3.076 37.253 3.273 ;
      RECT 37.081 3.079 37.167 3.273 ;
      RECT 36.995 3.083 37.081 3.274 ;
      RECT 36.96 3.088 36.995 3.275 ;
      RECT 36.905 3.098 36.96 3.282 ;
      RECT 36.88 3.11 36.905 3.292 ;
      RECT 36.845 3.123 36.88 3.3 ;
      RECT 36.805 3.14 36.845 3.323 ;
      RECT 36.785 3.153 36.805 3.35 ;
      RECT 36.755 3.165 36.785 3.378 ;
      RECT 36.75 3.173 36.755 3.398 ;
      RECT 36.745 3.176 36.75 3.408 ;
      RECT 36.695 3.188 36.745 3.442 ;
      RECT 36.685 3.203 36.695 3.475 ;
      RECT 36.675 3.209 36.685 3.488 ;
      RECT 36.665 3.216 36.675 3.5 ;
      RECT 36.64 3.229 36.665 3.518 ;
      RECT 36.625 3.244 36.64 3.54 ;
      RECT 36.615 3.252 36.625 3.556 ;
      RECT 36.6 3.261 36.615 3.571 ;
      RECT 36.59 3.271 36.6 3.585 ;
      RECT 36.571 3.284 36.59 3.602 ;
      RECT 36.485 3.329 36.571 3.667 ;
      RECT 36.47 3.374 36.485 3.725 ;
      RECT 36.465 3.383 36.47 3.738 ;
      RECT 36.455 3.39 36.465 3.743 ;
      RECT 36.45 3.395 36.455 3.747 ;
      RECT 36.43 3.405 36.45 3.754 ;
      RECT 36.405 3.425 36.43 3.768 ;
      RECT 36.37 3.45 36.405 3.788 ;
      RECT 36.355 3.473 36.37 3.803 ;
      RECT 36.345 3.483 36.355 3.808 ;
      RECT 36.335 3.491 36.345 3.815 ;
      RECT 36.325 3.5 36.335 3.821 ;
      RECT 36.305 3.512 36.325 3.823 ;
      RECT 36.295 3.525 36.305 3.825 ;
      RECT 36.27 3.54 36.295 3.828 ;
      RECT 36.25 3.557 36.27 3.832 ;
      RECT 36.21 3.585 36.25 3.838 ;
      RECT 36.145 3.632 36.21 3.847 ;
      RECT 36.13 3.665 36.145 3.855 ;
      RECT 36.125 3.672 36.13 3.857 ;
      RECT 36.075 3.697 36.125 3.862 ;
      RECT 36.06 3.721 36.075 3.869 ;
      RECT 36.01 3.726 36.06 3.87 ;
      RECT 35.924 3.73 36.01 3.87 ;
      RECT 35.838 3.73 35.924 3.87 ;
      RECT 35.752 3.73 35.838 3.871 ;
      RECT 35.666 3.73 35.752 3.871 ;
      RECT 35.58 3.73 35.666 3.871 ;
      RECT 35.514 3.73 35.58 3.871 ;
      RECT 35.428 3.73 35.514 3.872 ;
      RECT 35.342 3.73 35.428 3.872 ;
      RECT 35.256 3.731 35.342 3.873 ;
      RECT 35.17 3.731 35.256 3.873 ;
      RECT 35.084 3.731 35.17 3.873 ;
      RECT 34.998 3.731 35.084 3.874 ;
      RECT 34.912 3.731 34.998 3.874 ;
      RECT 34.826 3.732 34.912 3.875 ;
      RECT 34.74 3.732 34.826 3.875 ;
      RECT 34.72 3.732 34.74 3.875 ;
      RECT 34.634 3.732 34.72 3.875 ;
      RECT 34.548 3.732 34.634 3.875 ;
      RECT 34.462 3.733 34.548 3.875 ;
      RECT 34.376 3.733 34.462 3.875 ;
      RECT 34.29 3.733 34.376 3.875 ;
      RECT 34.204 3.734 34.29 3.875 ;
      RECT 34.118 3.734 34.204 3.875 ;
      RECT 34.032 3.734 34.118 3.875 ;
      RECT 33.946 3.734 34.032 3.875 ;
      RECT 33.86 3.735 33.946 3.875 ;
      RECT 33.81 3.732 33.86 3.875 ;
      RECT 33.8 3.73 33.81 3.874 ;
      RECT 33.796 3.73 33.8 3.873 ;
      RECT 33.71 3.725 33.796 3.868 ;
      RECT 33.688 3.718 33.71 3.862 ;
      RECT 33.602 3.709 33.688 3.856 ;
      RECT 33.516 3.696 33.602 3.847 ;
      RECT 33.43 3.682 33.516 3.837 ;
      RECT 33.385 3.672 33.43 3.83 ;
      RECT 33.365 2.96 33.385 3.238 ;
      RECT 33.365 3.665 33.385 3.826 ;
      RECT 33.335 2.96 33.365 3.26 ;
      RECT 33.325 3.632 33.365 3.823 ;
      RECT 33.32 2.96 33.335 3.28 ;
      RECT 33.32 3.597 33.325 3.821 ;
      RECT 33.315 2.96 33.32 3.405 ;
      RECT 33.315 3.557 33.32 3.821 ;
      RECT 33.305 2.96 33.315 3.821 ;
      RECT 33.23 2.96 33.305 3.815 ;
      RECT 33.2 2.96 33.23 3.805 ;
      RECT 33.195 2.96 33.2 3.797 ;
      RECT 33.19 3.002 33.195 3.79 ;
      RECT 33.18 3.071 33.19 3.781 ;
      RECT 33.175 3.141 33.18 3.733 ;
      RECT 33.17 3.205 33.175 3.63 ;
      RECT 33.165 3.24 33.17 3.585 ;
      RECT 33.163 3.277 33.165 3.477 ;
      RECT 33.16 3.285 33.163 3.47 ;
      RECT 33.155 3.35 33.16 3.413 ;
      RECT 37.23 2.44 37.51 2.72 ;
      RECT 37.22 2.44 37.51 2.583 ;
      RECT 37.175 2.305 37.435 2.565 ;
      RECT 37.175 2.42 37.49 2.565 ;
      RECT 37.175 2.39 37.485 2.565 ;
      RECT 37.175 2.377 37.475 2.565 ;
      RECT 37.175 2.367 37.47 2.565 ;
      RECT 33.15 2.35 33.41 2.61 ;
      RECT 36.92 1.9 37.18 2.16 ;
      RECT 36.91 1.925 37.18 2.12 ;
      RECT 36.905 1.925 36.91 2.119 ;
      RECT 36.835 1.92 36.905 2.111 ;
      RECT 36.75 1.907 36.835 2.094 ;
      RECT 36.746 1.899 36.75 2.084 ;
      RECT 36.66 1.892 36.746 2.074 ;
      RECT 36.651 1.884 36.66 2.064 ;
      RECT 36.565 1.877 36.651 2.052 ;
      RECT 36.545 1.868 36.565 2.038 ;
      RECT 36.49 1.863 36.545 2.03 ;
      RECT 36.48 1.857 36.49 2.024 ;
      RECT 36.46 1.855 36.48 2.02 ;
      RECT 36.452 1.854 36.46 2.016 ;
      RECT 36.366 1.846 36.452 2.005 ;
      RECT 36.28 1.832 36.366 1.985 ;
      RECT 36.22 1.82 36.28 1.97 ;
      RECT 36.21 1.815 36.22 1.965 ;
      RECT 36.16 1.815 36.21 1.967 ;
      RECT 36.113 1.817 36.16 1.971 ;
      RECT 36.027 1.824 36.113 1.976 ;
      RECT 35.941 1.832 36.027 1.982 ;
      RECT 35.855 1.841 35.941 1.988 ;
      RECT 35.796 1.847 35.855 1.993 ;
      RECT 35.71 1.852 35.796 1.999 ;
      RECT 35.635 1.857 35.71 2.005 ;
      RECT 35.596 1.859 35.635 2.01 ;
      RECT 35.51 1.856 35.596 2.015 ;
      RECT 35.425 1.854 35.51 2.022 ;
      RECT 35.393 1.853 35.425 2.025 ;
      RECT 35.307 1.852 35.393 2.026 ;
      RECT 35.221 1.851 35.307 2.027 ;
      RECT 35.135 1.85 35.221 2.027 ;
      RECT 35.049 1.849 35.135 2.028 ;
      RECT 34.963 1.848 35.049 2.029 ;
      RECT 34.877 1.847 34.963 2.03 ;
      RECT 34.791 1.846 34.877 2.03 ;
      RECT 34.705 1.845 34.791 2.031 ;
      RECT 34.655 1.845 34.705 2.032 ;
      RECT 34.641 1.846 34.655 2.032 ;
      RECT 34.555 1.853 34.641 2.033 ;
      RECT 34.481 1.864 34.555 2.034 ;
      RECT 34.395 1.873 34.481 2.035 ;
      RECT 34.36 1.88 34.395 2.05 ;
      RECT 34.335 1.883 34.36 2.08 ;
      RECT 34.31 1.892 34.335 2.109 ;
      RECT 34.3 1.903 34.31 2.129 ;
      RECT 34.29 1.911 34.3 2.143 ;
      RECT 34.285 1.917 34.29 2.153 ;
      RECT 34.26 1.934 34.285 2.17 ;
      RECT 34.245 1.956 34.26 2.198 ;
      RECT 34.215 1.982 34.245 2.228 ;
      RECT 34.195 2.011 34.215 2.258 ;
      RECT 34.19 2.026 34.195 2.275 ;
      RECT 34.17 2.041 34.19 2.29 ;
      RECT 34.16 2.059 34.17 2.308 ;
      RECT 34.15 2.07 34.16 2.323 ;
      RECT 34.1 2.102 34.15 2.349 ;
      RECT 34.095 2.132 34.1 2.369 ;
      RECT 34.085 2.145 34.095 2.375 ;
      RECT 34.076 2.155 34.085 2.383 ;
      RECT 34.065 2.166 34.076 2.391 ;
      RECT 34.06 2.176 34.065 2.397 ;
      RECT 34.045 2.197 34.06 2.404 ;
      RECT 34.03 2.227 34.045 2.412 ;
      RECT 33.995 2.257 34.03 2.418 ;
      RECT 33.97 2.275 33.995 2.425 ;
      RECT 33.92 2.283 33.97 2.434 ;
      RECT 33.895 2.288 33.92 2.443 ;
      RECT 33.84 2.294 33.895 2.453 ;
      RECT 33.835 2.299 33.84 2.461 ;
      RECT 33.821 2.302 33.835 2.463 ;
      RECT 33.735 2.314 33.821 2.475 ;
      RECT 33.725 2.326 33.735 2.488 ;
      RECT 33.64 2.339 33.725 2.5 ;
      RECT 33.596 2.356 33.64 2.514 ;
      RECT 33.51 2.373 33.596 2.53 ;
      RECT 33.48 2.387 33.51 2.544 ;
      RECT 33.47 2.392 33.48 2.549 ;
      RECT 33.41 2.395 33.47 2.558 ;
      RECT 36.3 2.665 36.56 2.925 ;
      RECT 36.3 2.665 36.58 2.778 ;
      RECT 36.3 2.665 36.605 2.745 ;
      RECT 36.3 2.665 36.61 2.725 ;
      RECT 36.35 2.44 36.63 2.72 ;
      RECT 35.905 3.175 36.165 3.435 ;
      RECT 35.895 3.032 36.09 3.373 ;
      RECT 35.89 3.14 36.105 3.365 ;
      RECT 35.885 3.19 36.165 3.355 ;
      RECT 35.875 3.267 36.165 3.34 ;
      RECT 35.895 3.115 36.105 3.373 ;
      RECT 35.905 2.99 36.09 3.435 ;
      RECT 35.905 2.885 36.07 3.435 ;
      RECT 35.915 2.872 36.07 3.435 ;
      RECT 35.915 2.83 36.06 3.435 ;
      RECT 35.92 2.755 36.06 3.435 ;
      RECT 35.95 2.405 36.06 3.435 ;
      RECT 35.955 2.135 36.08 2.758 ;
      RECT 35.925 2.71 36.08 2.758 ;
      RECT 35.94 2.512 36.06 3.435 ;
      RECT 35.93 2.622 36.08 2.758 ;
      RECT 35.955 2.135 36.095 2.615 ;
      RECT 35.955 2.135 36.115 2.49 ;
      RECT 35.92 2.135 36.18 2.395 ;
      RECT 35.39 2.44 35.67 2.72 ;
      RECT 35.375 2.44 35.67 2.7 ;
      RECT 33.43 3.305 33.69 3.565 ;
      RECT 35.215 3.16 35.475 3.42 ;
      RECT 35.195 3.18 35.475 3.395 ;
      RECT 35.152 3.18 35.195 3.394 ;
      RECT 35.066 3.181 35.152 3.391 ;
      RECT 34.98 3.182 35.066 3.387 ;
      RECT 34.905 3.184 34.98 3.384 ;
      RECT 34.882 3.185 34.905 3.382 ;
      RECT 34.796 3.186 34.882 3.38 ;
      RECT 34.71 3.187 34.796 3.377 ;
      RECT 34.686 3.188 34.71 3.375 ;
      RECT 34.6 3.19 34.686 3.372 ;
      RECT 34.515 3.192 34.6 3.373 ;
      RECT 34.458 3.193 34.515 3.379 ;
      RECT 34.372 3.195 34.458 3.389 ;
      RECT 34.286 3.198 34.372 3.402 ;
      RECT 34.2 3.2 34.286 3.414 ;
      RECT 34.186 3.201 34.2 3.421 ;
      RECT 34.1 3.202 34.186 3.429 ;
      RECT 34.06 3.204 34.1 3.438 ;
      RECT 34.051 3.205 34.06 3.441 ;
      RECT 33.965 3.213 34.051 3.447 ;
      RECT 33.945 3.222 33.965 3.455 ;
      RECT 33.86 3.237 33.945 3.463 ;
      RECT 33.8 3.26 33.86 3.474 ;
      RECT 33.79 3.272 33.8 3.479 ;
      RECT 33.75 3.282 33.79 3.483 ;
      RECT 33.695 3.299 33.75 3.491 ;
      RECT 33.69 3.309 33.695 3.495 ;
      RECT 34.756 2.44 34.815 2.837 ;
      RECT 34.67 2.44 34.875 2.828 ;
      RECT 34.665 2.47 34.875 2.823 ;
      RECT 34.631 2.47 34.875 2.821 ;
      RECT 34.545 2.47 34.875 2.815 ;
      RECT 34.5 2.47 34.895 2.793 ;
      RECT 34.5 2.47 34.915 2.748 ;
      RECT 34.46 2.47 34.915 2.738 ;
      RECT 34.67 2.44 34.95 2.72 ;
      RECT 34.405 2.44 34.665 2.7 ;
      RECT 33.59 1.92 33.85 2.18 ;
      RECT 33.645 1.88 33.95 2.16 ;
      RECT 33.645 1.855 33.82 2.18 ;
      RECT 27.97 6.28 28.29 6.605 ;
      RECT 28 5.695 28.17 6.605 ;
      RECT 28 5.695 28.175 6.045 ;
      RECT 28 5.695 28.975 5.87 ;
      RECT 28.8 1.965 28.975 5.87 ;
      RECT 25.02 2.84 25.3 3.28 ;
      RECT 25.02 2.84 25.305 3.238 ;
      RECT 25.02 2.84 25.31 3.135 ;
      RECT 25.02 2.84 25.312 3.015 ;
      RECT 25.02 2.84 25.945 3.01 ;
      RECT 25.775 2.025 25.945 3.01 ;
      RECT 25.02 2.805 25.28 3.28 ;
      RECT 28.745 1.965 29.095 2.315 ;
      RECT 27.18 0.915 27.35 2.21 ;
      RECT 25.775 2.025 29.095 2.195 ;
      RECT 15.28 0.885 15.63 1.235 ;
      RECT 15.28 0.915 27.35 1.085 ;
      RECT 28.77 6.655 29.095 6.98 ;
      RECT 27.655 6.745 29.095 6.915 ;
      RECT 27.655 2.395 27.815 6.915 ;
      RECT 27.97 2.365 28.29 2.685 ;
      RECT 27.655 2.395 28.29 2.565 ;
      RECT 26.92 5.855 27.27 6.205 ;
      RECT 26.99 2.705 27.165 6.205 ;
      RECT 26.915 2.705 27.265 3.055 ;
      RECT 16.38 3 16.66 3.28 ;
      RECT 16.35 3 16.66 3.265 ;
      RECT 16.345 2.963 16.605 3.263 ;
      RECT 16.34 2.964 16.605 3.257 ;
      RECT 16.335 2.967 16.605 3.25 ;
      RECT 16.33 3 16.66 3.243 ;
      RECT 16.3 2.97 16.605 3.23 ;
      RECT 16.3 2.997 16.625 3.23 ;
      RECT 16.3 2.987 16.62 3.23 ;
      RECT 16.3 2.972 16.615 3.23 ;
      RECT 16.4 2.962 16.605 3.28 ;
      RECT 16.4 2.957 16.595 3.28 ;
      RECT 16.4 2.955 16.58 3.28 ;
      RECT 16.4 1.42 16.575 3.28 ;
      RECT 26.31 1.34 26.66 1.69 ;
      RECT 16.4 1.42 26.66 1.595 ;
      RECT 22.09 2.455 22.325 2.715 ;
      RECT 25.235 2.235 25.4 2.495 ;
      RECT 25.14 2.225 25.155 2.495 ;
      RECT 23.74 1.795 23.78 1.935 ;
      RECT 25.155 2.23 25.235 2.495 ;
      RECT 25.1 2.225 25.14 2.461 ;
      RECT 25.086 2.225 25.1 2.461 ;
      RECT 25 2.23 25.086 2.463 ;
      RECT 24.955 2.237 25 2.465 ;
      RECT 24.925 2.237 24.955 2.467 ;
      RECT 24.9 2.232 24.925 2.469 ;
      RECT 24.87 2.228 24.9 2.478 ;
      RECT 24.86 2.225 24.87 2.49 ;
      RECT 24.855 2.225 24.86 2.498 ;
      RECT 24.85 2.225 24.855 2.503 ;
      RECT 24.84 2.224 24.85 2.513 ;
      RECT 24.835 2.223 24.84 2.523 ;
      RECT 24.82 2.222 24.835 2.528 ;
      RECT 24.792 2.219 24.82 2.555 ;
      RECT 24.706 2.211 24.792 2.555 ;
      RECT 24.62 2.2 24.706 2.555 ;
      RECT 24.58 2.185 24.62 2.555 ;
      RECT 24.54 2.159 24.58 2.555 ;
      RECT 24.535 2.141 24.54 2.367 ;
      RECT 24.525 2.137 24.535 2.357 ;
      RECT 24.51 2.127 24.525 2.344 ;
      RECT 24.49 2.111 24.51 2.329 ;
      RECT 24.475 2.096 24.49 2.314 ;
      RECT 24.465 2.085 24.475 2.304 ;
      RECT 24.44 2.069 24.465 2.293 ;
      RECT 24.435 2.056 24.44 2.283 ;
      RECT 24.43 2.052 24.435 2.278 ;
      RECT 24.375 2.038 24.43 2.256 ;
      RECT 24.336 2.019 24.375 2.22 ;
      RECT 24.25 1.993 24.336 2.173 ;
      RECT 24.246 1.975 24.25 2.139 ;
      RECT 24.16 1.956 24.246 2.117 ;
      RECT 24.155 1.938 24.16 2.095 ;
      RECT 24.15 1.936 24.155 2.093 ;
      RECT 24.14 1.935 24.15 2.088 ;
      RECT 24.08 1.922 24.14 2.074 ;
      RECT 24.035 1.9 24.08 2.053 ;
      RECT 23.975 1.877 24.035 2.032 ;
      RECT 23.911 1.852 23.975 2.007 ;
      RECT 23.825 1.822 23.911 1.976 ;
      RECT 23.81 1.802 23.825 1.955 ;
      RECT 23.78 1.797 23.81 1.946 ;
      RECT 23.727 1.795 23.74 1.935 ;
      RECT 23.641 1.795 23.727 1.937 ;
      RECT 23.555 1.795 23.641 1.939 ;
      RECT 23.535 1.795 23.555 1.943 ;
      RECT 23.49 1.797 23.535 1.954 ;
      RECT 23.45 1.807 23.49 1.97 ;
      RECT 23.446 1.816 23.45 1.978 ;
      RECT 23.36 1.836 23.446 1.994 ;
      RECT 23.35 1.855 23.36 2.012 ;
      RECT 23.345 1.857 23.35 2.015 ;
      RECT 23.335 1.861 23.345 2.018 ;
      RECT 23.315 1.866 23.335 2.028 ;
      RECT 23.285 1.876 23.315 2.048 ;
      RECT 23.28 1.883 23.285 2.062 ;
      RECT 23.27 1.887 23.28 2.069 ;
      RECT 23.255 1.895 23.27 2.08 ;
      RECT 23.245 1.905 23.255 2.091 ;
      RECT 23.235 1.912 23.245 2.099 ;
      RECT 23.21 1.925 23.235 2.114 ;
      RECT 23.146 1.961 23.21 2.153 ;
      RECT 23.06 2.024 23.146 2.217 ;
      RECT 23.025 2.075 23.06 2.27 ;
      RECT 23.02 2.092 23.025 2.287 ;
      RECT 23.005 2.101 23.02 2.294 ;
      RECT 22.985 2.116 23.005 2.308 ;
      RECT 22.98 2.127 22.985 2.318 ;
      RECT 22.96 2.14 22.98 2.328 ;
      RECT 22.955 2.15 22.96 2.338 ;
      RECT 22.94 2.155 22.955 2.347 ;
      RECT 22.93 2.165 22.94 2.358 ;
      RECT 22.9 2.182 22.93 2.375 ;
      RECT 22.89 2.2 22.9 2.393 ;
      RECT 22.875 2.211 22.89 2.404 ;
      RECT 22.835 2.235 22.875 2.42 ;
      RECT 22.8 2.269 22.835 2.437 ;
      RECT 22.77 2.292 22.8 2.449 ;
      RECT 22.755 2.302 22.77 2.458 ;
      RECT 22.715 2.312 22.755 2.469 ;
      RECT 22.695 2.323 22.715 2.481 ;
      RECT 22.69 2.327 22.695 2.488 ;
      RECT 22.675 2.331 22.69 2.493 ;
      RECT 22.665 2.336 22.675 2.498 ;
      RECT 22.66 2.339 22.665 2.501 ;
      RECT 22.63 2.345 22.66 2.508 ;
      RECT 22.595 2.355 22.63 2.522 ;
      RECT 22.535 2.37 22.595 2.542 ;
      RECT 22.48 2.39 22.535 2.566 ;
      RECT 22.451 2.405 22.48 2.584 ;
      RECT 22.365 2.425 22.451 2.609 ;
      RECT 22.36 2.44 22.365 2.629 ;
      RECT 22.35 2.443 22.36 2.63 ;
      RECT 22.325 2.45 22.35 2.715 ;
      RECT 22.74 3.685 22.75 3.875 ;
      RECT 21 3.56 21.28 3.84 ;
      RECT 24.045 2.5 24.05 2.985 ;
      RECT 23.94 2.5 24 2.76 ;
      RECT 24.265 3.47 24.27 3.545 ;
      RECT 24.255 3.337 24.265 3.58 ;
      RECT 24.245 3.172 24.255 3.601 ;
      RECT 24.24 3.042 24.245 3.617 ;
      RECT 24.23 2.932 24.24 3.633 ;
      RECT 24.225 2.831 24.23 3.65 ;
      RECT 24.22 2.813 24.225 3.66 ;
      RECT 24.215 2.795 24.22 3.67 ;
      RECT 24.205 2.77 24.215 3.685 ;
      RECT 24.2 2.75 24.205 3.7 ;
      RECT 24.18 2.5 24.2 3.725 ;
      RECT 24.165 2.5 24.18 3.758 ;
      RECT 24.135 2.5 24.165 3.78 ;
      RECT 24.115 2.5 24.135 3.794 ;
      RECT 24.095 2.5 24.115 3.31 ;
      RECT 24.11 3.377 24.115 3.799 ;
      RECT 24.105 3.407 24.11 3.801 ;
      RECT 24.1 3.42 24.105 3.804 ;
      RECT 24.095 3.43 24.1 3.808 ;
      RECT 24.09 2.5 24.095 3.228 ;
      RECT 24.09 3.44 24.095 3.81 ;
      RECT 24.085 2.5 24.09 3.205 ;
      RECT 24.075 3.462 24.09 3.81 ;
      RECT 24.07 2.5 24.085 3.15 ;
      RECT 24.065 3.487 24.075 3.81 ;
      RECT 24.065 2.5 24.07 3.095 ;
      RECT 24.055 2.5 24.065 3.043 ;
      RECT 24.06 3.5 24.065 3.811 ;
      RECT 24.055 3.512 24.06 3.812 ;
      RECT 24.05 2.5 24.055 3.003 ;
      RECT 24.05 3.525 24.055 3.813 ;
      RECT 24.035 3.54 24.05 3.814 ;
      RECT 24.04 2.5 24.045 2.965 ;
      RECT 24.035 2.5 24.04 2.93 ;
      RECT 24.03 2.5 24.035 2.905 ;
      RECT 24.025 3.567 24.035 3.816 ;
      RECT 24.02 2.5 24.03 2.863 ;
      RECT 24.02 3.585 24.025 3.817 ;
      RECT 24.015 2.5 24.02 2.823 ;
      RECT 24.015 3.592 24.02 3.818 ;
      RECT 24.01 2.5 24.015 2.795 ;
      RECT 24.005 3.61 24.015 3.819 ;
      RECT 24 2.5 24.01 2.775 ;
      RECT 23.995 3.63 24.005 3.821 ;
      RECT 23.985 3.647 23.995 3.822 ;
      RECT 23.95 3.67 23.985 3.825 ;
      RECT 23.895 3.688 23.95 3.831 ;
      RECT 23.809 3.696 23.895 3.84 ;
      RECT 23.723 3.707 23.809 3.851 ;
      RECT 23.637 3.717 23.723 3.862 ;
      RECT 23.551 3.727 23.637 3.874 ;
      RECT 23.465 3.737 23.551 3.885 ;
      RECT 23.445 3.743 23.465 3.891 ;
      RECT 23.365 3.745 23.445 3.895 ;
      RECT 23.36 3.744 23.365 3.9 ;
      RECT 23.352 3.743 23.36 3.9 ;
      RECT 23.266 3.739 23.352 3.898 ;
      RECT 23.18 3.731 23.266 3.895 ;
      RECT 23.094 3.722 23.18 3.891 ;
      RECT 23.008 3.714 23.094 3.888 ;
      RECT 22.922 3.706 23.008 3.884 ;
      RECT 22.836 3.697 22.922 3.881 ;
      RECT 22.75 3.689 22.836 3.877 ;
      RECT 22.695 3.682 22.74 3.875 ;
      RECT 22.61 3.675 22.695 3.873 ;
      RECT 22.536 3.667 22.61 3.869 ;
      RECT 22.45 3.659 22.536 3.866 ;
      RECT 22.447 3.655 22.45 3.864 ;
      RECT 22.361 3.651 22.447 3.863 ;
      RECT 22.275 3.643 22.361 3.86 ;
      RECT 22.19 3.638 22.275 3.857 ;
      RECT 22.104 3.635 22.19 3.854 ;
      RECT 22.018 3.633 22.104 3.851 ;
      RECT 21.932 3.63 22.018 3.848 ;
      RECT 21.846 3.627 21.932 3.845 ;
      RECT 21.76 3.624 21.846 3.842 ;
      RECT 21.684 3.622 21.76 3.839 ;
      RECT 21.598 3.619 21.684 3.836 ;
      RECT 21.512 3.616 21.598 3.834 ;
      RECT 21.426 3.614 21.512 3.831 ;
      RECT 21.34 3.611 21.426 3.828 ;
      RECT 21.28 3.602 21.34 3.826 ;
      RECT 23.79 3.22 23.865 3.48 ;
      RECT 23.77 3.2 23.775 3.48 ;
      RECT 23.09 2.985 23.195 3.28 ;
      RECT 17.535 2.96 17.605 3.22 ;
      RECT 23.43 2.835 23.435 3.206 ;
      RECT 23.42 2.89 23.425 3.206 ;
      RECT 23.725 2.06 23.785 2.32 ;
      RECT 23.78 3.215 23.79 3.48 ;
      RECT 23.775 3.205 23.78 3.48 ;
      RECT 23.695 3.152 23.77 3.48 ;
      RECT 23.72 2.06 23.725 2.34 ;
      RECT 23.71 2.06 23.72 2.36 ;
      RECT 23.695 2.06 23.71 2.39 ;
      RECT 23.68 2.06 23.695 2.433 ;
      RECT 23.675 3.095 23.695 3.48 ;
      RECT 23.665 2.06 23.68 2.47 ;
      RECT 23.66 3.075 23.675 3.48 ;
      RECT 23.66 2.06 23.665 2.493 ;
      RECT 23.65 2.06 23.66 2.518 ;
      RECT 23.62 3.042 23.66 3.48 ;
      RECT 23.625 2.06 23.65 2.568 ;
      RECT 23.62 2.06 23.625 2.623 ;
      RECT 23.615 2.06 23.62 2.665 ;
      RECT 23.605 3.005 23.62 3.48 ;
      RECT 23.61 2.06 23.615 2.708 ;
      RECT 23.605 2.06 23.61 2.773 ;
      RECT 23.6 2.06 23.605 2.795 ;
      RECT 23.6 2.993 23.605 3.345 ;
      RECT 23.595 2.06 23.6 2.863 ;
      RECT 23.595 2.985 23.6 3.328 ;
      RECT 23.59 2.06 23.595 2.908 ;
      RECT 23.585 2.967 23.595 3.305 ;
      RECT 23.585 2.06 23.59 2.945 ;
      RECT 23.575 2.06 23.585 3.285 ;
      RECT 23.57 2.06 23.575 3.268 ;
      RECT 23.565 2.06 23.57 3.253 ;
      RECT 23.56 2.06 23.565 3.238 ;
      RECT 23.54 2.06 23.56 3.228 ;
      RECT 23.535 2.06 23.54 3.218 ;
      RECT 23.525 2.06 23.535 3.214 ;
      RECT 23.52 2.337 23.525 3.213 ;
      RECT 23.515 2.36 23.52 3.212 ;
      RECT 23.51 2.39 23.515 3.211 ;
      RECT 23.505 2.417 23.51 3.21 ;
      RECT 23.5 2.445 23.505 3.21 ;
      RECT 23.495 2.472 23.5 3.21 ;
      RECT 23.49 2.492 23.495 3.21 ;
      RECT 23.485 2.52 23.49 3.21 ;
      RECT 23.475 2.562 23.485 3.21 ;
      RECT 23.465 2.607 23.475 3.209 ;
      RECT 23.46 2.66 23.465 3.208 ;
      RECT 23.455 2.692 23.46 3.207 ;
      RECT 23.45 2.712 23.455 3.206 ;
      RECT 23.445 2.75 23.45 3.206 ;
      RECT 23.44 2.772 23.445 3.206 ;
      RECT 23.435 2.797 23.44 3.206 ;
      RECT 23.425 2.862 23.43 3.206 ;
      RECT 23.41 2.922 23.42 3.206 ;
      RECT 23.395 2.932 23.41 3.206 ;
      RECT 23.375 2.942 23.395 3.206 ;
      RECT 23.345 2.947 23.375 3.203 ;
      RECT 23.285 2.957 23.345 3.2 ;
      RECT 23.265 2.966 23.285 3.205 ;
      RECT 23.24 2.972 23.265 3.218 ;
      RECT 23.22 2.977 23.24 3.233 ;
      RECT 23.195 2.982 23.22 3.28 ;
      RECT 23.066 2.984 23.09 3.28 ;
      RECT 22.98 2.979 23.066 3.28 ;
      RECT 22.94 2.976 22.98 3.28 ;
      RECT 22.89 2.978 22.94 3.26 ;
      RECT 22.86 2.982 22.89 3.26 ;
      RECT 22.781 2.992 22.86 3.26 ;
      RECT 22.695 3.007 22.781 3.261 ;
      RECT 22.645 3.017 22.695 3.262 ;
      RECT 22.637 3.02 22.645 3.262 ;
      RECT 22.551 3.022 22.637 3.263 ;
      RECT 22.465 3.026 22.551 3.263 ;
      RECT 22.379 3.03 22.465 3.264 ;
      RECT 22.293 3.033 22.379 3.265 ;
      RECT 22.207 3.037 22.293 3.265 ;
      RECT 22.121 3.041 22.207 3.266 ;
      RECT 22.035 3.044 22.121 3.267 ;
      RECT 21.949 3.048 22.035 3.267 ;
      RECT 21.863 3.052 21.949 3.268 ;
      RECT 21.777 3.056 21.863 3.269 ;
      RECT 21.691 3.059 21.777 3.269 ;
      RECT 21.605 3.063 21.691 3.27 ;
      RECT 21.575 3.065 21.605 3.27 ;
      RECT 21.489 3.068 21.575 3.271 ;
      RECT 21.403 3.072 21.489 3.272 ;
      RECT 21.317 3.076 21.403 3.273 ;
      RECT 21.231 3.079 21.317 3.273 ;
      RECT 21.145 3.083 21.231 3.274 ;
      RECT 21.11 3.088 21.145 3.275 ;
      RECT 21.055 3.098 21.11 3.282 ;
      RECT 21.03 3.11 21.055 3.292 ;
      RECT 20.995 3.123 21.03 3.3 ;
      RECT 20.955 3.14 20.995 3.323 ;
      RECT 20.935 3.153 20.955 3.35 ;
      RECT 20.905 3.165 20.935 3.378 ;
      RECT 20.9 3.173 20.905 3.398 ;
      RECT 20.895 3.176 20.9 3.408 ;
      RECT 20.845 3.188 20.895 3.442 ;
      RECT 20.835 3.203 20.845 3.475 ;
      RECT 20.825 3.209 20.835 3.488 ;
      RECT 20.815 3.216 20.825 3.5 ;
      RECT 20.79 3.229 20.815 3.518 ;
      RECT 20.775 3.244 20.79 3.54 ;
      RECT 20.765 3.252 20.775 3.556 ;
      RECT 20.75 3.261 20.765 3.571 ;
      RECT 20.74 3.271 20.75 3.585 ;
      RECT 20.721 3.284 20.74 3.602 ;
      RECT 20.635 3.329 20.721 3.667 ;
      RECT 20.62 3.374 20.635 3.725 ;
      RECT 20.615 3.383 20.62 3.738 ;
      RECT 20.605 3.39 20.615 3.743 ;
      RECT 20.6 3.395 20.605 3.747 ;
      RECT 20.58 3.405 20.6 3.754 ;
      RECT 20.555 3.425 20.58 3.768 ;
      RECT 20.52 3.45 20.555 3.788 ;
      RECT 20.505 3.473 20.52 3.803 ;
      RECT 20.495 3.483 20.505 3.808 ;
      RECT 20.485 3.491 20.495 3.815 ;
      RECT 20.475 3.5 20.485 3.821 ;
      RECT 20.455 3.512 20.475 3.823 ;
      RECT 20.445 3.525 20.455 3.825 ;
      RECT 20.42 3.54 20.445 3.828 ;
      RECT 20.4 3.557 20.42 3.832 ;
      RECT 20.36 3.585 20.4 3.838 ;
      RECT 20.295 3.632 20.36 3.847 ;
      RECT 20.28 3.665 20.295 3.855 ;
      RECT 20.275 3.672 20.28 3.857 ;
      RECT 20.225 3.697 20.275 3.862 ;
      RECT 20.21 3.721 20.225 3.869 ;
      RECT 20.16 3.726 20.21 3.87 ;
      RECT 20.074 3.73 20.16 3.87 ;
      RECT 19.988 3.73 20.074 3.87 ;
      RECT 19.902 3.73 19.988 3.871 ;
      RECT 19.816 3.73 19.902 3.871 ;
      RECT 19.73 3.73 19.816 3.871 ;
      RECT 19.664 3.73 19.73 3.871 ;
      RECT 19.578 3.73 19.664 3.872 ;
      RECT 19.492 3.73 19.578 3.872 ;
      RECT 19.406 3.731 19.492 3.873 ;
      RECT 19.32 3.731 19.406 3.873 ;
      RECT 19.234 3.731 19.32 3.873 ;
      RECT 19.148 3.731 19.234 3.874 ;
      RECT 19.062 3.731 19.148 3.874 ;
      RECT 18.976 3.732 19.062 3.875 ;
      RECT 18.89 3.732 18.976 3.875 ;
      RECT 18.87 3.732 18.89 3.875 ;
      RECT 18.784 3.732 18.87 3.875 ;
      RECT 18.698 3.732 18.784 3.875 ;
      RECT 18.612 3.733 18.698 3.875 ;
      RECT 18.526 3.733 18.612 3.875 ;
      RECT 18.44 3.733 18.526 3.875 ;
      RECT 18.354 3.734 18.44 3.875 ;
      RECT 18.268 3.734 18.354 3.875 ;
      RECT 18.182 3.734 18.268 3.875 ;
      RECT 18.096 3.734 18.182 3.875 ;
      RECT 18.01 3.735 18.096 3.875 ;
      RECT 17.96 3.732 18.01 3.875 ;
      RECT 17.95 3.73 17.96 3.874 ;
      RECT 17.946 3.73 17.95 3.873 ;
      RECT 17.86 3.725 17.946 3.868 ;
      RECT 17.838 3.718 17.86 3.862 ;
      RECT 17.752 3.709 17.838 3.856 ;
      RECT 17.666 3.696 17.752 3.847 ;
      RECT 17.58 3.682 17.666 3.837 ;
      RECT 17.535 3.672 17.58 3.83 ;
      RECT 17.515 2.96 17.535 3.238 ;
      RECT 17.515 3.665 17.535 3.826 ;
      RECT 17.485 2.96 17.515 3.26 ;
      RECT 17.475 3.632 17.515 3.823 ;
      RECT 17.47 2.96 17.485 3.28 ;
      RECT 17.47 3.597 17.475 3.821 ;
      RECT 17.465 2.96 17.47 3.405 ;
      RECT 17.465 3.557 17.47 3.821 ;
      RECT 17.455 2.96 17.465 3.821 ;
      RECT 17.38 2.96 17.455 3.815 ;
      RECT 17.35 2.96 17.38 3.805 ;
      RECT 17.345 2.96 17.35 3.797 ;
      RECT 17.34 3.002 17.345 3.79 ;
      RECT 17.33 3.071 17.34 3.781 ;
      RECT 17.325 3.141 17.33 3.733 ;
      RECT 17.32 3.205 17.325 3.63 ;
      RECT 17.315 3.24 17.32 3.585 ;
      RECT 17.313 3.277 17.315 3.477 ;
      RECT 17.31 3.285 17.313 3.47 ;
      RECT 17.305 3.35 17.31 3.413 ;
      RECT 21.38 2.44 21.66 2.72 ;
      RECT 21.37 2.44 21.66 2.583 ;
      RECT 21.325 2.305 21.585 2.565 ;
      RECT 21.325 2.42 21.64 2.565 ;
      RECT 21.325 2.39 21.635 2.565 ;
      RECT 21.325 2.377 21.625 2.565 ;
      RECT 21.325 2.367 21.62 2.565 ;
      RECT 17.3 2.35 17.56 2.61 ;
      RECT 21.07 1.9 21.33 2.16 ;
      RECT 21.06 1.925 21.33 2.12 ;
      RECT 21.055 1.925 21.06 2.119 ;
      RECT 20.985 1.92 21.055 2.111 ;
      RECT 20.9 1.907 20.985 2.094 ;
      RECT 20.896 1.899 20.9 2.084 ;
      RECT 20.81 1.892 20.896 2.074 ;
      RECT 20.801 1.884 20.81 2.064 ;
      RECT 20.715 1.877 20.801 2.052 ;
      RECT 20.695 1.868 20.715 2.038 ;
      RECT 20.64 1.863 20.695 2.03 ;
      RECT 20.63 1.857 20.64 2.024 ;
      RECT 20.61 1.855 20.63 2.02 ;
      RECT 20.602 1.854 20.61 2.016 ;
      RECT 20.516 1.846 20.602 2.005 ;
      RECT 20.43 1.832 20.516 1.985 ;
      RECT 20.37 1.82 20.43 1.97 ;
      RECT 20.36 1.815 20.37 1.965 ;
      RECT 20.31 1.815 20.36 1.967 ;
      RECT 20.263 1.817 20.31 1.971 ;
      RECT 20.177 1.824 20.263 1.976 ;
      RECT 20.091 1.832 20.177 1.982 ;
      RECT 20.005 1.841 20.091 1.988 ;
      RECT 19.946 1.847 20.005 1.993 ;
      RECT 19.86 1.852 19.946 1.999 ;
      RECT 19.785 1.857 19.86 2.005 ;
      RECT 19.746 1.859 19.785 2.01 ;
      RECT 19.66 1.856 19.746 2.015 ;
      RECT 19.575 1.854 19.66 2.022 ;
      RECT 19.543 1.853 19.575 2.025 ;
      RECT 19.457 1.852 19.543 2.026 ;
      RECT 19.371 1.851 19.457 2.027 ;
      RECT 19.285 1.85 19.371 2.027 ;
      RECT 19.199 1.849 19.285 2.028 ;
      RECT 19.113 1.848 19.199 2.029 ;
      RECT 19.027 1.847 19.113 2.03 ;
      RECT 18.941 1.846 19.027 2.03 ;
      RECT 18.855 1.845 18.941 2.031 ;
      RECT 18.805 1.845 18.855 2.032 ;
      RECT 18.791 1.846 18.805 2.032 ;
      RECT 18.705 1.853 18.791 2.033 ;
      RECT 18.631 1.864 18.705 2.034 ;
      RECT 18.545 1.873 18.631 2.035 ;
      RECT 18.51 1.88 18.545 2.05 ;
      RECT 18.485 1.883 18.51 2.08 ;
      RECT 18.46 1.892 18.485 2.109 ;
      RECT 18.45 1.903 18.46 2.129 ;
      RECT 18.44 1.911 18.45 2.143 ;
      RECT 18.435 1.917 18.44 2.153 ;
      RECT 18.41 1.934 18.435 2.17 ;
      RECT 18.395 1.956 18.41 2.198 ;
      RECT 18.365 1.982 18.395 2.228 ;
      RECT 18.345 2.011 18.365 2.258 ;
      RECT 18.34 2.026 18.345 2.275 ;
      RECT 18.32 2.041 18.34 2.29 ;
      RECT 18.31 2.059 18.32 2.308 ;
      RECT 18.3 2.07 18.31 2.323 ;
      RECT 18.25 2.102 18.3 2.349 ;
      RECT 18.245 2.132 18.25 2.369 ;
      RECT 18.235 2.145 18.245 2.375 ;
      RECT 18.226 2.155 18.235 2.383 ;
      RECT 18.215 2.166 18.226 2.391 ;
      RECT 18.21 2.176 18.215 2.397 ;
      RECT 18.195 2.197 18.21 2.404 ;
      RECT 18.18 2.227 18.195 2.412 ;
      RECT 18.145 2.257 18.18 2.418 ;
      RECT 18.12 2.275 18.145 2.425 ;
      RECT 18.07 2.283 18.12 2.434 ;
      RECT 18.045 2.288 18.07 2.443 ;
      RECT 17.99 2.294 18.045 2.453 ;
      RECT 17.985 2.299 17.99 2.461 ;
      RECT 17.971 2.302 17.985 2.463 ;
      RECT 17.885 2.314 17.971 2.475 ;
      RECT 17.875 2.326 17.885 2.488 ;
      RECT 17.79 2.339 17.875 2.5 ;
      RECT 17.746 2.356 17.79 2.514 ;
      RECT 17.66 2.373 17.746 2.53 ;
      RECT 17.63 2.387 17.66 2.544 ;
      RECT 17.62 2.392 17.63 2.549 ;
      RECT 17.56 2.395 17.62 2.558 ;
      RECT 20.45 2.665 20.71 2.925 ;
      RECT 20.45 2.665 20.73 2.778 ;
      RECT 20.45 2.665 20.755 2.745 ;
      RECT 20.45 2.665 20.76 2.725 ;
      RECT 20.5 2.44 20.78 2.72 ;
      RECT 20.055 3.175 20.315 3.435 ;
      RECT 20.045 3.032 20.24 3.373 ;
      RECT 20.04 3.14 20.255 3.365 ;
      RECT 20.035 3.19 20.315 3.355 ;
      RECT 20.025 3.267 20.315 3.34 ;
      RECT 20.045 3.115 20.255 3.373 ;
      RECT 20.055 2.99 20.24 3.435 ;
      RECT 20.055 2.885 20.22 3.435 ;
      RECT 20.065 2.872 20.22 3.435 ;
      RECT 20.065 2.83 20.21 3.435 ;
      RECT 20.07 2.755 20.21 3.435 ;
      RECT 20.1 2.405 20.21 3.435 ;
      RECT 20.105 2.135 20.23 2.758 ;
      RECT 20.075 2.71 20.23 2.758 ;
      RECT 20.09 2.512 20.21 3.435 ;
      RECT 20.08 2.622 20.23 2.758 ;
      RECT 20.105 2.135 20.245 2.615 ;
      RECT 20.105 2.135 20.265 2.49 ;
      RECT 20.07 2.135 20.33 2.395 ;
      RECT 19.54 2.44 19.82 2.72 ;
      RECT 19.525 2.44 19.82 2.7 ;
      RECT 17.58 3.305 17.84 3.565 ;
      RECT 19.365 3.16 19.625 3.42 ;
      RECT 19.345 3.18 19.625 3.395 ;
      RECT 19.302 3.18 19.345 3.394 ;
      RECT 19.216 3.181 19.302 3.391 ;
      RECT 19.13 3.182 19.216 3.387 ;
      RECT 19.055 3.184 19.13 3.384 ;
      RECT 19.032 3.185 19.055 3.382 ;
      RECT 18.946 3.186 19.032 3.38 ;
      RECT 18.86 3.187 18.946 3.377 ;
      RECT 18.836 3.188 18.86 3.375 ;
      RECT 18.75 3.19 18.836 3.372 ;
      RECT 18.665 3.192 18.75 3.373 ;
      RECT 18.608 3.193 18.665 3.379 ;
      RECT 18.522 3.195 18.608 3.389 ;
      RECT 18.436 3.198 18.522 3.402 ;
      RECT 18.35 3.2 18.436 3.414 ;
      RECT 18.336 3.201 18.35 3.421 ;
      RECT 18.25 3.202 18.336 3.429 ;
      RECT 18.21 3.204 18.25 3.438 ;
      RECT 18.201 3.205 18.21 3.441 ;
      RECT 18.115 3.213 18.201 3.447 ;
      RECT 18.095 3.222 18.115 3.455 ;
      RECT 18.01 3.237 18.095 3.463 ;
      RECT 17.95 3.26 18.01 3.474 ;
      RECT 17.94 3.272 17.95 3.479 ;
      RECT 17.9 3.282 17.94 3.483 ;
      RECT 17.845 3.299 17.9 3.491 ;
      RECT 17.84 3.309 17.845 3.495 ;
      RECT 18.906 2.44 18.965 2.837 ;
      RECT 18.82 2.44 19.025 2.828 ;
      RECT 18.815 2.47 19.025 2.823 ;
      RECT 18.781 2.47 19.025 2.821 ;
      RECT 18.695 2.47 19.025 2.815 ;
      RECT 18.65 2.47 19.045 2.793 ;
      RECT 18.65 2.47 19.065 2.748 ;
      RECT 18.61 2.47 19.065 2.738 ;
      RECT 18.82 2.44 19.1 2.72 ;
      RECT 18.555 2.44 18.815 2.7 ;
      RECT 17.74 1.92 18 2.18 ;
      RECT 17.795 1.88 18.1 2.16 ;
      RECT 17.795 1.855 17.97 2.18 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 11.805 6.745 13.245 6.915 ;
      RECT 11.805 2.395 11.965 6.915 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 11.805 2.395 12.44 2.565 ;
      RECT 11.07 5.855 11.42 6.205 ;
      RECT 11.14 2.705 11.315 6.205 ;
      RECT 11.065 2.705 11.415 3.055 ;
      RECT 0.53 3 0.81 3.28 ;
      RECT 0.5 3 0.81 3.265 ;
      RECT 0.495 2.963 0.755 3.263 ;
      RECT 0.49 2.964 0.755 3.257 ;
      RECT 0.485 2.967 0.755 3.25 ;
      RECT 0.48 3 0.81 3.243 ;
      RECT 0.45 2.97 0.755 3.23 ;
      RECT 0.45 2.997 0.775 3.23 ;
      RECT 0.45 2.987 0.77 3.23 ;
      RECT 0.45 2.972 0.765 3.23 ;
      RECT 0.55 2.962 0.755 3.28 ;
      RECT 0.55 2.957 0.745 3.28 ;
      RECT 0.55 2.955 0.73 3.28 ;
      RECT 0.55 1.42 0.725 3.28 ;
      RECT 10.46 1.34 10.81 1.69 ;
      RECT 0.55 1.42 10.81 1.595 ;
      RECT 6.24 2.455 6.475 2.715 ;
      RECT 9.385 2.235 9.55 2.495 ;
      RECT 9.29 2.225 9.305 2.495 ;
      RECT 7.89 1.795 7.93 1.935 ;
      RECT 9.305 2.23 9.385 2.495 ;
      RECT 9.25 2.225 9.29 2.461 ;
      RECT 9.236 2.225 9.25 2.461 ;
      RECT 9.15 2.23 9.236 2.463 ;
      RECT 9.105 2.237 9.15 2.465 ;
      RECT 9.075 2.237 9.105 2.467 ;
      RECT 9.05 2.232 9.075 2.469 ;
      RECT 9.02 2.228 9.05 2.478 ;
      RECT 9.01 2.225 9.02 2.49 ;
      RECT 9.005 2.225 9.01 2.498 ;
      RECT 9 2.225 9.005 2.503 ;
      RECT 8.99 2.224 9 2.513 ;
      RECT 8.985 2.223 8.99 2.523 ;
      RECT 8.97 2.222 8.985 2.528 ;
      RECT 8.942 2.219 8.97 2.555 ;
      RECT 8.856 2.211 8.942 2.555 ;
      RECT 8.77 2.2 8.856 2.555 ;
      RECT 8.73 2.185 8.77 2.555 ;
      RECT 8.69 2.159 8.73 2.555 ;
      RECT 8.685 2.141 8.69 2.367 ;
      RECT 8.675 2.137 8.685 2.357 ;
      RECT 8.66 2.127 8.675 2.344 ;
      RECT 8.64 2.111 8.66 2.329 ;
      RECT 8.625 2.096 8.64 2.314 ;
      RECT 8.615 2.085 8.625 2.304 ;
      RECT 8.59 2.069 8.615 2.293 ;
      RECT 8.585 2.056 8.59 2.283 ;
      RECT 8.58 2.052 8.585 2.278 ;
      RECT 8.525 2.038 8.58 2.256 ;
      RECT 8.486 2.019 8.525 2.22 ;
      RECT 8.4 1.993 8.486 2.173 ;
      RECT 8.396 1.975 8.4 2.139 ;
      RECT 8.31 1.956 8.396 2.117 ;
      RECT 8.305 1.938 8.31 2.095 ;
      RECT 8.3 1.936 8.305 2.093 ;
      RECT 8.29 1.935 8.3 2.088 ;
      RECT 8.23 1.922 8.29 2.074 ;
      RECT 8.185 1.9 8.23 2.053 ;
      RECT 8.125 1.877 8.185 2.032 ;
      RECT 8.061 1.852 8.125 2.007 ;
      RECT 7.975 1.822 8.061 1.976 ;
      RECT 7.96 1.802 7.975 1.955 ;
      RECT 7.93 1.797 7.96 1.946 ;
      RECT 7.877 1.795 7.89 1.935 ;
      RECT 7.791 1.795 7.877 1.937 ;
      RECT 7.705 1.795 7.791 1.939 ;
      RECT 7.685 1.795 7.705 1.943 ;
      RECT 7.64 1.797 7.685 1.954 ;
      RECT 7.6 1.807 7.64 1.97 ;
      RECT 7.596 1.816 7.6 1.978 ;
      RECT 7.51 1.836 7.596 1.994 ;
      RECT 7.5 1.855 7.51 2.012 ;
      RECT 7.495 1.857 7.5 2.015 ;
      RECT 7.485 1.861 7.495 2.018 ;
      RECT 7.465 1.866 7.485 2.028 ;
      RECT 7.435 1.876 7.465 2.048 ;
      RECT 7.43 1.883 7.435 2.062 ;
      RECT 7.42 1.887 7.43 2.069 ;
      RECT 7.405 1.895 7.42 2.08 ;
      RECT 7.395 1.905 7.405 2.091 ;
      RECT 7.385 1.912 7.395 2.099 ;
      RECT 7.36 1.925 7.385 2.114 ;
      RECT 7.296 1.961 7.36 2.153 ;
      RECT 7.21 2.024 7.296 2.217 ;
      RECT 7.175 2.075 7.21 2.27 ;
      RECT 7.17 2.092 7.175 2.287 ;
      RECT 7.155 2.101 7.17 2.294 ;
      RECT 7.135 2.116 7.155 2.308 ;
      RECT 7.13 2.127 7.135 2.318 ;
      RECT 7.11 2.14 7.13 2.328 ;
      RECT 7.105 2.15 7.11 2.338 ;
      RECT 7.09 2.155 7.105 2.347 ;
      RECT 7.08 2.165 7.09 2.358 ;
      RECT 7.05 2.182 7.08 2.375 ;
      RECT 7.04 2.2 7.05 2.393 ;
      RECT 7.025 2.211 7.04 2.404 ;
      RECT 6.985 2.235 7.025 2.42 ;
      RECT 6.95 2.269 6.985 2.437 ;
      RECT 6.92 2.292 6.95 2.449 ;
      RECT 6.905 2.302 6.92 2.458 ;
      RECT 6.865 2.312 6.905 2.469 ;
      RECT 6.845 2.323 6.865 2.481 ;
      RECT 6.84 2.327 6.845 2.488 ;
      RECT 6.825 2.331 6.84 2.493 ;
      RECT 6.815 2.336 6.825 2.498 ;
      RECT 6.81 2.339 6.815 2.501 ;
      RECT 6.78 2.345 6.81 2.508 ;
      RECT 6.745 2.355 6.78 2.522 ;
      RECT 6.685 2.37 6.745 2.542 ;
      RECT 6.63 2.39 6.685 2.566 ;
      RECT 6.601 2.405 6.63 2.584 ;
      RECT 6.515 2.425 6.601 2.609 ;
      RECT 6.51 2.44 6.515 2.629 ;
      RECT 6.5 2.443 6.51 2.63 ;
      RECT 6.475 2.45 6.5 2.715 ;
      RECT 6.89 3.685 6.9 3.875 ;
      RECT 5.15 3.56 5.43 3.84 ;
      RECT 8.195 2.5 8.2 2.985 ;
      RECT 8.09 2.5 8.15 2.76 ;
      RECT 8.415 3.47 8.42 3.545 ;
      RECT 8.405 3.337 8.415 3.58 ;
      RECT 8.395 3.172 8.405 3.601 ;
      RECT 8.39 3.042 8.395 3.617 ;
      RECT 8.38 2.932 8.39 3.633 ;
      RECT 8.375 2.831 8.38 3.65 ;
      RECT 8.37 2.813 8.375 3.66 ;
      RECT 8.365 2.795 8.37 3.67 ;
      RECT 8.355 2.77 8.365 3.685 ;
      RECT 8.35 2.75 8.355 3.7 ;
      RECT 8.33 2.5 8.35 3.725 ;
      RECT 8.315 2.5 8.33 3.758 ;
      RECT 8.285 2.5 8.315 3.78 ;
      RECT 8.265 2.5 8.285 3.794 ;
      RECT 8.245 2.5 8.265 3.31 ;
      RECT 8.26 3.377 8.265 3.799 ;
      RECT 8.255 3.407 8.26 3.801 ;
      RECT 8.25 3.42 8.255 3.804 ;
      RECT 8.245 3.43 8.25 3.808 ;
      RECT 8.24 2.5 8.245 3.228 ;
      RECT 8.24 3.44 8.245 3.81 ;
      RECT 8.235 2.5 8.24 3.205 ;
      RECT 8.225 3.462 8.24 3.81 ;
      RECT 8.22 2.5 8.235 3.15 ;
      RECT 8.215 3.487 8.225 3.81 ;
      RECT 8.215 2.5 8.22 3.095 ;
      RECT 8.205 2.5 8.215 3.043 ;
      RECT 8.21 3.5 8.215 3.811 ;
      RECT 8.205 3.512 8.21 3.812 ;
      RECT 8.2 2.5 8.205 3.003 ;
      RECT 8.2 3.525 8.205 3.813 ;
      RECT 8.185 3.54 8.2 3.814 ;
      RECT 8.19 2.5 8.195 2.965 ;
      RECT 8.185 2.5 8.19 2.93 ;
      RECT 8.18 2.5 8.185 2.905 ;
      RECT 8.175 3.567 8.185 3.816 ;
      RECT 8.17 2.5 8.18 2.863 ;
      RECT 8.17 3.585 8.175 3.817 ;
      RECT 8.165 2.5 8.17 2.823 ;
      RECT 8.165 3.592 8.17 3.818 ;
      RECT 8.16 2.5 8.165 2.795 ;
      RECT 8.155 3.61 8.165 3.819 ;
      RECT 8.15 2.5 8.16 2.775 ;
      RECT 8.145 3.63 8.155 3.821 ;
      RECT 8.135 3.647 8.145 3.822 ;
      RECT 8.1 3.67 8.135 3.825 ;
      RECT 8.045 3.688 8.1 3.831 ;
      RECT 7.959 3.696 8.045 3.84 ;
      RECT 7.873 3.707 7.959 3.851 ;
      RECT 7.787 3.717 7.873 3.862 ;
      RECT 7.701 3.727 7.787 3.874 ;
      RECT 7.615 3.737 7.701 3.885 ;
      RECT 7.595 3.743 7.615 3.891 ;
      RECT 7.515 3.745 7.595 3.895 ;
      RECT 7.51 3.744 7.515 3.9 ;
      RECT 7.502 3.743 7.51 3.9 ;
      RECT 7.416 3.739 7.502 3.898 ;
      RECT 7.33 3.731 7.416 3.895 ;
      RECT 7.244 3.722 7.33 3.891 ;
      RECT 7.158 3.714 7.244 3.888 ;
      RECT 7.072 3.706 7.158 3.884 ;
      RECT 6.986 3.697 7.072 3.881 ;
      RECT 6.9 3.689 6.986 3.877 ;
      RECT 6.845 3.682 6.89 3.875 ;
      RECT 6.76 3.675 6.845 3.873 ;
      RECT 6.686 3.667 6.76 3.869 ;
      RECT 6.6 3.659 6.686 3.866 ;
      RECT 6.597 3.655 6.6 3.864 ;
      RECT 6.511 3.651 6.597 3.863 ;
      RECT 6.425 3.643 6.511 3.86 ;
      RECT 6.34 3.638 6.425 3.857 ;
      RECT 6.254 3.635 6.34 3.854 ;
      RECT 6.168 3.633 6.254 3.851 ;
      RECT 6.082 3.63 6.168 3.848 ;
      RECT 5.996 3.627 6.082 3.845 ;
      RECT 5.91 3.624 5.996 3.842 ;
      RECT 5.834 3.622 5.91 3.839 ;
      RECT 5.748 3.619 5.834 3.836 ;
      RECT 5.662 3.616 5.748 3.834 ;
      RECT 5.576 3.614 5.662 3.831 ;
      RECT 5.49 3.611 5.576 3.828 ;
      RECT 5.43 3.602 5.49 3.826 ;
      RECT 7.94 3.22 8.015 3.48 ;
      RECT 7.92 3.2 7.925 3.48 ;
      RECT 7.24 2.985 7.345 3.28 ;
      RECT 1.685 2.96 1.755 3.22 ;
      RECT 7.58 2.835 7.585 3.206 ;
      RECT 7.57 2.89 7.575 3.206 ;
      RECT 7.875 2.06 7.935 2.32 ;
      RECT 7.93 3.215 7.94 3.48 ;
      RECT 7.925 3.205 7.93 3.48 ;
      RECT 7.845 3.152 7.92 3.48 ;
      RECT 7.87 2.06 7.875 2.34 ;
      RECT 7.86 2.06 7.87 2.36 ;
      RECT 7.845 2.06 7.86 2.39 ;
      RECT 7.83 2.06 7.845 2.433 ;
      RECT 7.825 3.095 7.845 3.48 ;
      RECT 7.815 2.06 7.83 2.47 ;
      RECT 7.81 3.075 7.825 3.48 ;
      RECT 7.81 2.06 7.815 2.493 ;
      RECT 7.8 2.06 7.81 2.518 ;
      RECT 7.77 3.042 7.81 3.48 ;
      RECT 7.775 2.06 7.8 2.568 ;
      RECT 7.77 2.06 7.775 2.623 ;
      RECT 7.765 2.06 7.77 2.665 ;
      RECT 7.755 3.005 7.77 3.48 ;
      RECT 7.76 2.06 7.765 2.708 ;
      RECT 7.755 2.06 7.76 2.773 ;
      RECT 7.75 2.06 7.755 2.795 ;
      RECT 7.75 2.993 7.755 3.345 ;
      RECT 7.745 2.06 7.75 2.863 ;
      RECT 7.745 2.985 7.75 3.328 ;
      RECT 7.74 2.06 7.745 2.908 ;
      RECT 7.735 2.967 7.745 3.305 ;
      RECT 7.735 2.06 7.74 2.945 ;
      RECT 7.725 2.06 7.735 3.285 ;
      RECT 7.72 2.06 7.725 3.268 ;
      RECT 7.715 2.06 7.72 3.253 ;
      RECT 7.71 2.06 7.715 3.238 ;
      RECT 7.69 2.06 7.71 3.228 ;
      RECT 7.685 2.06 7.69 3.218 ;
      RECT 7.675 2.06 7.685 3.214 ;
      RECT 7.67 2.337 7.675 3.213 ;
      RECT 7.665 2.36 7.67 3.212 ;
      RECT 7.66 2.39 7.665 3.211 ;
      RECT 7.655 2.417 7.66 3.21 ;
      RECT 7.65 2.445 7.655 3.21 ;
      RECT 7.645 2.472 7.65 3.21 ;
      RECT 7.64 2.492 7.645 3.21 ;
      RECT 7.635 2.52 7.64 3.21 ;
      RECT 7.625 2.562 7.635 3.21 ;
      RECT 7.615 2.607 7.625 3.209 ;
      RECT 7.61 2.66 7.615 3.208 ;
      RECT 7.605 2.692 7.61 3.207 ;
      RECT 7.6 2.712 7.605 3.206 ;
      RECT 7.595 2.75 7.6 3.206 ;
      RECT 7.59 2.772 7.595 3.206 ;
      RECT 7.585 2.797 7.59 3.206 ;
      RECT 7.575 2.862 7.58 3.206 ;
      RECT 7.56 2.922 7.57 3.206 ;
      RECT 7.545 2.932 7.56 3.206 ;
      RECT 7.525 2.942 7.545 3.206 ;
      RECT 7.495 2.947 7.525 3.203 ;
      RECT 7.435 2.957 7.495 3.2 ;
      RECT 7.415 2.966 7.435 3.205 ;
      RECT 7.39 2.972 7.415 3.218 ;
      RECT 7.37 2.977 7.39 3.233 ;
      RECT 7.345 2.982 7.37 3.28 ;
      RECT 7.216 2.984 7.24 3.28 ;
      RECT 7.13 2.979 7.216 3.28 ;
      RECT 7.09 2.976 7.13 3.28 ;
      RECT 7.04 2.978 7.09 3.26 ;
      RECT 7.01 2.982 7.04 3.26 ;
      RECT 6.931 2.992 7.01 3.26 ;
      RECT 6.845 3.007 6.931 3.261 ;
      RECT 6.795 3.017 6.845 3.262 ;
      RECT 6.787 3.02 6.795 3.262 ;
      RECT 6.701 3.022 6.787 3.263 ;
      RECT 6.615 3.026 6.701 3.263 ;
      RECT 6.529 3.03 6.615 3.264 ;
      RECT 6.443 3.033 6.529 3.265 ;
      RECT 6.357 3.037 6.443 3.265 ;
      RECT 6.271 3.041 6.357 3.266 ;
      RECT 6.185 3.044 6.271 3.267 ;
      RECT 6.099 3.048 6.185 3.267 ;
      RECT 6.013 3.052 6.099 3.268 ;
      RECT 5.927 3.056 6.013 3.269 ;
      RECT 5.841 3.059 5.927 3.269 ;
      RECT 5.755 3.063 5.841 3.27 ;
      RECT 5.725 3.065 5.755 3.27 ;
      RECT 5.639 3.068 5.725 3.271 ;
      RECT 5.553 3.072 5.639 3.272 ;
      RECT 5.467 3.076 5.553 3.273 ;
      RECT 5.381 3.079 5.467 3.273 ;
      RECT 5.295 3.083 5.381 3.274 ;
      RECT 5.26 3.088 5.295 3.275 ;
      RECT 5.205 3.098 5.26 3.282 ;
      RECT 5.18 3.11 5.205 3.292 ;
      RECT 5.145 3.123 5.18 3.3 ;
      RECT 5.105 3.14 5.145 3.323 ;
      RECT 5.085 3.153 5.105 3.35 ;
      RECT 5.055 3.165 5.085 3.378 ;
      RECT 5.05 3.173 5.055 3.398 ;
      RECT 5.045 3.176 5.05 3.408 ;
      RECT 4.995 3.188 5.045 3.442 ;
      RECT 4.985 3.203 4.995 3.475 ;
      RECT 4.975 3.209 4.985 3.488 ;
      RECT 4.965 3.216 4.975 3.5 ;
      RECT 4.94 3.229 4.965 3.518 ;
      RECT 4.925 3.244 4.94 3.54 ;
      RECT 4.915 3.252 4.925 3.556 ;
      RECT 4.9 3.261 4.915 3.571 ;
      RECT 4.89 3.271 4.9 3.585 ;
      RECT 4.871 3.284 4.89 3.602 ;
      RECT 4.785 3.329 4.871 3.667 ;
      RECT 4.77 3.374 4.785 3.725 ;
      RECT 4.765 3.383 4.77 3.738 ;
      RECT 4.755 3.39 4.765 3.743 ;
      RECT 4.75 3.395 4.755 3.747 ;
      RECT 4.73 3.405 4.75 3.754 ;
      RECT 4.705 3.425 4.73 3.768 ;
      RECT 4.67 3.45 4.705 3.788 ;
      RECT 4.655 3.473 4.67 3.803 ;
      RECT 4.645 3.483 4.655 3.808 ;
      RECT 4.635 3.491 4.645 3.815 ;
      RECT 4.625 3.5 4.635 3.821 ;
      RECT 4.605 3.512 4.625 3.823 ;
      RECT 4.595 3.525 4.605 3.825 ;
      RECT 4.57 3.54 4.595 3.828 ;
      RECT 4.55 3.557 4.57 3.832 ;
      RECT 4.51 3.585 4.55 3.838 ;
      RECT 4.445 3.632 4.51 3.847 ;
      RECT 4.43 3.665 4.445 3.855 ;
      RECT 4.425 3.672 4.43 3.857 ;
      RECT 4.375 3.697 4.425 3.862 ;
      RECT 4.36 3.721 4.375 3.869 ;
      RECT 4.31 3.726 4.36 3.87 ;
      RECT 4.224 3.73 4.31 3.87 ;
      RECT 4.138 3.73 4.224 3.87 ;
      RECT 4.052 3.73 4.138 3.871 ;
      RECT 3.966 3.73 4.052 3.871 ;
      RECT 3.88 3.73 3.966 3.871 ;
      RECT 3.814 3.73 3.88 3.871 ;
      RECT 3.728 3.73 3.814 3.872 ;
      RECT 3.642 3.73 3.728 3.872 ;
      RECT 3.556 3.731 3.642 3.873 ;
      RECT 3.47 3.731 3.556 3.873 ;
      RECT 3.384 3.731 3.47 3.873 ;
      RECT 3.298 3.731 3.384 3.874 ;
      RECT 3.212 3.731 3.298 3.874 ;
      RECT 3.126 3.732 3.212 3.875 ;
      RECT 3.04 3.732 3.126 3.875 ;
      RECT 3.02 3.732 3.04 3.875 ;
      RECT 2.934 3.732 3.02 3.875 ;
      RECT 2.848 3.732 2.934 3.875 ;
      RECT 2.762 3.733 2.848 3.875 ;
      RECT 2.676 3.733 2.762 3.875 ;
      RECT 2.59 3.733 2.676 3.875 ;
      RECT 2.504 3.734 2.59 3.875 ;
      RECT 2.418 3.734 2.504 3.875 ;
      RECT 2.332 3.734 2.418 3.875 ;
      RECT 2.246 3.734 2.332 3.875 ;
      RECT 2.16 3.735 2.246 3.875 ;
      RECT 2.11 3.732 2.16 3.875 ;
      RECT 2.1 3.73 2.11 3.874 ;
      RECT 2.096 3.73 2.1 3.873 ;
      RECT 2.01 3.725 2.096 3.868 ;
      RECT 1.988 3.718 2.01 3.862 ;
      RECT 1.902 3.709 1.988 3.856 ;
      RECT 1.816 3.696 1.902 3.847 ;
      RECT 1.73 3.682 1.816 3.837 ;
      RECT 1.685 3.672 1.73 3.83 ;
      RECT 1.665 2.96 1.685 3.238 ;
      RECT 1.665 3.665 1.685 3.826 ;
      RECT 1.635 2.96 1.665 3.26 ;
      RECT 1.625 3.632 1.665 3.823 ;
      RECT 1.62 2.96 1.635 3.28 ;
      RECT 1.62 3.597 1.625 3.821 ;
      RECT 1.615 2.96 1.62 3.405 ;
      RECT 1.615 3.557 1.62 3.821 ;
      RECT 1.605 2.96 1.615 3.821 ;
      RECT 1.53 2.96 1.605 3.815 ;
      RECT 1.5 2.96 1.53 3.805 ;
      RECT 1.495 2.96 1.5 3.797 ;
      RECT 1.49 3.002 1.495 3.79 ;
      RECT 1.48 3.071 1.49 3.781 ;
      RECT 1.475 3.141 1.48 3.733 ;
      RECT 1.47 3.205 1.475 3.63 ;
      RECT 1.465 3.24 1.47 3.585 ;
      RECT 1.463 3.277 1.465 3.477 ;
      RECT 1.46 3.285 1.463 3.47 ;
      RECT 1.455 3.35 1.46 3.413 ;
      RECT 5.53 2.44 5.81 2.72 ;
      RECT 5.52 2.44 5.81 2.583 ;
      RECT 5.475 2.305 5.735 2.565 ;
      RECT 5.475 2.42 5.79 2.565 ;
      RECT 5.475 2.39 5.785 2.565 ;
      RECT 5.475 2.377 5.775 2.565 ;
      RECT 5.475 2.367 5.77 2.565 ;
      RECT 1.45 2.35 1.71 2.61 ;
      RECT 5.22 1.9 5.48 2.16 ;
      RECT 5.21 1.925 5.48 2.12 ;
      RECT 5.205 1.925 5.21 2.119 ;
      RECT 5.135 1.92 5.205 2.111 ;
      RECT 5.05 1.907 5.135 2.094 ;
      RECT 5.046 1.899 5.05 2.084 ;
      RECT 4.96 1.892 5.046 2.074 ;
      RECT 4.951 1.884 4.96 2.064 ;
      RECT 4.865 1.877 4.951 2.052 ;
      RECT 4.845 1.868 4.865 2.038 ;
      RECT 4.79 1.863 4.845 2.03 ;
      RECT 4.78 1.857 4.79 2.024 ;
      RECT 4.76 1.855 4.78 2.02 ;
      RECT 4.752 1.854 4.76 2.016 ;
      RECT 4.666 1.846 4.752 2.005 ;
      RECT 4.58 1.832 4.666 1.985 ;
      RECT 4.52 1.82 4.58 1.97 ;
      RECT 4.51 1.815 4.52 1.965 ;
      RECT 4.46 1.815 4.51 1.967 ;
      RECT 4.413 1.817 4.46 1.971 ;
      RECT 4.327 1.824 4.413 1.976 ;
      RECT 4.241 1.832 4.327 1.982 ;
      RECT 4.155 1.841 4.241 1.988 ;
      RECT 4.096 1.847 4.155 1.993 ;
      RECT 4.01 1.852 4.096 1.999 ;
      RECT 3.935 1.857 4.01 2.005 ;
      RECT 3.896 1.859 3.935 2.01 ;
      RECT 3.81 1.856 3.896 2.015 ;
      RECT 3.725 1.854 3.81 2.022 ;
      RECT 3.693 1.853 3.725 2.025 ;
      RECT 3.607 1.852 3.693 2.026 ;
      RECT 3.521 1.851 3.607 2.027 ;
      RECT 3.435 1.85 3.521 2.027 ;
      RECT 3.349 1.849 3.435 2.028 ;
      RECT 3.263 1.848 3.349 2.029 ;
      RECT 3.177 1.847 3.263 2.03 ;
      RECT 3.091 1.846 3.177 2.03 ;
      RECT 3.005 1.845 3.091 2.031 ;
      RECT 2.955 1.845 3.005 2.032 ;
      RECT 2.941 1.846 2.955 2.032 ;
      RECT 2.855 1.853 2.941 2.033 ;
      RECT 2.781 1.864 2.855 2.034 ;
      RECT 2.695 1.873 2.781 2.035 ;
      RECT 2.66 1.88 2.695 2.05 ;
      RECT 2.635 1.883 2.66 2.08 ;
      RECT 2.61 1.892 2.635 2.109 ;
      RECT 2.6 1.903 2.61 2.129 ;
      RECT 2.59 1.911 2.6 2.143 ;
      RECT 2.585 1.917 2.59 2.153 ;
      RECT 2.56 1.934 2.585 2.17 ;
      RECT 2.545 1.956 2.56 2.198 ;
      RECT 2.515 1.982 2.545 2.228 ;
      RECT 2.495 2.011 2.515 2.258 ;
      RECT 2.49 2.026 2.495 2.275 ;
      RECT 2.47 2.041 2.49 2.29 ;
      RECT 2.46 2.059 2.47 2.308 ;
      RECT 2.45 2.07 2.46 2.323 ;
      RECT 2.4 2.102 2.45 2.349 ;
      RECT 2.395 2.132 2.4 2.369 ;
      RECT 2.385 2.145 2.395 2.375 ;
      RECT 2.376 2.155 2.385 2.383 ;
      RECT 2.365 2.166 2.376 2.391 ;
      RECT 2.36 2.176 2.365 2.397 ;
      RECT 2.345 2.197 2.36 2.404 ;
      RECT 2.33 2.227 2.345 2.412 ;
      RECT 2.295 2.257 2.33 2.418 ;
      RECT 2.27 2.275 2.295 2.425 ;
      RECT 2.22 2.283 2.27 2.434 ;
      RECT 2.195 2.288 2.22 2.443 ;
      RECT 2.14 2.294 2.195 2.453 ;
      RECT 2.135 2.299 2.14 2.461 ;
      RECT 2.121 2.302 2.135 2.463 ;
      RECT 2.035 2.314 2.121 2.475 ;
      RECT 2.025 2.326 2.035 2.488 ;
      RECT 1.94 2.339 2.025 2.5 ;
      RECT 1.896 2.356 1.94 2.514 ;
      RECT 1.81 2.373 1.896 2.53 ;
      RECT 1.78 2.387 1.81 2.544 ;
      RECT 1.77 2.392 1.78 2.549 ;
      RECT 1.71 2.395 1.77 2.558 ;
      RECT 4.6 2.665 4.86 2.925 ;
      RECT 4.6 2.665 4.88 2.778 ;
      RECT 4.6 2.665 4.905 2.745 ;
      RECT 4.6 2.665 4.91 2.725 ;
      RECT 4.65 2.44 4.93 2.72 ;
      RECT 4.205 3.175 4.465 3.435 ;
      RECT 4.195 3.032 4.39 3.373 ;
      RECT 4.19 3.14 4.405 3.365 ;
      RECT 4.185 3.19 4.465 3.355 ;
      RECT 4.175 3.267 4.465 3.34 ;
      RECT 4.195 3.115 4.405 3.373 ;
      RECT 4.205 2.99 4.39 3.435 ;
      RECT 4.205 2.885 4.37 3.435 ;
      RECT 4.215 2.872 4.37 3.435 ;
      RECT 4.215 2.83 4.36 3.435 ;
      RECT 4.22 2.755 4.36 3.435 ;
      RECT 4.25 2.405 4.36 3.435 ;
      RECT 4.255 2.135 4.38 2.758 ;
      RECT 4.225 2.71 4.38 2.758 ;
      RECT 4.24 2.512 4.36 3.435 ;
      RECT 4.23 2.622 4.38 2.758 ;
      RECT 4.255 2.135 4.395 2.615 ;
      RECT 4.255 2.135 4.415 2.49 ;
      RECT 4.22 2.135 4.48 2.395 ;
      RECT 3.69 2.44 3.97 2.72 ;
      RECT 3.675 2.44 3.97 2.7 ;
      RECT 1.73 3.305 1.99 3.565 ;
      RECT 3.515 3.16 3.775 3.42 ;
      RECT 3.495 3.18 3.775 3.395 ;
      RECT 3.452 3.18 3.495 3.394 ;
      RECT 3.366 3.181 3.452 3.391 ;
      RECT 3.28 3.182 3.366 3.387 ;
      RECT 3.205 3.184 3.28 3.384 ;
      RECT 3.182 3.185 3.205 3.382 ;
      RECT 3.096 3.186 3.182 3.38 ;
      RECT 3.01 3.187 3.096 3.377 ;
      RECT 2.986 3.188 3.01 3.375 ;
      RECT 2.9 3.19 2.986 3.372 ;
      RECT 2.815 3.192 2.9 3.373 ;
      RECT 2.758 3.193 2.815 3.379 ;
      RECT 2.672 3.195 2.758 3.389 ;
      RECT 2.586 3.198 2.672 3.402 ;
      RECT 2.5 3.2 2.586 3.414 ;
      RECT 2.486 3.201 2.5 3.421 ;
      RECT 2.4 3.202 2.486 3.429 ;
      RECT 2.36 3.204 2.4 3.438 ;
      RECT 2.351 3.205 2.36 3.441 ;
      RECT 2.265 3.213 2.351 3.447 ;
      RECT 2.245 3.222 2.265 3.455 ;
      RECT 2.16 3.237 2.245 3.463 ;
      RECT 2.1 3.26 2.16 3.474 ;
      RECT 2.09 3.272 2.1 3.479 ;
      RECT 2.05 3.282 2.09 3.483 ;
      RECT 1.995 3.299 2.05 3.491 ;
      RECT 1.99 3.309 1.995 3.495 ;
      RECT 3.056 2.44 3.115 2.837 ;
      RECT 2.97 2.44 3.175 2.828 ;
      RECT 2.965 2.47 3.175 2.823 ;
      RECT 2.931 2.47 3.175 2.821 ;
      RECT 2.845 2.47 3.175 2.815 ;
      RECT 2.8 2.47 3.195 2.793 ;
      RECT 2.8 2.47 3.215 2.748 ;
      RECT 2.76 2.47 3.215 2.738 ;
      RECT 2.97 2.44 3.25 2.72 ;
      RECT 2.705 2.44 2.965 2.7 ;
      RECT 1.89 1.92 2.15 2.18 ;
      RECT 1.945 1.88 2.25 2.16 ;
      RECT 1.945 1.855 2.12 2.18 ;
    LAYER via1 ;
      RECT 78.755 2.265 78.905 2.415 ;
      RECT 76.41 6.74 76.56 6.89 ;
      RECT 76.395 2.065 76.545 2.215 ;
      RECT 75.605 2.45 75.755 2.6 ;
      RECT 75.605 6.37 75.755 6.52 ;
      RECT 74.57 5.955 74.72 6.105 ;
      RECT 74.565 2.805 74.715 2.955 ;
      RECT 73.96 1.44 74.11 1.59 ;
      RECT 72.745 2.29 72.895 2.44 ;
      RECT 72.625 2.86 72.775 3.01 ;
      RECT 71.545 2.555 71.695 2.705 ;
      RECT 71.21 3.275 71.36 3.425 ;
      RECT 71.13 2.115 71.28 2.265 ;
      RECT 69.695 2.51 69.845 2.66 ;
      RECT 68.93 2.36 69.08 2.51 ;
      RECT 68.675 1.955 68.825 2.105 ;
      RECT 68.055 2.72 68.205 2.87 ;
      RECT 67.675 2.19 67.825 2.34 ;
      RECT 67.66 3.23 67.81 3.38 ;
      RECT 67.13 2.495 67.28 2.645 ;
      RECT 66.97 3.215 67.12 3.365 ;
      RECT 66.16 2.495 66.31 2.645 ;
      RECT 65.345 1.975 65.495 2.125 ;
      RECT 65.185 3.36 65.335 3.51 ;
      RECT 64.95 3.015 65.1 3.165 ;
      RECT 64.905 2.405 65.055 2.555 ;
      RECT 63.905 3.025 64.055 3.175 ;
      RECT 62.93 0.985 63.08 1.135 ;
      RECT 60.56 6.74 60.71 6.89 ;
      RECT 60.545 2.065 60.695 2.215 ;
      RECT 59.755 2.45 59.905 2.6 ;
      RECT 59.755 6.37 59.905 6.52 ;
      RECT 58.72 5.955 58.87 6.105 ;
      RECT 58.715 2.805 58.865 2.955 ;
      RECT 58.11 1.44 58.26 1.59 ;
      RECT 56.895 2.29 57.045 2.44 ;
      RECT 56.775 2.86 56.925 3.01 ;
      RECT 55.695 2.555 55.845 2.705 ;
      RECT 55.36 3.275 55.51 3.425 ;
      RECT 55.28 2.115 55.43 2.265 ;
      RECT 53.845 2.51 53.995 2.66 ;
      RECT 53.08 2.36 53.23 2.51 ;
      RECT 52.825 1.955 52.975 2.105 ;
      RECT 52.205 2.72 52.355 2.87 ;
      RECT 51.825 2.19 51.975 2.34 ;
      RECT 51.81 3.23 51.96 3.38 ;
      RECT 51.28 2.495 51.43 2.645 ;
      RECT 51.12 3.215 51.27 3.365 ;
      RECT 50.31 2.495 50.46 2.645 ;
      RECT 49.495 1.975 49.645 2.125 ;
      RECT 49.335 3.36 49.485 3.51 ;
      RECT 49.1 3.015 49.25 3.165 ;
      RECT 49.055 2.405 49.205 2.555 ;
      RECT 48.055 3.025 48.205 3.175 ;
      RECT 47.08 0.985 47.23 1.135 ;
      RECT 44.71 6.74 44.86 6.89 ;
      RECT 44.695 2.065 44.845 2.215 ;
      RECT 43.905 2.45 44.055 2.6 ;
      RECT 43.905 6.37 44.055 6.52 ;
      RECT 42.87 5.955 43.02 6.105 ;
      RECT 42.865 2.805 43.015 2.955 ;
      RECT 42.26 1.44 42.41 1.59 ;
      RECT 41.045 2.29 41.195 2.44 ;
      RECT 40.925 2.86 41.075 3.01 ;
      RECT 39.845 2.555 39.995 2.705 ;
      RECT 39.51 3.275 39.66 3.425 ;
      RECT 39.43 2.115 39.58 2.265 ;
      RECT 37.995 2.51 38.145 2.66 ;
      RECT 37.23 2.36 37.38 2.51 ;
      RECT 36.975 1.955 37.125 2.105 ;
      RECT 36.355 2.72 36.505 2.87 ;
      RECT 35.975 2.19 36.125 2.34 ;
      RECT 35.96 3.23 36.11 3.38 ;
      RECT 35.43 2.495 35.58 2.645 ;
      RECT 35.27 3.215 35.42 3.365 ;
      RECT 34.46 2.495 34.61 2.645 ;
      RECT 33.645 1.975 33.795 2.125 ;
      RECT 33.485 3.36 33.635 3.51 ;
      RECT 33.25 3.015 33.4 3.165 ;
      RECT 33.205 2.405 33.355 2.555 ;
      RECT 32.205 3.025 32.355 3.175 ;
      RECT 31.23 0.985 31.38 1.135 ;
      RECT 28.86 6.74 29.01 6.89 ;
      RECT 28.845 2.065 28.995 2.215 ;
      RECT 28.055 2.45 28.205 2.6 ;
      RECT 28.055 6.37 28.205 6.52 ;
      RECT 27.02 5.955 27.17 6.105 ;
      RECT 27.015 2.805 27.165 2.955 ;
      RECT 26.41 1.44 26.56 1.59 ;
      RECT 25.195 2.29 25.345 2.44 ;
      RECT 25.075 2.86 25.225 3.01 ;
      RECT 23.995 2.555 24.145 2.705 ;
      RECT 23.66 3.275 23.81 3.425 ;
      RECT 23.58 2.115 23.73 2.265 ;
      RECT 22.145 2.51 22.295 2.66 ;
      RECT 21.38 2.36 21.53 2.51 ;
      RECT 21.125 1.955 21.275 2.105 ;
      RECT 20.505 2.72 20.655 2.87 ;
      RECT 20.125 2.19 20.275 2.34 ;
      RECT 20.11 3.23 20.26 3.38 ;
      RECT 19.58 2.495 19.73 2.645 ;
      RECT 19.42 3.215 19.57 3.365 ;
      RECT 18.61 2.495 18.76 2.645 ;
      RECT 17.795 1.975 17.945 2.125 ;
      RECT 17.635 3.36 17.785 3.51 ;
      RECT 17.4 3.015 17.55 3.165 ;
      RECT 17.355 2.405 17.505 2.555 ;
      RECT 16.355 3.025 16.505 3.175 ;
      RECT 15.38 0.985 15.53 1.135 ;
      RECT 13.01 6.74 13.16 6.89 ;
      RECT 12.995 2.065 13.145 2.215 ;
      RECT 12.205 2.45 12.355 2.6 ;
      RECT 12.205 6.37 12.355 6.52 ;
      RECT 11.17 5.955 11.32 6.105 ;
      RECT 11.165 2.805 11.315 2.955 ;
      RECT 10.56 1.44 10.71 1.59 ;
      RECT 9.345 2.29 9.495 2.44 ;
      RECT 9.225 2.86 9.375 3.01 ;
      RECT 8.145 2.555 8.295 2.705 ;
      RECT 7.81 3.275 7.96 3.425 ;
      RECT 7.73 2.115 7.88 2.265 ;
      RECT 6.295 2.51 6.445 2.66 ;
      RECT 5.53 2.36 5.68 2.51 ;
      RECT 5.275 1.955 5.425 2.105 ;
      RECT 4.655 2.72 4.805 2.87 ;
      RECT 4.275 2.19 4.425 2.34 ;
      RECT 4.26 3.23 4.41 3.38 ;
      RECT 3.73 2.495 3.88 2.645 ;
      RECT 3.57 3.215 3.72 3.365 ;
      RECT 2.76 2.495 2.91 2.645 ;
      RECT 1.945 1.975 2.095 2.125 ;
      RECT 1.785 3.36 1.935 3.51 ;
      RECT 1.55 3.015 1.7 3.165 ;
      RECT 1.505 2.405 1.655 2.555 ;
      RECT 0.505 3.025 0.655 3.175 ;
    LAYER met1 ;
      RECT 63.655 1.26 73.315 1.74 ;
      RECT 47.805 1.26 57.465 1.74 ;
      RECT 31.955 1.26 41.615 1.74 ;
      RECT 16.105 1.26 25.765 1.74 ;
      RECT 0.255 1.26 9.915 1.74 ;
      RECT 63.655 1.26 73.37 1.59 ;
      RECT 47.805 1.26 57.52 1.59 ;
      RECT 31.955 1.26 41.67 1.59 ;
      RECT 16.105 1.26 25.82 1.59 ;
      RECT 0.255 1.26 9.97 1.59 ;
      RECT 63.77 0 73.485 1.585 ;
      RECT 47.92 0 57.635 1.585 ;
      RECT 32.07 0 41.785 1.585 ;
      RECT 16.22 0 25.935 1.585 ;
      RECT 0.37 0 10.085 1.585 ;
      RECT 0 0 79.25 0.305 ;
      RECT 63.19 4.135 63.69 4.75 ;
      RECT 0.005 4.305 79.25 4.745 ;
      RECT 0.255 4.135 79.25 4.745 ;
      RECT 63.655 3.98 73.315 4.745 ;
      RECT 47.34 4.13 57.465 4.745 ;
      RECT 47.805 3.98 57.465 4.745 ;
      RECT 31.955 3.98 41.615 4.745 ;
      RECT 16.105 3.98 25.765 4.745 ;
      RECT 0.255 3.98 9.915 4.745 ;
      RECT 78.65 2.365 78.94 2.595 ;
      RECT 78.655 2.165 79.005 2.515 ;
      RECT 78.71 0.885 78.88 2.595 ;
      RECT 78.65 0.885 78.94 1.115 ;
      RECT 78.65 7.765 78.94 7.995 ;
      RECT 78.71 6.285 78.88 7.995 ;
      RECT 78.65 6.285 78.94 6.515 ;
      RECT 78.24 2.735 78.57 2.965 ;
      RECT 78.24 2.765 78.74 2.935 ;
      RECT 78.24 2.395 78.43 2.965 ;
      RECT 77.66 2.365 77.95 2.595 ;
      RECT 77.66 2.395 78.43 2.565 ;
      RECT 77.72 0.885 77.89 2.595 ;
      RECT 77.66 0.885 77.95 1.115 ;
      RECT 77.66 7.765 77.95 7.995 ;
      RECT 77.72 6.285 77.89 7.995 ;
      RECT 77.66 6.285 77.95 6.515 ;
      RECT 77.66 6.325 78.51 6.485 ;
      RECT 78.34 5.915 78.51 6.485 ;
      RECT 77.66 6.32 78.05 6.485 ;
      RECT 78.28 5.915 78.57 6.145 ;
      RECT 78.28 5.945 78.74 6.115 ;
      RECT 77.29 2.735 77.58 2.965 ;
      RECT 77.29 2.765 77.75 2.935 ;
      RECT 77.35 1.655 77.515 2.965 ;
      RECT 75.865 1.625 76.155 1.855 ;
      RECT 75.865 1.655 77.515 1.825 ;
      RECT 75.925 0.885 76.095 1.855 ;
      RECT 75.865 0.885 76.155 1.115 ;
      RECT 75.865 7.765 76.155 7.995 ;
      RECT 75.925 7.025 76.095 7.995 ;
      RECT 75.925 7.12 77.515 7.29 ;
      RECT 77.345 5.915 77.515 7.29 ;
      RECT 75.865 7.025 76.155 7.255 ;
      RECT 77.29 5.915 77.58 6.145 ;
      RECT 77.29 5.945 77.75 6.115 ;
      RECT 76.295 1.965 76.645 2.315 ;
      RECT 76.125 2.025 76.645 2.195 ;
      RECT 76.32 6.655 76.645 6.98 ;
      RECT 76.295 6.655 76.645 6.885 ;
      RECT 76.125 6.685 76.645 6.855 ;
      RECT 75.52 2.365 75.84 2.685 ;
      RECT 75.49 2.365 75.84 2.595 ;
      RECT 73.96 2.395 75.84 2.565 ;
      RECT 73.96 1.34 74.13 2.565 ;
      RECT 73.86 1.34 74.21 1.69 ;
      RECT 75.52 6.28 75.84 6.605 ;
      RECT 75.49 6.285 75.84 6.515 ;
      RECT 75.32 6.315 75.84 6.485 ;
      RECT 74.465 2.705 74.815 3.055 ;
      RECT 74.465 2.765 74.955 2.935 ;
      RECT 74.47 5.855 74.82 6.205 ;
      RECT 74.47 5.945 74.955 6.115 ;
      RECT 72.155 2.465 72.34 2.675 ;
      RECT 72.145 2.47 72.355 2.668 ;
      RECT 72.145 2.47 72.441 2.645 ;
      RECT 72.145 2.47 72.5 2.62 ;
      RECT 72.145 2.47 72.555 2.6 ;
      RECT 72.145 2.47 72.565 2.588 ;
      RECT 72.145 2.47 72.76 2.527 ;
      RECT 72.145 2.47 72.79 2.51 ;
      RECT 72.145 2.47 72.81 2.5 ;
      RECT 72.69 2.235 72.95 2.495 ;
      RECT 72.675 2.325 72.69 2.542 ;
      RECT 72.21 2.457 72.95 2.495 ;
      RECT 72.661 2.336 72.675 2.548 ;
      RECT 72.25 2.45 72.95 2.495 ;
      RECT 72.575 2.376 72.661 2.567 ;
      RECT 72.5 2.437 72.95 2.495 ;
      RECT 72.57 2.412 72.575 2.584 ;
      RECT 72.555 2.422 72.95 2.495 ;
      RECT 72.565 2.417 72.57 2.586 ;
      RECT 72.86 2.922 72.865 3.014 ;
      RECT 72.855 2.9 72.86 3.031 ;
      RECT 72.85 2.89 72.855 3.043 ;
      RECT 72.84 2.881 72.85 3.053 ;
      RECT 72.835 2.876 72.84 3.061 ;
      RECT 72.83 2.735 72.835 3.064 ;
      RECT 72.796 2.735 72.83 3.075 ;
      RECT 72.71 2.735 72.796 3.11 ;
      RECT 72.63 2.735 72.71 3.158 ;
      RECT 72.601 2.735 72.63 3.182 ;
      RECT 72.515 2.735 72.601 3.188 ;
      RECT 72.51 2.919 72.515 3.193 ;
      RECT 72.475 2.93 72.51 3.196 ;
      RECT 72.45 2.945 72.475 3.2 ;
      RECT 72.436 2.954 72.45 3.202 ;
      RECT 72.35 2.981 72.436 3.208 ;
      RECT 72.285 3.022 72.35 3.217 ;
      RECT 72.27 3.042 72.285 3.222 ;
      RECT 72.24 3.052 72.27 3.225 ;
      RECT 72.235 3.062 72.24 3.228 ;
      RECT 72.205 3.067 72.235 3.23 ;
      RECT 72.185 3.072 72.205 3.234 ;
      RECT 72.1 3.075 72.185 3.241 ;
      RECT 72.085 3.072 72.1 3.247 ;
      RECT 72.075 3.069 72.085 3.249 ;
      RECT 72.055 3.066 72.075 3.251 ;
      RECT 72.035 3.062 72.055 3.252 ;
      RECT 72.02 3.058 72.035 3.254 ;
      RECT 72.01 3.055 72.02 3.255 ;
      RECT 71.97 3.049 72.01 3.253 ;
      RECT 71.96 3.044 71.97 3.251 ;
      RECT 71.945 3.041 71.96 3.247 ;
      RECT 71.92 3.036 71.945 3.24 ;
      RECT 71.87 3.027 71.92 3.228 ;
      RECT 71.8 3.013 71.87 3.21 ;
      RECT 71.742 2.998 71.8 3.192 ;
      RECT 71.656 2.981 71.742 3.172 ;
      RECT 71.57 2.96 71.656 3.147 ;
      RECT 71.52 2.945 71.57 3.128 ;
      RECT 71.516 2.939 71.52 3.12 ;
      RECT 71.43 2.929 71.516 3.107 ;
      RECT 71.395 2.914 71.43 3.09 ;
      RECT 71.38 2.907 71.395 3.083 ;
      RECT 71.32 2.895 71.38 3.071 ;
      RECT 71.3 2.882 71.32 3.059 ;
      RECT 71.26 2.873 71.3 3.051 ;
      RECT 71.255 2.865 71.26 3.044 ;
      RECT 71.175 2.855 71.255 3.03 ;
      RECT 71.16 2.842 71.175 3.015 ;
      RECT 71.155 2.84 71.16 3.013 ;
      RECT 71.076 2.828 71.155 3 ;
      RECT 70.99 2.803 71.076 2.975 ;
      RECT 70.975 2.772 70.99 2.96 ;
      RECT 70.96 2.747 70.975 2.956 ;
      RECT 70.945 2.74 70.96 2.952 ;
      RECT 70.77 2.745 70.775 2.948 ;
      RECT 70.765 2.75 70.77 2.943 ;
      RECT 70.775 2.74 70.945 2.95 ;
      RECT 71.49 2.5 71.595 2.76 ;
      RECT 72.305 2.025 72.31 2.25 ;
      RECT 72.435 2.025 72.49 2.235 ;
      RECT 72.49 2.03 72.5 2.228 ;
      RECT 72.396 2.025 72.435 2.238 ;
      RECT 72.31 2.025 72.396 2.245 ;
      RECT 72.29 2.03 72.305 2.251 ;
      RECT 72.28 2.07 72.29 2.253 ;
      RECT 72.25 2.08 72.28 2.255 ;
      RECT 72.245 2.085 72.25 2.257 ;
      RECT 72.22 2.09 72.245 2.259 ;
      RECT 72.205 2.095 72.22 2.261 ;
      RECT 72.19 2.097 72.205 2.263 ;
      RECT 72.185 2.102 72.19 2.265 ;
      RECT 72.135 2.11 72.185 2.268 ;
      RECT 72.11 2.119 72.135 2.273 ;
      RECT 72.1 2.126 72.11 2.278 ;
      RECT 72.095 2.129 72.1 2.282 ;
      RECT 72.075 2.132 72.095 2.291 ;
      RECT 72.045 2.14 72.075 2.311 ;
      RECT 72.016 2.153 72.045 2.333 ;
      RECT 71.93 2.187 72.016 2.377 ;
      RECT 71.925 2.213 71.93 2.415 ;
      RECT 71.92 2.217 71.925 2.424 ;
      RECT 71.885 2.23 71.92 2.457 ;
      RECT 71.875 2.244 71.885 2.495 ;
      RECT 71.87 2.248 71.875 2.508 ;
      RECT 71.865 2.252 71.87 2.513 ;
      RECT 71.855 2.26 71.865 2.525 ;
      RECT 71.85 2.267 71.855 2.54 ;
      RECT 71.825 2.28 71.85 2.565 ;
      RECT 71.785 2.309 71.825 2.62 ;
      RECT 71.77 2.334 71.785 2.675 ;
      RECT 71.76 2.345 71.77 2.698 ;
      RECT 71.755 2.352 71.76 2.71 ;
      RECT 71.75 2.356 71.755 2.718 ;
      RECT 71.695 2.384 71.75 2.76 ;
      RECT 71.675 2.42 71.695 2.76 ;
      RECT 71.66 2.435 71.675 2.76 ;
      RECT 71.605 2.467 71.66 2.76 ;
      RECT 71.595 2.497 71.605 2.76 ;
      RECT 71.205 2.112 71.39 2.35 ;
      RECT 71.19 2.114 71.4 2.345 ;
      RECT 71.075 2.06 71.335 2.32 ;
      RECT 71.07 2.097 71.335 2.274 ;
      RECT 71.065 2.107 71.335 2.271 ;
      RECT 71.06 2.147 71.4 2.265 ;
      RECT 71.055 2.18 71.4 2.255 ;
      RECT 71.065 2.122 71.415 2.193 ;
      RECT 71.362 3.22 71.375 3.75 ;
      RECT 71.276 3.22 71.375 3.749 ;
      RECT 71.276 3.22 71.38 3.748 ;
      RECT 71.19 3.22 71.38 3.746 ;
      RECT 71.185 3.22 71.38 3.743 ;
      RECT 71.185 3.22 71.39 3.741 ;
      RECT 71.18 3.512 71.39 3.738 ;
      RECT 71.18 3.522 71.395 3.735 ;
      RECT 71.18 3.59 71.4 3.731 ;
      RECT 71.17 3.595 71.4 3.73 ;
      RECT 71.17 3.687 71.405 3.727 ;
      RECT 71.155 3.22 71.415 3.48 ;
      RECT 70.385 2.21 70.43 3.745 ;
      RECT 70.585 2.21 70.615 2.425 ;
      RECT 68.96 1.95 69.08 2.16 ;
      RECT 68.62 1.9 68.88 2.16 ;
      RECT 68.62 1.945 68.915 2.15 ;
      RECT 70.625 2.226 70.63 2.28 ;
      RECT 70.62 2.219 70.625 2.413 ;
      RECT 70.615 2.213 70.62 2.42 ;
      RECT 70.57 2.21 70.585 2.433 ;
      RECT 70.565 2.21 70.57 2.455 ;
      RECT 70.56 2.21 70.565 2.503 ;
      RECT 70.555 2.21 70.56 2.523 ;
      RECT 70.545 2.21 70.555 2.63 ;
      RECT 70.54 2.21 70.545 2.693 ;
      RECT 70.535 2.21 70.54 2.75 ;
      RECT 70.53 2.21 70.535 2.758 ;
      RECT 70.515 2.21 70.53 2.865 ;
      RECT 70.505 2.21 70.515 3 ;
      RECT 70.495 2.21 70.505 3.11 ;
      RECT 70.485 2.21 70.495 3.167 ;
      RECT 70.48 2.21 70.485 3.207 ;
      RECT 70.475 2.21 70.48 3.243 ;
      RECT 70.465 2.21 70.475 3.283 ;
      RECT 70.46 2.21 70.465 3.325 ;
      RECT 70.44 2.21 70.46 3.39 ;
      RECT 70.445 3.535 70.45 3.715 ;
      RECT 70.44 3.517 70.445 3.723 ;
      RECT 70.435 2.21 70.44 3.453 ;
      RECT 70.435 3.497 70.44 3.73 ;
      RECT 70.43 2.21 70.435 3.74 ;
      RECT 70.375 2.21 70.385 2.51 ;
      RECT 70.38 2.757 70.385 3.745 ;
      RECT 70.375 2.822 70.38 3.745 ;
      RECT 70.37 2.211 70.375 2.5 ;
      RECT 70.365 2.887 70.375 3.745 ;
      RECT 70.36 2.212 70.37 2.49 ;
      RECT 70.35 3 70.365 3.745 ;
      RECT 70.355 2.213 70.36 2.48 ;
      RECT 70.335 2.214 70.355 2.458 ;
      RECT 70.34 3.097 70.35 3.745 ;
      RECT 70.335 3.172 70.34 3.745 ;
      RECT 70.325 2.213 70.335 2.435 ;
      RECT 70.33 3.215 70.335 3.745 ;
      RECT 70.325 3.242 70.33 3.745 ;
      RECT 70.315 2.211 70.325 2.423 ;
      RECT 70.32 3.285 70.325 3.745 ;
      RECT 70.315 3.312 70.32 3.745 ;
      RECT 70.305 2.21 70.315 2.41 ;
      RECT 70.31 3.327 70.315 3.745 ;
      RECT 70.27 3.385 70.31 3.745 ;
      RECT 70.3 2.209 70.305 2.395 ;
      RECT 70.295 2.207 70.3 2.388 ;
      RECT 70.285 2.204 70.295 2.378 ;
      RECT 70.28 2.201 70.285 2.363 ;
      RECT 70.265 2.197 70.28 2.356 ;
      RECT 70.26 3.44 70.27 3.745 ;
      RECT 70.26 2.194 70.265 2.351 ;
      RECT 70.245 2.19 70.26 2.345 ;
      RECT 70.255 3.457 70.26 3.745 ;
      RECT 70.245 3.52 70.255 3.745 ;
      RECT 70.165 2.175 70.245 2.325 ;
      RECT 70.24 3.527 70.245 3.74 ;
      RECT 70.235 3.535 70.24 3.73 ;
      RECT 70.155 2.161 70.165 2.309 ;
      RECT 70.14 2.157 70.155 2.307 ;
      RECT 70.13 2.152 70.14 2.303 ;
      RECT 70.105 2.145 70.13 2.295 ;
      RECT 70.1 2.14 70.105 2.29 ;
      RECT 70.09 2.14 70.1 2.288 ;
      RECT 70.08 2.138 70.09 2.286 ;
      RECT 70.05 2.13 70.08 2.28 ;
      RECT 70.035 2.122 70.05 2.273 ;
      RECT 70.015 2.117 70.035 2.266 ;
      RECT 70.01 2.113 70.015 2.261 ;
      RECT 69.98 2.106 70.01 2.255 ;
      RECT 69.955 2.097 69.98 2.245 ;
      RECT 69.925 2.09 69.955 2.237 ;
      RECT 69.9 2.08 69.925 2.228 ;
      RECT 69.885 2.072 69.9 2.222 ;
      RECT 69.86 2.067 69.885 2.217 ;
      RECT 69.85 2.063 69.86 2.212 ;
      RECT 69.83 2.058 69.85 2.207 ;
      RECT 69.795 2.053 69.83 2.2 ;
      RECT 69.735 2.048 69.795 2.193 ;
      RECT 69.722 2.044 69.735 2.191 ;
      RECT 69.636 2.039 69.722 2.188 ;
      RECT 69.55 2.029 69.636 2.184 ;
      RECT 69.509 2.022 69.55 2.181 ;
      RECT 69.423 2.015 69.509 2.178 ;
      RECT 69.337 2.005 69.423 2.174 ;
      RECT 69.251 1.995 69.337 2.169 ;
      RECT 69.165 1.985 69.251 2.165 ;
      RECT 69.155 1.97 69.165 2.163 ;
      RECT 69.145 1.955 69.155 2.163 ;
      RECT 69.08 1.95 69.145 2.162 ;
      RECT 68.915 1.947 68.96 2.155 ;
      RECT 70.16 2.852 70.165 3.043 ;
      RECT 70.155 2.847 70.16 3.05 ;
      RECT 70.141 2.845 70.155 3.056 ;
      RECT 70.055 2.845 70.141 3.058 ;
      RECT 70.051 2.845 70.055 3.061 ;
      RECT 69.965 2.845 70.051 3.079 ;
      RECT 69.955 2.85 69.965 3.098 ;
      RECT 69.945 2.905 69.955 3.102 ;
      RECT 69.92 2.92 69.945 3.109 ;
      RECT 69.88 2.94 69.92 3.122 ;
      RECT 69.875 2.952 69.88 3.132 ;
      RECT 69.86 2.958 69.875 3.137 ;
      RECT 69.855 2.963 69.86 3.141 ;
      RECT 69.835 2.97 69.855 3.146 ;
      RECT 69.765 2.995 69.835 3.163 ;
      RECT 69.725 3.023 69.765 3.183 ;
      RECT 69.72 3.033 69.725 3.191 ;
      RECT 69.7 3.04 69.72 3.193 ;
      RECT 69.695 3.047 69.7 3.196 ;
      RECT 69.665 3.055 69.695 3.199 ;
      RECT 69.66 3.06 69.665 3.203 ;
      RECT 69.586 3.064 69.66 3.211 ;
      RECT 69.5 3.073 69.586 3.227 ;
      RECT 69.496 3.078 69.5 3.236 ;
      RECT 69.41 3.083 69.496 3.246 ;
      RECT 69.37 3.091 69.41 3.258 ;
      RECT 69.32 3.097 69.37 3.265 ;
      RECT 69.235 3.106 69.32 3.28 ;
      RECT 69.16 3.117 69.235 3.298 ;
      RECT 69.125 3.124 69.16 3.308 ;
      RECT 69.05 3.132 69.125 3.313 ;
      RECT 68.995 3.141 69.05 3.313 ;
      RECT 68.97 3.146 68.995 3.311 ;
      RECT 68.96 3.149 68.97 3.309 ;
      RECT 68.925 3.151 68.96 3.307 ;
      RECT 68.895 3.153 68.925 3.303 ;
      RECT 68.85 3.152 68.895 3.299 ;
      RECT 68.83 3.147 68.85 3.296 ;
      RECT 68.78 3.132 68.83 3.293 ;
      RECT 68.77 3.117 68.78 3.288 ;
      RECT 68.72 3.102 68.77 3.278 ;
      RECT 68.67 3.077 68.72 3.258 ;
      RECT 68.66 3.062 68.67 3.24 ;
      RECT 68.655 3.06 68.66 3.234 ;
      RECT 68.635 3.055 68.655 3.229 ;
      RECT 68.63 3.047 68.635 3.223 ;
      RECT 68.615 3.041 68.63 3.216 ;
      RECT 68.61 3.036 68.615 3.208 ;
      RECT 68.59 3.031 68.61 3.2 ;
      RECT 68.575 3.024 68.59 3.193 ;
      RECT 68.56 3.018 68.575 3.184 ;
      RECT 68.555 3.012 68.56 3.177 ;
      RECT 68.51 2.987 68.555 3.163 ;
      RECT 68.495 2.957 68.51 3.145 ;
      RECT 68.48 2.94 68.495 3.136 ;
      RECT 68.455 2.92 68.48 3.124 ;
      RECT 68.415 2.89 68.455 3.104 ;
      RECT 68.405 2.86 68.415 3.089 ;
      RECT 68.39 2.85 68.405 3.082 ;
      RECT 68.335 2.815 68.39 3.061 ;
      RECT 68.32 2.778 68.335 3.04 ;
      RECT 68.31 2.765 68.32 3.032 ;
      RECT 68.26 2.735 68.31 3.014 ;
      RECT 68.245 2.665 68.26 2.995 ;
      RECT 68.2 2.665 68.245 2.978 ;
      RECT 68.175 2.665 68.2 2.96 ;
      RECT 68.165 2.665 68.175 2.953 ;
      RECT 68.086 2.665 68.165 2.946 ;
      RECT 68 2.665 68.086 2.938 ;
      RECT 67.985 2.697 68 2.933 ;
      RECT 67.91 2.707 67.985 2.929 ;
      RECT 67.89 2.717 67.91 2.924 ;
      RECT 67.865 2.717 67.89 2.921 ;
      RECT 67.855 2.707 67.865 2.92 ;
      RECT 67.845 2.68 67.855 2.919 ;
      RECT 67.805 2.675 67.845 2.917 ;
      RECT 67.76 2.675 67.805 2.913 ;
      RECT 67.735 2.675 67.76 2.908 ;
      RECT 67.685 2.675 67.735 2.895 ;
      RECT 67.645 2.68 67.655 2.88 ;
      RECT 67.655 2.675 67.685 2.885 ;
      RECT 69.64 2.455 69.9 2.715 ;
      RECT 69.635 2.477 69.9 2.673 ;
      RECT 68.875 2.305 69.095 2.67 ;
      RECT 68.857 2.392 69.095 2.669 ;
      RECT 68.84 2.397 69.095 2.666 ;
      RECT 68.84 2.397 69.115 2.665 ;
      RECT 68.81 2.407 69.115 2.663 ;
      RECT 68.805 2.422 69.115 2.659 ;
      RECT 68.805 2.422 69.12 2.658 ;
      RECT 68.8 2.48 69.12 2.656 ;
      RECT 68.8 2.48 69.13 2.653 ;
      RECT 68.795 2.545 69.13 2.648 ;
      RECT 68.875 2.305 69.135 2.565 ;
      RECT 67.62 2.135 67.88 2.395 ;
      RECT 67.62 2.178 67.966 2.369 ;
      RECT 67.62 2.178 68.01 2.368 ;
      RECT 67.62 2.178 68.03 2.366 ;
      RECT 67.62 2.178 68.13 2.365 ;
      RECT 67.62 2.178 68.15 2.363 ;
      RECT 67.62 2.178 68.16 2.358 ;
      RECT 68.03 2.145 68.22 2.355 ;
      RECT 68.03 2.147 68.225 2.353 ;
      RECT 68.02 2.152 68.23 2.345 ;
      RECT 67.966 2.176 68.23 2.345 ;
      RECT 68.01 2.17 68.02 2.367 ;
      RECT 68.02 2.15 68.225 2.353 ;
      RECT 66.975 3.21 67.18 3.44 ;
      RECT 66.915 3.16 66.97 3.42 ;
      RECT 66.975 3.16 67.175 3.44 ;
      RECT 67.945 3.475 67.95 3.502 ;
      RECT 67.935 3.385 67.945 3.507 ;
      RECT 67.93 3.307 67.935 3.513 ;
      RECT 67.92 3.297 67.93 3.52 ;
      RECT 67.915 3.287 67.92 3.526 ;
      RECT 67.905 3.282 67.915 3.528 ;
      RECT 67.89 3.274 67.905 3.536 ;
      RECT 67.875 3.265 67.89 3.548 ;
      RECT 67.865 3.257 67.875 3.558 ;
      RECT 67.83 3.175 67.865 3.576 ;
      RECT 67.795 3.175 67.83 3.595 ;
      RECT 67.78 3.175 67.795 3.603 ;
      RECT 67.725 3.175 67.78 3.603 ;
      RECT 67.691 3.175 67.725 3.594 ;
      RECT 67.605 3.175 67.691 3.57 ;
      RECT 67.595 3.235 67.605 3.552 ;
      RECT 67.555 3.237 67.595 3.543 ;
      RECT 67.55 3.239 67.555 3.533 ;
      RECT 67.53 3.241 67.55 3.528 ;
      RECT 67.52 3.244 67.53 3.523 ;
      RECT 67.51 3.245 67.52 3.518 ;
      RECT 67.486 3.246 67.51 3.51 ;
      RECT 67.4 3.251 67.486 3.488 ;
      RECT 67.345 3.25 67.4 3.461 ;
      RECT 67.33 3.243 67.345 3.448 ;
      RECT 67.295 3.238 67.33 3.444 ;
      RECT 67.24 3.23 67.295 3.443 ;
      RECT 67.18 3.217 67.24 3.441 ;
      RECT 66.97 3.16 66.975 3.428 ;
      RECT 67.045 2.53 67.23 2.74 ;
      RECT 67.035 2.535 67.245 2.733 ;
      RECT 67.075 2.44 67.335 2.7 ;
      RECT 67.03 2.597 67.335 2.623 ;
      RECT 66.375 2.39 66.38 3.19 ;
      RECT 66.32 2.44 66.35 3.19 ;
      RECT 66.31 2.44 66.315 2.75 ;
      RECT 66.295 2.44 66.3 2.745 ;
      RECT 65.84 2.485 65.855 2.7 ;
      RECT 65.77 2.485 65.855 2.695 ;
      RECT 67.035 2.065 67.105 2.275 ;
      RECT 67.105 2.072 67.115 2.27 ;
      RECT 67.001 2.065 67.035 2.282 ;
      RECT 66.915 2.065 67.001 2.306 ;
      RECT 66.905 2.07 66.915 2.325 ;
      RECT 66.9 2.082 66.905 2.328 ;
      RECT 66.885 2.097 66.9 2.332 ;
      RECT 66.88 2.115 66.885 2.336 ;
      RECT 66.84 2.125 66.88 2.345 ;
      RECT 66.825 2.132 66.84 2.357 ;
      RECT 66.81 2.137 66.825 2.362 ;
      RECT 66.795 2.14 66.81 2.367 ;
      RECT 66.785 2.142 66.795 2.371 ;
      RECT 66.75 2.149 66.785 2.379 ;
      RECT 66.715 2.157 66.75 2.393 ;
      RECT 66.705 2.163 66.715 2.402 ;
      RECT 66.7 2.165 66.705 2.404 ;
      RECT 66.68 2.168 66.7 2.41 ;
      RECT 66.65 2.175 66.68 2.421 ;
      RECT 66.64 2.181 66.65 2.428 ;
      RECT 66.615 2.184 66.64 2.435 ;
      RECT 66.605 2.188 66.615 2.443 ;
      RECT 66.6 2.189 66.605 2.465 ;
      RECT 66.595 2.19 66.6 2.48 ;
      RECT 66.59 2.191 66.595 2.495 ;
      RECT 66.585 2.192 66.59 2.51 ;
      RECT 66.58 2.193 66.585 2.54 ;
      RECT 66.57 2.195 66.58 2.573 ;
      RECT 66.555 2.199 66.57 2.62 ;
      RECT 66.545 2.202 66.555 2.665 ;
      RECT 66.54 2.205 66.545 2.693 ;
      RECT 66.53 2.207 66.54 2.72 ;
      RECT 66.525 2.21 66.53 2.755 ;
      RECT 66.495 2.215 66.525 2.813 ;
      RECT 66.49 2.22 66.495 2.898 ;
      RECT 66.485 2.222 66.49 2.933 ;
      RECT 66.48 2.224 66.485 3.015 ;
      RECT 66.475 2.226 66.48 3.103 ;
      RECT 66.465 2.228 66.475 3.185 ;
      RECT 66.45 2.242 66.465 3.19 ;
      RECT 66.415 2.287 66.45 3.19 ;
      RECT 66.405 2.327 66.415 3.19 ;
      RECT 66.39 2.355 66.405 3.19 ;
      RECT 66.385 2.372 66.39 3.19 ;
      RECT 66.38 2.38 66.385 3.19 ;
      RECT 66.37 2.395 66.375 3.19 ;
      RECT 66.365 2.402 66.37 3.19 ;
      RECT 66.355 2.422 66.365 3.19 ;
      RECT 66.35 2.435 66.355 3.19 ;
      RECT 66.315 2.44 66.32 2.775 ;
      RECT 66.3 2.83 66.32 3.19 ;
      RECT 66.3 2.44 66.31 2.748 ;
      RECT 66.295 2.87 66.3 3.19 ;
      RECT 66.245 2.44 66.295 2.743 ;
      RECT 66.29 2.907 66.295 3.19 ;
      RECT 66.28 2.93 66.29 3.19 ;
      RECT 66.275 2.975 66.28 3.19 ;
      RECT 66.265 2.985 66.275 3.183 ;
      RECT 66.191 2.44 66.245 2.737 ;
      RECT 66.105 2.44 66.191 2.73 ;
      RECT 66.056 2.487 66.105 2.723 ;
      RECT 65.97 2.495 66.056 2.716 ;
      RECT 65.955 2.492 65.97 2.711 ;
      RECT 65.941 2.485 65.955 2.71 ;
      RECT 65.855 2.485 65.941 2.705 ;
      RECT 65.76 2.49 65.77 2.69 ;
      RECT 65.35 1.92 65.365 2.32 ;
      RECT 65.545 1.92 65.55 2.18 ;
      RECT 65.29 1.92 65.335 2.18 ;
      RECT 65.745 3.225 65.75 3.43 ;
      RECT 65.74 3.215 65.745 3.435 ;
      RECT 65.735 3.202 65.74 3.44 ;
      RECT 65.73 3.182 65.735 3.44 ;
      RECT 65.705 3.135 65.73 3.44 ;
      RECT 65.67 3.05 65.705 3.44 ;
      RECT 65.665 2.987 65.67 3.44 ;
      RECT 65.66 2.972 65.665 3.44 ;
      RECT 65.645 2.932 65.66 3.44 ;
      RECT 65.64 2.907 65.645 3.44 ;
      RECT 65.63 2.89 65.64 3.44 ;
      RECT 65.595 2.812 65.63 3.44 ;
      RECT 65.59 2.755 65.595 3.44 ;
      RECT 65.585 2.742 65.59 3.44 ;
      RECT 65.575 2.72 65.585 3.44 ;
      RECT 65.565 2.685 65.575 3.44 ;
      RECT 65.555 2.655 65.565 3.44 ;
      RECT 65.545 2.57 65.555 3.083 ;
      RECT 65.552 3.215 65.555 3.44 ;
      RECT 65.55 3.225 65.552 3.44 ;
      RECT 65.54 3.235 65.55 3.435 ;
      RECT 65.535 1.92 65.545 2.315 ;
      RECT 65.54 2.447 65.545 3.058 ;
      RECT 65.535 2.345 65.54 3.041 ;
      RECT 65.525 1.92 65.535 3.017 ;
      RECT 65.52 1.92 65.525 2.988 ;
      RECT 65.515 1.92 65.52 2.978 ;
      RECT 65.495 1.92 65.515 2.94 ;
      RECT 65.49 1.92 65.495 2.898 ;
      RECT 65.485 1.92 65.49 2.878 ;
      RECT 65.455 1.92 65.485 2.828 ;
      RECT 65.445 1.92 65.455 2.775 ;
      RECT 65.44 1.92 65.445 2.748 ;
      RECT 65.435 1.92 65.44 2.733 ;
      RECT 65.425 1.92 65.435 2.71 ;
      RECT 65.415 1.92 65.425 2.685 ;
      RECT 65.41 1.92 65.415 2.625 ;
      RECT 65.4 1.92 65.41 2.563 ;
      RECT 65.395 1.92 65.4 2.483 ;
      RECT 65.39 1.92 65.395 2.448 ;
      RECT 65.385 1.92 65.39 2.423 ;
      RECT 65.38 1.92 65.385 2.408 ;
      RECT 65.375 1.92 65.38 2.378 ;
      RECT 65.37 1.92 65.375 2.355 ;
      RECT 65.365 1.92 65.37 2.328 ;
      RECT 65.335 1.92 65.35 2.315 ;
      RECT 64.49 3.455 64.675 3.665 ;
      RECT 64.48 3.46 64.69 3.658 ;
      RECT 64.48 3.46 64.71 3.63 ;
      RECT 64.48 3.46 64.725 3.609 ;
      RECT 64.48 3.46 64.74 3.607 ;
      RECT 64.48 3.46 64.75 3.606 ;
      RECT 64.48 3.46 64.78 3.603 ;
      RECT 65.13 3.305 65.39 3.565 ;
      RECT 65.09 3.352 65.39 3.548 ;
      RECT 65.081 3.36 65.09 3.551 ;
      RECT 64.675 3.453 65.39 3.548 ;
      RECT 64.995 3.378 65.081 3.558 ;
      RECT 64.69 3.45 65.39 3.548 ;
      RECT 64.936 3.4 64.995 3.57 ;
      RECT 64.71 3.446 65.39 3.548 ;
      RECT 64.85 3.412 64.936 3.581 ;
      RECT 64.725 3.442 65.39 3.548 ;
      RECT 64.795 3.425 64.85 3.593 ;
      RECT 64.74 3.44 65.39 3.548 ;
      RECT 64.78 3.431 64.795 3.599 ;
      RECT 64.75 3.436 65.39 3.548 ;
      RECT 64.895 2.96 65.155 3.22 ;
      RECT 64.895 2.98 65.265 3.19 ;
      RECT 64.895 2.985 65.275 3.185 ;
      RECT 65.086 2.399 65.165 2.63 ;
      RECT 65 2.402 65.215 2.625 ;
      RECT 64.995 2.402 65.215 2.62 ;
      RECT 64.995 2.407 65.225 2.618 ;
      RECT 64.97 2.407 65.225 2.615 ;
      RECT 64.97 2.415 65.235 2.613 ;
      RECT 64.85 2.35 65.11 2.61 ;
      RECT 64.85 2.397 65.16 2.61 ;
      RECT 64.105 2.97 64.11 3.23 ;
      RECT 63.935 2.74 63.94 3.23 ;
      RECT 63.82 2.98 63.825 3.205 ;
      RECT 64.53 2.075 64.535 2.285 ;
      RECT 64.535 2.08 64.55 2.28 ;
      RECT 64.47 2.075 64.53 2.293 ;
      RECT 64.455 2.075 64.47 2.303 ;
      RECT 64.405 2.075 64.455 2.32 ;
      RECT 64.385 2.075 64.405 2.343 ;
      RECT 64.37 2.075 64.385 2.355 ;
      RECT 64.35 2.075 64.37 2.365 ;
      RECT 64.34 2.08 64.35 2.374 ;
      RECT 64.335 2.09 64.34 2.379 ;
      RECT 64.33 2.102 64.335 2.383 ;
      RECT 64.32 2.125 64.33 2.388 ;
      RECT 64.315 2.14 64.32 2.392 ;
      RECT 64.31 2.157 64.315 2.395 ;
      RECT 64.305 2.165 64.31 2.398 ;
      RECT 64.295 2.17 64.305 2.402 ;
      RECT 64.29 2.177 64.295 2.407 ;
      RECT 64.28 2.182 64.29 2.411 ;
      RECT 64.255 2.194 64.28 2.422 ;
      RECT 64.235 2.211 64.255 2.438 ;
      RECT 64.21 2.228 64.235 2.46 ;
      RECT 64.175 2.251 64.21 2.518 ;
      RECT 64.155 2.273 64.175 2.58 ;
      RECT 64.15 2.283 64.155 2.615 ;
      RECT 64.14 2.29 64.15 2.653 ;
      RECT 64.135 2.297 64.14 2.673 ;
      RECT 64.13 2.308 64.135 2.71 ;
      RECT 64.125 2.316 64.13 2.775 ;
      RECT 64.115 2.327 64.125 2.828 ;
      RECT 64.11 2.345 64.115 2.898 ;
      RECT 64.105 2.355 64.11 2.935 ;
      RECT 64.1 2.365 64.105 3.23 ;
      RECT 64.095 2.377 64.1 3.23 ;
      RECT 64.09 2.387 64.095 3.23 ;
      RECT 64.08 2.397 64.09 3.23 ;
      RECT 64.07 2.42 64.08 3.23 ;
      RECT 64.055 2.455 64.07 3.23 ;
      RECT 64.015 2.517 64.055 3.23 ;
      RECT 64.01 2.57 64.015 3.23 ;
      RECT 63.985 2.605 64.01 3.23 ;
      RECT 63.97 2.65 63.985 3.23 ;
      RECT 63.965 2.672 63.97 3.23 ;
      RECT 63.955 2.685 63.965 3.23 ;
      RECT 63.945 2.71 63.955 3.23 ;
      RECT 63.94 2.732 63.945 3.23 ;
      RECT 63.915 2.77 63.935 3.23 ;
      RECT 63.875 2.827 63.915 3.23 ;
      RECT 63.87 2.877 63.875 3.23 ;
      RECT 63.865 2.895 63.87 3.23 ;
      RECT 63.86 2.907 63.865 3.23 ;
      RECT 63.85 2.925 63.86 3.23 ;
      RECT 63.84 2.945 63.85 3.205 ;
      RECT 63.835 2.962 63.84 3.205 ;
      RECT 63.825 2.975 63.835 3.205 ;
      RECT 63.795 2.985 63.82 3.205 ;
      RECT 63.785 2.992 63.795 3.205 ;
      RECT 63.77 3.002 63.785 3.2 ;
      RECT 62.8 2.365 63.09 2.595 ;
      RECT 62.86 0.885 63.03 2.595 ;
      RECT 62.83 0.885 63.18 1.235 ;
      RECT 62.8 0.885 63.18 1.115 ;
      RECT 62.8 7.765 63.09 7.995 ;
      RECT 62.86 6.285 63.03 7.995 ;
      RECT 62.8 6.285 63.09 6.515 ;
      RECT 62.39 2.735 62.72 2.965 ;
      RECT 62.39 2.765 62.89 2.935 ;
      RECT 62.39 2.395 62.58 2.965 ;
      RECT 61.81 2.365 62.1 2.595 ;
      RECT 61.81 2.395 62.58 2.565 ;
      RECT 61.87 0.885 62.04 2.595 ;
      RECT 61.81 0.885 62.1 1.115 ;
      RECT 61.81 7.765 62.1 7.995 ;
      RECT 61.87 6.285 62.04 7.995 ;
      RECT 61.81 6.285 62.1 6.515 ;
      RECT 61.81 6.325 62.66 6.485 ;
      RECT 62.49 5.915 62.66 6.485 ;
      RECT 61.81 6.32 62.2 6.485 ;
      RECT 62.43 5.915 62.72 6.145 ;
      RECT 62.43 5.945 62.89 6.115 ;
      RECT 61.44 2.735 61.73 2.965 ;
      RECT 61.44 2.765 61.9 2.935 ;
      RECT 61.5 1.655 61.665 2.965 ;
      RECT 60.015 1.625 60.305 1.855 ;
      RECT 60.015 1.655 61.665 1.825 ;
      RECT 60.075 0.885 60.245 1.855 ;
      RECT 60.015 0.885 60.305 1.115 ;
      RECT 60.015 7.765 60.305 7.995 ;
      RECT 60.075 7.025 60.245 7.995 ;
      RECT 60.075 7.12 61.665 7.29 ;
      RECT 61.495 5.915 61.665 7.29 ;
      RECT 60.015 7.025 60.305 7.255 ;
      RECT 61.44 5.915 61.73 6.145 ;
      RECT 61.44 5.945 61.9 6.115 ;
      RECT 60.445 1.965 60.795 2.315 ;
      RECT 60.275 2.025 60.795 2.195 ;
      RECT 60.47 6.655 60.795 6.98 ;
      RECT 60.445 6.655 60.795 6.885 ;
      RECT 60.275 6.685 60.795 6.855 ;
      RECT 59.67 2.365 59.99 2.685 ;
      RECT 59.64 2.365 59.99 2.595 ;
      RECT 58.11 2.395 59.99 2.565 ;
      RECT 58.11 1.34 58.28 2.565 ;
      RECT 58.01 1.34 58.36 1.69 ;
      RECT 59.67 6.28 59.99 6.605 ;
      RECT 59.64 6.285 59.99 6.515 ;
      RECT 59.47 6.315 59.99 6.485 ;
      RECT 58.615 2.705 58.965 3.055 ;
      RECT 58.615 2.765 59.105 2.935 ;
      RECT 58.62 5.855 58.97 6.205 ;
      RECT 58.62 5.945 59.105 6.115 ;
      RECT 56.305 2.465 56.49 2.675 ;
      RECT 56.295 2.47 56.505 2.668 ;
      RECT 56.295 2.47 56.591 2.645 ;
      RECT 56.295 2.47 56.65 2.62 ;
      RECT 56.295 2.47 56.705 2.6 ;
      RECT 56.295 2.47 56.715 2.588 ;
      RECT 56.295 2.47 56.91 2.527 ;
      RECT 56.295 2.47 56.94 2.51 ;
      RECT 56.295 2.47 56.96 2.5 ;
      RECT 56.84 2.235 57.1 2.495 ;
      RECT 56.825 2.325 56.84 2.542 ;
      RECT 56.36 2.457 57.1 2.495 ;
      RECT 56.811 2.336 56.825 2.548 ;
      RECT 56.4 2.45 57.1 2.495 ;
      RECT 56.725 2.376 56.811 2.567 ;
      RECT 56.65 2.437 57.1 2.495 ;
      RECT 56.72 2.412 56.725 2.584 ;
      RECT 56.705 2.422 57.1 2.495 ;
      RECT 56.715 2.417 56.72 2.586 ;
      RECT 57.01 2.922 57.015 3.014 ;
      RECT 57.005 2.9 57.01 3.031 ;
      RECT 57 2.89 57.005 3.043 ;
      RECT 56.99 2.881 57 3.053 ;
      RECT 56.985 2.876 56.99 3.061 ;
      RECT 56.98 2.735 56.985 3.064 ;
      RECT 56.946 2.735 56.98 3.075 ;
      RECT 56.86 2.735 56.946 3.11 ;
      RECT 56.78 2.735 56.86 3.158 ;
      RECT 56.751 2.735 56.78 3.182 ;
      RECT 56.665 2.735 56.751 3.188 ;
      RECT 56.66 2.919 56.665 3.193 ;
      RECT 56.625 2.93 56.66 3.196 ;
      RECT 56.6 2.945 56.625 3.2 ;
      RECT 56.586 2.954 56.6 3.202 ;
      RECT 56.5 2.981 56.586 3.208 ;
      RECT 56.435 3.022 56.5 3.217 ;
      RECT 56.42 3.042 56.435 3.222 ;
      RECT 56.39 3.052 56.42 3.225 ;
      RECT 56.385 3.062 56.39 3.228 ;
      RECT 56.355 3.067 56.385 3.23 ;
      RECT 56.335 3.072 56.355 3.234 ;
      RECT 56.25 3.075 56.335 3.241 ;
      RECT 56.235 3.072 56.25 3.247 ;
      RECT 56.225 3.069 56.235 3.249 ;
      RECT 56.205 3.066 56.225 3.251 ;
      RECT 56.185 3.062 56.205 3.252 ;
      RECT 56.17 3.058 56.185 3.254 ;
      RECT 56.16 3.055 56.17 3.255 ;
      RECT 56.12 3.049 56.16 3.253 ;
      RECT 56.11 3.044 56.12 3.251 ;
      RECT 56.095 3.041 56.11 3.247 ;
      RECT 56.07 3.036 56.095 3.24 ;
      RECT 56.02 3.027 56.07 3.228 ;
      RECT 55.95 3.013 56.02 3.21 ;
      RECT 55.892 2.998 55.95 3.192 ;
      RECT 55.806 2.981 55.892 3.172 ;
      RECT 55.72 2.96 55.806 3.147 ;
      RECT 55.67 2.945 55.72 3.128 ;
      RECT 55.666 2.939 55.67 3.12 ;
      RECT 55.58 2.929 55.666 3.107 ;
      RECT 55.545 2.914 55.58 3.09 ;
      RECT 55.53 2.907 55.545 3.083 ;
      RECT 55.47 2.895 55.53 3.071 ;
      RECT 55.45 2.882 55.47 3.059 ;
      RECT 55.41 2.873 55.45 3.051 ;
      RECT 55.405 2.865 55.41 3.044 ;
      RECT 55.325 2.855 55.405 3.03 ;
      RECT 55.31 2.842 55.325 3.015 ;
      RECT 55.305 2.84 55.31 3.013 ;
      RECT 55.226 2.828 55.305 3 ;
      RECT 55.14 2.803 55.226 2.975 ;
      RECT 55.125 2.772 55.14 2.96 ;
      RECT 55.11 2.747 55.125 2.956 ;
      RECT 55.095 2.74 55.11 2.952 ;
      RECT 54.92 2.745 54.925 2.948 ;
      RECT 54.915 2.75 54.92 2.943 ;
      RECT 54.925 2.74 55.095 2.95 ;
      RECT 55.64 2.5 55.745 2.76 ;
      RECT 56.455 2.025 56.46 2.25 ;
      RECT 56.585 2.025 56.64 2.235 ;
      RECT 56.64 2.03 56.65 2.228 ;
      RECT 56.546 2.025 56.585 2.238 ;
      RECT 56.46 2.025 56.546 2.245 ;
      RECT 56.44 2.03 56.455 2.251 ;
      RECT 56.43 2.07 56.44 2.253 ;
      RECT 56.4 2.08 56.43 2.255 ;
      RECT 56.395 2.085 56.4 2.257 ;
      RECT 56.37 2.09 56.395 2.259 ;
      RECT 56.355 2.095 56.37 2.261 ;
      RECT 56.34 2.097 56.355 2.263 ;
      RECT 56.335 2.102 56.34 2.265 ;
      RECT 56.285 2.11 56.335 2.268 ;
      RECT 56.26 2.119 56.285 2.273 ;
      RECT 56.25 2.126 56.26 2.278 ;
      RECT 56.245 2.129 56.25 2.282 ;
      RECT 56.225 2.132 56.245 2.291 ;
      RECT 56.195 2.14 56.225 2.311 ;
      RECT 56.166 2.153 56.195 2.333 ;
      RECT 56.08 2.187 56.166 2.377 ;
      RECT 56.075 2.213 56.08 2.415 ;
      RECT 56.07 2.217 56.075 2.424 ;
      RECT 56.035 2.23 56.07 2.457 ;
      RECT 56.025 2.244 56.035 2.495 ;
      RECT 56.02 2.248 56.025 2.508 ;
      RECT 56.015 2.252 56.02 2.513 ;
      RECT 56.005 2.26 56.015 2.525 ;
      RECT 56 2.267 56.005 2.54 ;
      RECT 55.975 2.28 56 2.565 ;
      RECT 55.935 2.309 55.975 2.62 ;
      RECT 55.92 2.334 55.935 2.675 ;
      RECT 55.91 2.345 55.92 2.698 ;
      RECT 55.905 2.352 55.91 2.71 ;
      RECT 55.9 2.356 55.905 2.718 ;
      RECT 55.845 2.384 55.9 2.76 ;
      RECT 55.825 2.42 55.845 2.76 ;
      RECT 55.81 2.435 55.825 2.76 ;
      RECT 55.755 2.467 55.81 2.76 ;
      RECT 55.745 2.497 55.755 2.76 ;
      RECT 55.355 2.112 55.54 2.35 ;
      RECT 55.34 2.114 55.55 2.345 ;
      RECT 55.225 2.06 55.485 2.32 ;
      RECT 55.22 2.097 55.485 2.274 ;
      RECT 55.215 2.107 55.485 2.271 ;
      RECT 55.21 2.147 55.55 2.265 ;
      RECT 55.205 2.18 55.55 2.255 ;
      RECT 55.215 2.122 55.565 2.193 ;
      RECT 55.512 3.22 55.525 3.75 ;
      RECT 55.426 3.22 55.525 3.749 ;
      RECT 55.426 3.22 55.53 3.748 ;
      RECT 55.34 3.22 55.53 3.746 ;
      RECT 55.335 3.22 55.53 3.743 ;
      RECT 55.335 3.22 55.54 3.741 ;
      RECT 55.33 3.512 55.54 3.738 ;
      RECT 55.33 3.522 55.545 3.735 ;
      RECT 55.33 3.59 55.55 3.731 ;
      RECT 55.32 3.595 55.55 3.73 ;
      RECT 55.32 3.687 55.555 3.727 ;
      RECT 55.305 3.22 55.565 3.48 ;
      RECT 54.535 2.21 54.58 3.745 ;
      RECT 54.735 2.21 54.765 2.425 ;
      RECT 53.11 1.95 53.23 2.16 ;
      RECT 52.77 1.9 53.03 2.16 ;
      RECT 52.77 1.945 53.065 2.15 ;
      RECT 54.775 2.226 54.78 2.28 ;
      RECT 54.77 2.219 54.775 2.413 ;
      RECT 54.765 2.213 54.77 2.42 ;
      RECT 54.72 2.21 54.735 2.433 ;
      RECT 54.715 2.21 54.72 2.455 ;
      RECT 54.71 2.21 54.715 2.503 ;
      RECT 54.705 2.21 54.71 2.523 ;
      RECT 54.695 2.21 54.705 2.63 ;
      RECT 54.69 2.21 54.695 2.693 ;
      RECT 54.685 2.21 54.69 2.75 ;
      RECT 54.68 2.21 54.685 2.758 ;
      RECT 54.665 2.21 54.68 2.865 ;
      RECT 54.655 2.21 54.665 3 ;
      RECT 54.645 2.21 54.655 3.11 ;
      RECT 54.635 2.21 54.645 3.167 ;
      RECT 54.63 2.21 54.635 3.207 ;
      RECT 54.625 2.21 54.63 3.243 ;
      RECT 54.615 2.21 54.625 3.283 ;
      RECT 54.61 2.21 54.615 3.325 ;
      RECT 54.59 2.21 54.61 3.39 ;
      RECT 54.595 3.535 54.6 3.715 ;
      RECT 54.59 3.517 54.595 3.723 ;
      RECT 54.585 2.21 54.59 3.453 ;
      RECT 54.585 3.497 54.59 3.73 ;
      RECT 54.58 2.21 54.585 3.74 ;
      RECT 54.525 2.21 54.535 2.51 ;
      RECT 54.53 2.757 54.535 3.745 ;
      RECT 54.525 2.822 54.53 3.745 ;
      RECT 54.52 2.211 54.525 2.5 ;
      RECT 54.515 2.887 54.525 3.745 ;
      RECT 54.51 2.212 54.52 2.49 ;
      RECT 54.5 3 54.515 3.745 ;
      RECT 54.505 2.213 54.51 2.48 ;
      RECT 54.485 2.214 54.505 2.458 ;
      RECT 54.49 3.097 54.5 3.745 ;
      RECT 54.485 3.172 54.49 3.745 ;
      RECT 54.475 2.213 54.485 2.435 ;
      RECT 54.48 3.215 54.485 3.745 ;
      RECT 54.475 3.242 54.48 3.745 ;
      RECT 54.465 2.211 54.475 2.423 ;
      RECT 54.47 3.285 54.475 3.745 ;
      RECT 54.465 3.312 54.47 3.745 ;
      RECT 54.455 2.21 54.465 2.41 ;
      RECT 54.46 3.327 54.465 3.745 ;
      RECT 54.42 3.385 54.46 3.745 ;
      RECT 54.45 2.209 54.455 2.395 ;
      RECT 54.445 2.207 54.45 2.388 ;
      RECT 54.435 2.204 54.445 2.378 ;
      RECT 54.43 2.201 54.435 2.363 ;
      RECT 54.415 2.197 54.43 2.356 ;
      RECT 54.41 3.44 54.42 3.745 ;
      RECT 54.41 2.194 54.415 2.351 ;
      RECT 54.395 2.19 54.41 2.345 ;
      RECT 54.405 3.457 54.41 3.745 ;
      RECT 54.395 3.52 54.405 3.745 ;
      RECT 54.315 2.175 54.395 2.325 ;
      RECT 54.39 3.527 54.395 3.74 ;
      RECT 54.385 3.535 54.39 3.73 ;
      RECT 54.305 2.161 54.315 2.309 ;
      RECT 54.29 2.157 54.305 2.307 ;
      RECT 54.28 2.152 54.29 2.303 ;
      RECT 54.255 2.145 54.28 2.295 ;
      RECT 54.25 2.14 54.255 2.29 ;
      RECT 54.24 2.14 54.25 2.288 ;
      RECT 54.23 2.138 54.24 2.286 ;
      RECT 54.2 2.13 54.23 2.28 ;
      RECT 54.185 2.122 54.2 2.273 ;
      RECT 54.165 2.117 54.185 2.266 ;
      RECT 54.16 2.113 54.165 2.261 ;
      RECT 54.13 2.106 54.16 2.255 ;
      RECT 54.105 2.097 54.13 2.245 ;
      RECT 54.075 2.09 54.105 2.237 ;
      RECT 54.05 2.08 54.075 2.228 ;
      RECT 54.035 2.072 54.05 2.222 ;
      RECT 54.01 2.067 54.035 2.217 ;
      RECT 54 2.063 54.01 2.212 ;
      RECT 53.98 2.058 54 2.207 ;
      RECT 53.945 2.053 53.98 2.2 ;
      RECT 53.885 2.048 53.945 2.193 ;
      RECT 53.872 2.044 53.885 2.191 ;
      RECT 53.786 2.039 53.872 2.188 ;
      RECT 53.7 2.029 53.786 2.184 ;
      RECT 53.659 2.022 53.7 2.181 ;
      RECT 53.573 2.015 53.659 2.178 ;
      RECT 53.487 2.005 53.573 2.174 ;
      RECT 53.401 1.995 53.487 2.169 ;
      RECT 53.315 1.985 53.401 2.165 ;
      RECT 53.305 1.97 53.315 2.163 ;
      RECT 53.295 1.955 53.305 2.163 ;
      RECT 53.23 1.95 53.295 2.162 ;
      RECT 53.065 1.947 53.11 2.155 ;
      RECT 54.31 2.852 54.315 3.043 ;
      RECT 54.305 2.847 54.31 3.05 ;
      RECT 54.291 2.845 54.305 3.056 ;
      RECT 54.205 2.845 54.291 3.058 ;
      RECT 54.201 2.845 54.205 3.061 ;
      RECT 54.115 2.845 54.201 3.079 ;
      RECT 54.105 2.85 54.115 3.098 ;
      RECT 54.095 2.905 54.105 3.102 ;
      RECT 54.07 2.92 54.095 3.109 ;
      RECT 54.03 2.94 54.07 3.122 ;
      RECT 54.025 2.952 54.03 3.132 ;
      RECT 54.01 2.958 54.025 3.137 ;
      RECT 54.005 2.963 54.01 3.141 ;
      RECT 53.985 2.97 54.005 3.146 ;
      RECT 53.915 2.995 53.985 3.163 ;
      RECT 53.875 3.023 53.915 3.183 ;
      RECT 53.87 3.033 53.875 3.191 ;
      RECT 53.85 3.04 53.87 3.193 ;
      RECT 53.845 3.047 53.85 3.196 ;
      RECT 53.815 3.055 53.845 3.199 ;
      RECT 53.81 3.06 53.815 3.203 ;
      RECT 53.736 3.064 53.81 3.211 ;
      RECT 53.65 3.073 53.736 3.227 ;
      RECT 53.646 3.078 53.65 3.236 ;
      RECT 53.56 3.083 53.646 3.246 ;
      RECT 53.52 3.091 53.56 3.258 ;
      RECT 53.47 3.097 53.52 3.265 ;
      RECT 53.385 3.106 53.47 3.28 ;
      RECT 53.31 3.117 53.385 3.298 ;
      RECT 53.275 3.124 53.31 3.308 ;
      RECT 53.2 3.132 53.275 3.313 ;
      RECT 53.145 3.141 53.2 3.313 ;
      RECT 53.12 3.146 53.145 3.311 ;
      RECT 53.11 3.149 53.12 3.309 ;
      RECT 53.075 3.151 53.11 3.307 ;
      RECT 53.045 3.153 53.075 3.303 ;
      RECT 53 3.152 53.045 3.299 ;
      RECT 52.98 3.147 53 3.296 ;
      RECT 52.93 3.132 52.98 3.293 ;
      RECT 52.92 3.117 52.93 3.288 ;
      RECT 52.87 3.102 52.92 3.278 ;
      RECT 52.82 3.077 52.87 3.258 ;
      RECT 52.81 3.062 52.82 3.24 ;
      RECT 52.805 3.06 52.81 3.234 ;
      RECT 52.785 3.055 52.805 3.229 ;
      RECT 52.78 3.047 52.785 3.223 ;
      RECT 52.765 3.041 52.78 3.216 ;
      RECT 52.76 3.036 52.765 3.208 ;
      RECT 52.74 3.031 52.76 3.2 ;
      RECT 52.725 3.024 52.74 3.193 ;
      RECT 52.71 3.018 52.725 3.184 ;
      RECT 52.705 3.012 52.71 3.177 ;
      RECT 52.66 2.987 52.705 3.163 ;
      RECT 52.645 2.957 52.66 3.145 ;
      RECT 52.63 2.94 52.645 3.136 ;
      RECT 52.605 2.92 52.63 3.124 ;
      RECT 52.565 2.89 52.605 3.104 ;
      RECT 52.555 2.86 52.565 3.089 ;
      RECT 52.54 2.85 52.555 3.082 ;
      RECT 52.485 2.815 52.54 3.061 ;
      RECT 52.47 2.778 52.485 3.04 ;
      RECT 52.46 2.765 52.47 3.032 ;
      RECT 52.41 2.735 52.46 3.014 ;
      RECT 52.395 2.665 52.41 2.995 ;
      RECT 52.35 2.665 52.395 2.978 ;
      RECT 52.325 2.665 52.35 2.96 ;
      RECT 52.315 2.665 52.325 2.953 ;
      RECT 52.236 2.665 52.315 2.946 ;
      RECT 52.15 2.665 52.236 2.938 ;
      RECT 52.135 2.697 52.15 2.933 ;
      RECT 52.06 2.707 52.135 2.929 ;
      RECT 52.04 2.717 52.06 2.924 ;
      RECT 52.015 2.717 52.04 2.921 ;
      RECT 52.005 2.707 52.015 2.92 ;
      RECT 51.995 2.68 52.005 2.919 ;
      RECT 51.955 2.675 51.995 2.917 ;
      RECT 51.91 2.675 51.955 2.913 ;
      RECT 51.885 2.675 51.91 2.908 ;
      RECT 51.835 2.675 51.885 2.895 ;
      RECT 51.795 2.68 51.805 2.88 ;
      RECT 51.805 2.675 51.835 2.885 ;
      RECT 53.79 2.455 54.05 2.715 ;
      RECT 53.785 2.477 54.05 2.673 ;
      RECT 53.025 2.305 53.245 2.67 ;
      RECT 53.007 2.392 53.245 2.669 ;
      RECT 52.99 2.397 53.245 2.666 ;
      RECT 52.99 2.397 53.265 2.665 ;
      RECT 52.96 2.407 53.265 2.663 ;
      RECT 52.955 2.422 53.265 2.659 ;
      RECT 52.955 2.422 53.27 2.658 ;
      RECT 52.95 2.48 53.27 2.656 ;
      RECT 52.95 2.48 53.28 2.653 ;
      RECT 52.945 2.545 53.28 2.648 ;
      RECT 53.025 2.305 53.285 2.565 ;
      RECT 51.77 2.135 52.03 2.395 ;
      RECT 51.77 2.178 52.116 2.369 ;
      RECT 51.77 2.178 52.16 2.368 ;
      RECT 51.77 2.178 52.18 2.366 ;
      RECT 51.77 2.178 52.28 2.365 ;
      RECT 51.77 2.178 52.3 2.363 ;
      RECT 51.77 2.178 52.31 2.358 ;
      RECT 52.18 2.145 52.37 2.355 ;
      RECT 52.18 2.147 52.375 2.353 ;
      RECT 52.17 2.152 52.38 2.345 ;
      RECT 52.116 2.176 52.38 2.345 ;
      RECT 52.16 2.17 52.17 2.367 ;
      RECT 52.17 2.15 52.375 2.353 ;
      RECT 51.125 3.21 51.33 3.44 ;
      RECT 51.065 3.16 51.12 3.42 ;
      RECT 51.125 3.16 51.325 3.44 ;
      RECT 52.095 3.475 52.1 3.502 ;
      RECT 52.085 3.385 52.095 3.507 ;
      RECT 52.08 3.307 52.085 3.513 ;
      RECT 52.07 3.297 52.08 3.52 ;
      RECT 52.065 3.287 52.07 3.526 ;
      RECT 52.055 3.282 52.065 3.528 ;
      RECT 52.04 3.274 52.055 3.536 ;
      RECT 52.025 3.265 52.04 3.548 ;
      RECT 52.015 3.257 52.025 3.558 ;
      RECT 51.98 3.175 52.015 3.576 ;
      RECT 51.945 3.175 51.98 3.595 ;
      RECT 51.93 3.175 51.945 3.603 ;
      RECT 51.875 3.175 51.93 3.603 ;
      RECT 51.841 3.175 51.875 3.594 ;
      RECT 51.755 3.175 51.841 3.57 ;
      RECT 51.745 3.235 51.755 3.552 ;
      RECT 51.705 3.237 51.745 3.543 ;
      RECT 51.7 3.239 51.705 3.533 ;
      RECT 51.68 3.241 51.7 3.528 ;
      RECT 51.67 3.244 51.68 3.523 ;
      RECT 51.66 3.245 51.67 3.518 ;
      RECT 51.636 3.246 51.66 3.51 ;
      RECT 51.55 3.251 51.636 3.488 ;
      RECT 51.495 3.25 51.55 3.461 ;
      RECT 51.48 3.243 51.495 3.448 ;
      RECT 51.445 3.238 51.48 3.444 ;
      RECT 51.39 3.23 51.445 3.443 ;
      RECT 51.33 3.217 51.39 3.441 ;
      RECT 51.12 3.16 51.125 3.428 ;
      RECT 51.195 2.53 51.38 2.74 ;
      RECT 51.185 2.535 51.395 2.733 ;
      RECT 51.225 2.44 51.485 2.7 ;
      RECT 51.18 2.597 51.485 2.623 ;
      RECT 50.525 2.39 50.53 3.19 ;
      RECT 50.47 2.44 50.5 3.19 ;
      RECT 50.46 2.44 50.465 2.75 ;
      RECT 50.445 2.44 50.45 2.745 ;
      RECT 49.99 2.485 50.005 2.7 ;
      RECT 49.92 2.485 50.005 2.695 ;
      RECT 51.185 2.065 51.255 2.275 ;
      RECT 51.255 2.072 51.265 2.27 ;
      RECT 51.151 2.065 51.185 2.282 ;
      RECT 51.065 2.065 51.151 2.306 ;
      RECT 51.055 2.07 51.065 2.325 ;
      RECT 51.05 2.082 51.055 2.328 ;
      RECT 51.035 2.097 51.05 2.332 ;
      RECT 51.03 2.115 51.035 2.336 ;
      RECT 50.99 2.125 51.03 2.345 ;
      RECT 50.975 2.132 50.99 2.357 ;
      RECT 50.96 2.137 50.975 2.362 ;
      RECT 50.945 2.14 50.96 2.367 ;
      RECT 50.935 2.142 50.945 2.371 ;
      RECT 50.9 2.149 50.935 2.379 ;
      RECT 50.865 2.157 50.9 2.393 ;
      RECT 50.855 2.163 50.865 2.402 ;
      RECT 50.85 2.165 50.855 2.404 ;
      RECT 50.83 2.168 50.85 2.41 ;
      RECT 50.8 2.175 50.83 2.421 ;
      RECT 50.79 2.181 50.8 2.428 ;
      RECT 50.765 2.184 50.79 2.435 ;
      RECT 50.755 2.188 50.765 2.443 ;
      RECT 50.75 2.189 50.755 2.465 ;
      RECT 50.745 2.19 50.75 2.48 ;
      RECT 50.74 2.191 50.745 2.495 ;
      RECT 50.735 2.192 50.74 2.51 ;
      RECT 50.73 2.193 50.735 2.54 ;
      RECT 50.72 2.195 50.73 2.573 ;
      RECT 50.705 2.199 50.72 2.62 ;
      RECT 50.695 2.202 50.705 2.665 ;
      RECT 50.69 2.205 50.695 2.693 ;
      RECT 50.68 2.207 50.69 2.72 ;
      RECT 50.675 2.21 50.68 2.755 ;
      RECT 50.645 2.215 50.675 2.813 ;
      RECT 50.64 2.22 50.645 2.898 ;
      RECT 50.635 2.222 50.64 2.933 ;
      RECT 50.63 2.224 50.635 3.015 ;
      RECT 50.625 2.226 50.63 3.103 ;
      RECT 50.615 2.228 50.625 3.185 ;
      RECT 50.6 2.242 50.615 3.19 ;
      RECT 50.565 2.287 50.6 3.19 ;
      RECT 50.555 2.327 50.565 3.19 ;
      RECT 50.54 2.355 50.555 3.19 ;
      RECT 50.535 2.372 50.54 3.19 ;
      RECT 50.53 2.38 50.535 3.19 ;
      RECT 50.52 2.395 50.525 3.19 ;
      RECT 50.515 2.402 50.52 3.19 ;
      RECT 50.505 2.422 50.515 3.19 ;
      RECT 50.5 2.435 50.505 3.19 ;
      RECT 50.465 2.44 50.47 2.775 ;
      RECT 50.45 2.83 50.47 3.19 ;
      RECT 50.45 2.44 50.46 2.748 ;
      RECT 50.445 2.87 50.45 3.19 ;
      RECT 50.395 2.44 50.445 2.743 ;
      RECT 50.44 2.907 50.445 3.19 ;
      RECT 50.43 2.93 50.44 3.19 ;
      RECT 50.425 2.975 50.43 3.19 ;
      RECT 50.415 2.985 50.425 3.183 ;
      RECT 50.341 2.44 50.395 2.737 ;
      RECT 50.255 2.44 50.341 2.73 ;
      RECT 50.206 2.487 50.255 2.723 ;
      RECT 50.12 2.495 50.206 2.716 ;
      RECT 50.105 2.492 50.12 2.711 ;
      RECT 50.091 2.485 50.105 2.71 ;
      RECT 50.005 2.485 50.091 2.705 ;
      RECT 49.91 2.49 49.92 2.69 ;
      RECT 49.5 1.92 49.515 2.32 ;
      RECT 49.695 1.92 49.7 2.18 ;
      RECT 49.44 1.92 49.485 2.18 ;
      RECT 49.895 3.225 49.9 3.43 ;
      RECT 49.89 3.215 49.895 3.435 ;
      RECT 49.885 3.202 49.89 3.44 ;
      RECT 49.88 3.182 49.885 3.44 ;
      RECT 49.855 3.135 49.88 3.44 ;
      RECT 49.82 3.05 49.855 3.44 ;
      RECT 49.815 2.987 49.82 3.44 ;
      RECT 49.81 2.972 49.815 3.44 ;
      RECT 49.795 2.932 49.81 3.44 ;
      RECT 49.79 2.907 49.795 3.44 ;
      RECT 49.78 2.89 49.79 3.44 ;
      RECT 49.745 2.812 49.78 3.44 ;
      RECT 49.74 2.755 49.745 3.44 ;
      RECT 49.735 2.742 49.74 3.44 ;
      RECT 49.725 2.72 49.735 3.44 ;
      RECT 49.715 2.685 49.725 3.44 ;
      RECT 49.705 2.655 49.715 3.44 ;
      RECT 49.695 2.57 49.705 3.083 ;
      RECT 49.702 3.215 49.705 3.44 ;
      RECT 49.7 3.225 49.702 3.44 ;
      RECT 49.69 3.235 49.7 3.435 ;
      RECT 49.685 1.92 49.695 2.315 ;
      RECT 49.69 2.447 49.695 3.058 ;
      RECT 49.685 2.345 49.69 3.041 ;
      RECT 49.675 1.92 49.685 3.017 ;
      RECT 49.67 1.92 49.675 2.988 ;
      RECT 49.665 1.92 49.67 2.978 ;
      RECT 49.645 1.92 49.665 2.94 ;
      RECT 49.64 1.92 49.645 2.898 ;
      RECT 49.635 1.92 49.64 2.878 ;
      RECT 49.605 1.92 49.635 2.828 ;
      RECT 49.595 1.92 49.605 2.775 ;
      RECT 49.59 1.92 49.595 2.748 ;
      RECT 49.585 1.92 49.59 2.733 ;
      RECT 49.575 1.92 49.585 2.71 ;
      RECT 49.565 1.92 49.575 2.685 ;
      RECT 49.56 1.92 49.565 2.625 ;
      RECT 49.55 1.92 49.56 2.563 ;
      RECT 49.545 1.92 49.55 2.483 ;
      RECT 49.54 1.92 49.545 2.448 ;
      RECT 49.535 1.92 49.54 2.423 ;
      RECT 49.53 1.92 49.535 2.408 ;
      RECT 49.525 1.92 49.53 2.378 ;
      RECT 49.52 1.92 49.525 2.355 ;
      RECT 49.515 1.92 49.52 2.328 ;
      RECT 49.485 1.92 49.5 2.315 ;
      RECT 48.64 3.455 48.825 3.665 ;
      RECT 48.63 3.46 48.84 3.658 ;
      RECT 48.63 3.46 48.86 3.63 ;
      RECT 48.63 3.46 48.875 3.609 ;
      RECT 48.63 3.46 48.89 3.607 ;
      RECT 48.63 3.46 48.9 3.606 ;
      RECT 48.63 3.46 48.93 3.603 ;
      RECT 49.28 3.305 49.54 3.565 ;
      RECT 49.24 3.352 49.54 3.548 ;
      RECT 49.231 3.36 49.24 3.551 ;
      RECT 48.825 3.453 49.54 3.548 ;
      RECT 49.145 3.378 49.231 3.558 ;
      RECT 48.84 3.45 49.54 3.548 ;
      RECT 49.086 3.4 49.145 3.57 ;
      RECT 48.86 3.446 49.54 3.548 ;
      RECT 49 3.412 49.086 3.581 ;
      RECT 48.875 3.442 49.54 3.548 ;
      RECT 48.945 3.425 49 3.593 ;
      RECT 48.89 3.44 49.54 3.548 ;
      RECT 48.93 3.431 48.945 3.599 ;
      RECT 48.9 3.436 49.54 3.548 ;
      RECT 49.045 2.96 49.305 3.22 ;
      RECT 49.045 2.98 49.415 3.19 ;
      RECT 49.045 2.985 49.425 3.185 ;
      RECT 49.236 2.399 49.315 2.63 ;
      RECT 49.15 2.402 49.365 2.625 ;
      RECT 49.145 2.402 49.365 2.62 ;
      RECT 49.145 2.407 49.375 2.618 ;
      RECT 49.12 2.407 49.375 2.615 ;
      RECT 49.12 2.415 49.385 2.613 ;
      RECT 49 2.35 49.26 2.61 ;
      RECT 49 2.397 49.31 2.61 ;
      RECT 48.255 2.97 48.26 3.23 ;
      RECT 48.085 2.74 48.09 3.23 ;
      RECT 47.97 2.98 47.975 3.205 ;
      RECT 48.68 2.075 48.685 2.285 ;
      RECT 48.685 2.08 48.7 2.28 ;
      RECT 48.62 2.075 48.68 2.293 ;
      RECT 48.605 2.075 48.62 2.303 ;
      RECT 48.555 2.075 48.605 2.32 ;
      RECT 48.535 2.075 48.555 2.343 ;
      RECT 48.52 2.075 48.535 2.355 ;
      RECT 48.5 2.075 48.52 2.365 ;
      RECT 48.49 2.08 48.5 2.374 ;
      RECT 48.485 2.09 48.49 2.379 ;
      RECT 48.48 2.102 48.485 2.383 ;
      RECT 48.47 2.125 48.48 2.388 ;
      RECT 48.465 2.14 48.47 2.392 ;
      RECT 48.46 2.157 48.465 2.395 ;
      RECT 48.455 2.165 48.46 2.398 ;
      RECT 48.445 2.17 48.455 2.402 ;
      RECT 48.44 2.177 48.445 2.407 ;
      RECT 48.43 2.182 48.44 2.411 ;
      RECT 48.405 2.194 48.43 2.422 ;
      RECT 48.385 2.211 48.405 2.438 ;
      RECT 48.36 2.228 48.385 2.46 ;
      RECT 48.325 2.251 48.36 2.518 ;
      RECT 48.305 2.273 48.325 2.58 ;
      RECT 48.3 2.283 48.305 2.615 ;
      RECT 48.29 2.29 48.3 2.653 ;
      RECT 48.285 2.297 48.29 2.673 ;
      RECT 48.28 2.308 48.285 2.71 ;
      RECT 48.275 2.316 48.28 2.775 ;
      RECT 48.265 2.327 48.275 2.828 ;
      RECT 48.26 2.345 48.265 2.898 ;
      RECT 48.255 2.355 48.26 2.935 ;
      RECT 48.25 2.365 48.255 3.23 ;
      RECT 48.245 2.377 48.25 3.23 ;
      RECT 48.24 2.387 48.245 3.23 ;
      RECT 48.23 2.397 48.24 3.23 ;
      RECT 48.22 2.42 48.23 3.23 ;
      RECT 48.205 2.455 48.22 3.23 ;
      RECT 48.165 2.517 48.205 3.23 ;
      RECT 48.16 2.57 48.165 3.23 ;
      RECT 48.135 2.605 48.16 3.23 ;
      RECT 48.12 2.65 48.135 3.23 ;
      RECT 48.115 2.672 48.12 3.23 ;
      RECT 48.105 2.685 48.115 3.23 ;
      RECT 48.095 2.71 48.105 3.23 ;
      RECT 48.09 2.732 48.095 3.23 ;
      RECT 48.065 2.77 48.085 3.23 ;
      RECT 48.025 2.827 48.065 3.23 ;
      RECT 48.02 2.877 48.025 3.23 ;
      RECT 48.015 2.895 48.02 3.23 ;
      RECT 48.01 2.907 48.015 3.23 ;
      RECT 48 2.925 48.01 3.23 ;
      RECT 47.99 2.945 48 3.205 ;
      RECT 47.985 2.962 47.99 3.205 ;
      RECT 47.975 2.975 47.985 3.205 ;
      RECT 47.945 2.985 47.97 3.205 ;
      RECT 47.935 2.992 47.945 3.205 ;
      RECT 47.92 3.002 47.935 3.2 ;
      RECT 46.95 2.365 47.24 2.595 ;
      RECT 47.01 0.885 47.18 2.595 ;
      RECT 46.98 0.885 47.33 1.235 ;
      RECT 46.95 0.885 47.33 1.115 ;
      RECT 46.95 7.765 47.24 7.995 ;
      RECT 47.01 6.285 47.18 7.995 ;
      RECT 46.95 6.285 47.24 6.515 ;
      RECT 46.54 2.735 46.87 2.965 ;
      RECT 46.54 2.765 47.04 2.935 ;
      RECT 46.54 2.395 46.73 2.965 ;
      RECT 45.96 2.365 46.25 2.595 ;
      RECT 45.96 2.395 46.73 2.565 ;
      RECT 46.02 0.885 46.19 2.595 ;
      RECT 45.96 0.885 46.25 1.115 ;
      RECT 45.96 7.765 46.25 7.995 ;
      RECT 46.02 6.285 46.19 7.995 ;
      RECT 45.96 6.285 46.25 6.515 ;
      RECT 45.96 6.325 46.81 6.485 ;
      RECT 46.64 5.915 46.81 6.485 ;
      RECT 45.96 6.32 46.35 6.485 ;
      RECT 46.58 5.915 46.87 6.145 ;
      RECT 46.58 5.945 47.04 6.115 ;
      RECT 45.59 2.735 45.88 2.965 ;
      RECT 45.59 2.765 46.05 2.935 ;
      RECT 45.65 1.655 45.815 2.965 ;
      RECT 44.165 1.625 44.455 1.855 ;
      RECT 44.165 1.655 45.815 1.825 ;
      RECT 44.225 0.885 44.395 1.855 ;
      RECT 44.165 0.885 44.455 1.115 ;
      RECT 44.165 7.765 44.455 7.995 ;
      RECT 44.225 7.025 44.395 7.995 ;
      RECT 44.225 7.12 45.815 7.29 ;
      RECT 45.645 5.915 45.815 7.29 ;
      RECT 44.165 7.025 44.455 7.255 ;
      RECT 45.59 5.915 45.88 6.145 ;
      RECT 45.59 5.945 46.05 6.115 ;
      RECT 44.595 1.965 44.945 2.315 ;
      RECT 44.425 2.025 44.945 2.195 ;
      RECT 44.62 6.655 44.945 6.98 ;
      RECT 44.595 6.655 44.945 6.885 ;
      RECT 44.425 6.685 44.945 6.855 ;
      RECT 43.82 2.365 44.14 2.685 ;
      RECT 43.79 2.365 44.14 2.595 ;
      RECT 42.26 2.395 44.14 2.565 ;
      RECT 42.26 1.34 42.43 2.565 ;
      RECT 42.16 1.34 42.51 1.69 ;
      RECT 43.82 6.28 44.14 6.605 ;
      RECT 43.79 6.285 44.14 6.515 ;
      RECT 43.62 6.315 44.14 6.485 ;
      RECT 42.765 2.705 43.115 3.055 ;
      RECT 42.765 2.765 43.255 2.935 ;
      RECT 42.77 5.855 43.12 6.205 ;
      RECT 42.77 5.945 43.255 6.115 ;
      RECT 40.455 2.465 40.64 2.675 ;
      RECT 40.445 2.47 40.655 2.668 ;
      RECT 40.445 2.47 40.741 2.645 ;
      RECT 40.445 2.47 40.8 2.62 ;
      RECT 40.445 2.47 40.855 2.6 ;
      RECT 40.445 2.47 40.865 2.588 ;
      RECT 40.445 2.47 41.06 2.527 ;
      RECT 40.445 2.47 41.09 2.51 ;
      RECT 40.445 2.47 41.11 2.5 ;
      RECT 40.99 2.235 41.25 2.495 ;
      RECT 40.975 2.325 40.99 2.542 ;
      RECT 40.51 2.457 41.25 2.495 ;
      RECT 40.961 2.336 40.975 2.548 ;
      RECT 40.55 2.45 41.25 2.495 ;
      RECT 40.875 2.376 40.961 2.567 ;
      RECT 40.8 2.437 41.25 2.495 ;
      RECT 40.87 2.412 40.875 2.584 ;
      RECT 40.855 2.422 41.25 2.495 ;
      RECT 40.865 2.417 40.87 2.586 ;
      RECT 41.16 2.922 41.165 3.014 ;
      RECT 41.155 2.9 41.16 3.031 ;
      RECT 41.15 2.89 41.155 3.043 ;
      RECT 41.14 2.881 41.15 3.053 ;
      RECT 41.135 2.876 41.14 3.061 ;
      RECT 41.13 2.735 41.135 3.064 ;
      RECT 41.096 2.735 41.13 3.075 ;
      RECT 41.01 2.735 41.096 3.11 ;
      RECT 40.93 2.735 41.01 3.158 ;
      RECT 40.901 2.735 40.93 3.182 ;
      RECT 40.815 2.735 40.901 3.188 ;
      RECT 40.81 2.919 40.815 3.193 ;
      RECT 40.775 2.93 40.81 3.196 ;
      RECT 40.75 2.945 40.775 3.2 ;
      RECT 40.736 2.954 40.75 3.202 ;
      RECT 40.65 2.981 40.736 3.208 ;
      RECT 40.585 3.022 40.65 3.217 ;
      RECT 40.57 3.042 40.585 3.222 ;
      RECT 40.54 3.052 40.57 3.225 ;
      RECT 40.535 3.062 40.54 3.228 ;
      RECT 40.505 3.067 40.535 3.23 ;
      RECT 40.485 3.072 40.505 3.234 ;
      RECT 40.4 3.075 40.485 3.241 ;
      RECT 40.385 3.072 40.4 3.247 ;
      RECT 40.375 3.069 40.385 3.249 ;
      RECT 40.355 3.066 40.375 3.251 ;
      RECT 40.335 3.062 40.355 3.252 ;
      RECT 40.32 3.058 40.335 3.254 ;
      RECT 40.31 3.055 40.32 3.255 ;
      RECT 40.27 3.049 40.31 3.253 ;
      RECT 40.26 3.044 40.27 3.251 ;
      RECT 40.245 3.041 40.26 3.247 ;
      RECT 40.22 3.036 40.245 3.24 ;
      RECT 40.17 3.027 40.22 3.228 ;
      RECT 40.1 3.013 40.17 3.21 ;
      RECT 40.042 2.998 40.1 3.192 ;
      RECT 39.956 2.981 40.042 3.172 ;
      RECT 39.87 2.96 39.956 3.147 ;
      RECT 39.82 2.945 39.87 3.128 ;
      RECT 39.816 2.939 39.82 3.12 ;
      RECT 39.73 2.929 39.816 3.107 ;
      RECT 39.695 2.914 39.73 3.09 ;
      RECT 39.68 2.907 39.695 3.083 ;
      RECT 39.62 2.895 39.68 3.071 ;
      RECT 39.6 2.882 39.62 3.059 ;
      RECT 39.56 2.873 39.6 3.051 ;
      RECT 39.555 2.865 39.56 3.044 ;
      RECT 39.475 2.855 39.555 3.03 ;
      RECT 39.46 2.842 39.475 3.015 ;
      RECT 39.455 2.84 39.46 3.013 ;
      RECT 39.376 2.828 39.455 3 ;
      RECT 39.29 2.803 39.376 2.975 ;
      RECT 39.275 2.772 39.29 2.96 ;
      RECT 39.26 2.747 39.275 2.956 ;
      RECT 39.245 2.74 39.26 2.952 ;
      RECT 39.07 2.745 39.075 2.948 ;
      RECT 39.065 2.75 39.07 2.943 ;
      RECT 39.075 2.74 39.245 2.95 ;
      RECT 39.79 2.5 39.895 2.76 ;
      RECT 40.605 2.025 40.61 2.25 ;
      RECT 40.735 2.025 40.79 2.235 ;
      RECT 40.79 2.03 40.8 2.228 ;
      RECT 40.696 2.025 40.735 2.238 ;
      RECT 40.61 2.025 40.696 2.245 ;
      RECT 40.59 2.03 40.605 2.251 ;
      RECT 40.58 2.07 40.59 2.253 ;
      RECT 40.55 2.08 40.58 2.255 ;
      RECT 40.545 2.085 40.55 2.257 ;
      RECT 40.52 2.09 40.545 2.259 ;
      RECT 40.505 2.095 40.52 2.261 ;
      RECT 40.49 2.097 40.505 2.263 ;
      RECT 40.485 2.102 40.49 2.265 ;
      RECT 40.435 2.11 40.485 2.268 ;
      RECT 40.41 2.119 40.435 2.273 ;
      RECT 40.4 2.126 40.41 2.278 ;
      RECT 40.395 2.129 40.4 2.282 ;
      RECT 40.375 2.132 40.395 2.291 ;
      RECT 40.345 2.14 40.375 2.311 ;
      RECT 40.316 2.153 40.345 2.333 ;
      RECT 40.23 2.187 40.316 2.377 ;
      RECT 40.225 2.213 40.23 2.415 ;
      RECT 40.22 2.217 40.225 2.424 ;
      RECT 40.185 2.23 40.22 2.457 ;
      RECT 40.175 2.244 40.185 2.495 ;
      RECT 40.17 2.248 40.175 2.508 ;
      RECT 40.165 2.252 40.17 2.513 ;
      RECT 40.155 2.26 40.165 2.525 ;
      RECT 40.15 2.267 40.155 2.54 ;
      RECT 40.125 2.28 40.15 2.565 ;
      RECT 40.085 2.309 40.125 2.62 ;
      RECT 40.07 2.334 40.085 2.675 ;
      RECT 40.06 2.345 40.07 2.698 ;
      RECT 40.055 2.352 40.06 2.71 ;
      RECT 40.05 2.356 40.055 2.718 ;
      RECT 39.995 2.384 40.05 2.76 ;
      RECT 39.975 2.42 39.995 2.76 ;
      RECT 39.96 2.435 39.975 2.76 ;
      RECT 39.905 2.467 39.96 2.76 ;
      RECT 39.895 2.497 39.905 2.76 ;
      RECT 39.505 2.112 39.69 2.35 ;
      RECT 39.49 2.114 39.7 2.345 ;
      RECT 39.375 2.06 39.635 2.32 ;
      RECT 39.37 2.097 39.635 2.274 ;
      RECT 39.365 2.107 39.635 2.271 ;
      RECT 39.36 2.147 39.7 2.265 ;
      RECT 39.355 2.18 39.7 2.255 ;
      RECT 39.365 2.122 39.715 2.193 ;
      RECT 39.662 3.22 39.675 3.75 ;
      RECT 39.576 3.22 39.675 3.749 ;
      RECT 39.576 3.22 39.68 3.748 ;
      RECT 39.49 3.22 39.68 3.746 ;
      RECT 39.485 3.22 39.68 3.743 ;
      RECT 39.485 3.22 39.69 3.741 ;
      RECT 39.48 3.512 39.69 3.738 ;
      RECT 39.48 3.522 39.695 3.735 ;
      RECT 39.48 3.59 39.7 3.731 ;
      RECT 39.47 3.595 39.7 3.73 ;
      RECT 39.47 3.687 39.705 3.727 ;
      RECT 39.455 3.22 39.715 3.48 ;
      RECT 38.685 2.21 38.73 3.745 ;
      RECT 38.885 2.21 38.915 2.425 ;
      RECT 37.26 1.95 37.38 2.16 ;
      RECT 36.92 1.9 37.18 2.16 ;
      RECT 36.92 1.945 37.215 2.15 ;
      RECT 38.925 2.226 38.93 2.28 ;
      RECT 38.92 2.219 38.925 2.413 ;
      RECT 38.915 2.213 38.92 2.42 ;
      RECT 38.87 2.21 38.885 2.433 ;
      RECT 38.865 2.21 38.87 2.455 ;
      RECT 38.86 2.21 38.865 2.503 ;
      RECT 38.855 2.21 38.86 2.523 ;
      RECT 38.845 2.21 38.855 2.63 ;
      RECT 38.84 2.21 38.845 2.693 ;
      RECT 38.835 2.21 38.84 2.75 ;
      RECT 38.83 2.21 38.835 2.758 ;
      RECT 38.815 2.21 38.83 2.865 ;
      RECT 38.805 2.21 38.815 3 ;
      RECT 38.795 2.21 38.805 3.11 ;
      RECT 38.785 2.21 38.795 3.167 ;
      RECT 38.78 2.21 38.785 3.207 ;
      RECT 38.775 2.21 38.78 3.243 ;
      RECT 38.765 2.21 38.775 3.283 ;
      RECT 38.76 2.21 38.765 3.325 ;
      RECT 38.74 2.21 38.76 3.39 ;
      RECT 38.745 3.535 38.75 3.715 ;
      RECT 38.74 3.517 38.745 3.723 ;
      RECT 38.735 2.21 38.74 3.453 ;
      RECT 38.735 3.497 38.74 3.73 ;
      RECT 38.73 2.21 38.735 3.74 ;
      RECT 38.675 2.21 38.685 2.51 ;
      RECT 38.68 2.757 38.685 3.745 ;
      RECT 38.675 2.822 38.68 3.745 ;
      RECT 38.67 2.211 38.675 2.5 ;
      RECT 38.665 2.887 38.675 3.745 ;
      RECT 38.66 2.212 38.67 2.49 ;
      RECT 38.65 3 38.665 3.745 ;
      RECT 38.655 2.213 38.66 2.48 ;
      RECT 38.635 2.214 38.655 2.458 ;
      RECT 38.64 3.097 38.65 3.745 ;
      RECT 38.635 3.172 38.64 3.745 ;
      RECT 38.625 2.213 38.635 2.435 ;
      RECT 38.63 3.215 38.635 3.745 ;
      RECT 38.625 3.242 38.63 3.745 ;
      RECT 38.615 2.211 38.625 2.423 ;
      RECT 38.62 3.285 38.625 3.745 ;
      RECT 38.615 3.312 38.62 3.745 ;
      RECT 38.605 2.21 38.615 2.41 ;
      RECT 38.61 3.327 38.615 3.745 ;
      RECT 38.57 3.385 38.61 3.745 ;
      RECT 38.6 2.209 38.605 2.395 ;
      RECT 38.595 2.207 38.6 2.388 ;
      RECT 38.585 2.204 38.595 2.378 ;
      RECT 38.58 2.201 38.585 2.363 ;
      RECT 38.565 2.197 38.58 2.356 ;
      RECT 38.56 3.44 38.57 3.745 ;
      RECT 38.56 2.194 38.565 2.351 ;
      RECT 38.545 2.19 38.56 2.345 ;
      RECT 38.555 3.457 38.56 3.745 ;
      RECT 38.545 3.52 38.555 3.745 ;
      RECT 38.465 2.175 38.545 2.325 ;
      RECT 38.54 3.527 38.545 3.74 ;
      RECT 38.535 3.535 38.54 3.73 ;
      RECT 38.455 2.161 38.465 2.309 ;
      RECT 38.44 2.157 38.455 2.307 ;
      RECT 38.43 2.152 38.44 2.303 ;
      RECT 38.405 2.145 38.43 2.295 ;
      RECT 38.4 2.14 38.405 2.29 ;
      RECT 38.39 2.14 38.4 2.288 ;
      RECT 38.38 2.138 38.39 2.286 ;
      RECT 38.35 2.13 38.38 2.28 ;
      RECT 38.335 2.122 38.35 2.273 ;
      RECT 38.315 2.117 38.335 2.266 ;
      RECT 38.31 2.113 38.315 2.261 ;
      RECT 38.28 2.106 38.31 2.255 ;
      RECT 38.255 2.097 38.28 2.245 ;
      RECT 38.225 2.09 38.255 2.237 ;
      RECT 38.2 2.08 38.225 2.228 ;
      RECT 38.185 2.072 38.2 2.222 ;
      RECT 38.16 2.067 38.185 2.217 ;
      RECT 38.15 2.063 38.16 2.212 ;
      RECT 38.13 2.058 38.15 2.207 ;
      RECT 38.095 2.053 38.13 2.2 ;
      RECT 38.035 2.048 38.095 2.193 ;
      RECT 38.022 2.044 38.035 2.191 ;
      RECT 37.936 2.039 38.022 2.188 ;
      RECT 37.85 2.029 37.936 2.184 ;
      RECT 37.809 2.022 37.85 2.181 ;
      RECT 37.723 2.015 37.809 2.178 ;
      RECT 37.637 2.005 37.723 2.174 ;
      RECT 37.551 1.995 37.637 2.169 ;
      RECT 37.465 1.985 37.551 2.165 ;
      RECT 37.455 1.97 37.465 2.163 ;
      RECT 37.445 1.955 37.455 2.163 ;
      RECT 37.38 1.95 37.445 2.162 ;
      RECT 37.215 1.947 37.26 2.155 ;
      RECT 38.46 2.852 38.465 3.043 ;
      RECT 38.455 2.847 38.46 3.05 ;
      RECT 38.441 2.845 38.455 3.056 ;
      RECT 38.355 2.845 38.441 3.058 ;
      RECT 38.351 2.845 38.355 3.061 ;
      RECT 38.265 2.845 38.351 3.079 ;
      RECT 38.255 2.85 38.265 3.098 ;
      RECT 38.245 2.905 38.255 3.102 ;
      RECT 38.22 2.92 38.245 3.109 ;
      RECT 38.18 2.94 38.22 3.122 ;
      RECT 38.175 2.952 38.18 3.132 ;
      RECT 38.16 2.958 38.175 3.137 ;
      RECT 38.155 2.963 38.16 3.141 ;
      RECT 38.135 2.97 38.155 3.146 ;
      RECT 38.065 2.995 38.135 3.163 ;
      RECT 38.025 3.023 38.065 3.183 ;
      RECT 38.02 3.033 38.025 3.191 ;
      RECT 38 3.04 38.02 3.193 ;
      RECT 37.995 3.047 38 3.196 ;
      RECT 37.965 3.055 37.995 3.199 ;
      RECT 37.96 3.06 37.965 3.203 ;
      RECT 37.886 3.064 37.96 3.211 ;
      RECT 37.8 3.073 37.886 3.227 ;
      RECT 37.796 3.078 37.8 3.236 ;
      RECT 37.71 3.083 37.796 3.246 ;
      RECT 37.67 3.091 37.71 3.258 ;
      RECT 37.62 3.097 37.67 3.265 ;
      RECT 37.535 3.106 37.62 3.28 ;
      RECT 37.46 3.117 37.535 3.298 ;
      RECT 37.425 3.124 37.46 3.308 ;
      RECT 37.35 3.132 37.425 3.313 ;
      RECT 37.295 3.141 37.35 3.313 ;
      RECT 37.27 3.146 37.295 3.311 ;
      RECT 37.26 3.149 37.27 3.309 ;
      RECT 37.225 3.151 37.26 3.307 ;
      RECT 37.195 3.153 37.225 3.303 ;
      RECT 37.15 3.152 37.195 3.299 ;
      RECT 37.13 3.147 37.15 3.296 ;
      RECT 37.08 3.132 37.13 3.293 ;
      RECT 37.07 3.117 37.08 3.288 ;
      RECT 37.02 3.102 37.07 3.278 ;
      RECT 36.97 3.077 37.02 3.258 ;
      RECT 36.96 3.062 36.97 3.24 ;
      RECT 36.955 3.06 36.96 3.234 ;
      RECT 36.935 3.055 36.955 3.229 ;
      RECT 36.93 3.047 36.935 3.223 ;
      RECT 36.915 3.041 36.93 3.216 ;
      RECT 36.91 3.036 36.915 3.208 ;
      RECT 36.89 3.031 36.91 3.2 ;
      RECT 36.875 3.024 36.89 3.193 ;
      RECT 36.86 3.018 36.875 3.184 ;
      RECT 36.855 3.012 36.86 3.177 ;
      RECT 36.81 2.987 36.855 3.163 ;
      RECT 36.795 2.957 36.81 3.145 ;
      RECT 36.78 2.94 36.795 3.136 ;
      RECT 36.755 2.92 36.78 3.124 ;
      RECT 36.715 2.89 36.755 3.104 ;
      RECT 36.705 2.86 36.715 3.089 ;
      RECT 36.69 2.85 36.705 3.082 ;
      RECT 36.635 2.815 36.69 3.061 ;
      RECT 36.62 2.778 36.635 3.04 ;
      RECT 36.61 2.765 36.62 3.032 ;
      RECT 36.56 2.735 36.61 3.014 ;
      RECT 36.545 2.665 36.56 2.995 ;
      RECT 36.5 2.665 36.545 2.978 ;
      RECT 36.475 2.665 36.5 2.96 ;
      RECT 36.465 2.665 36.475 2.953 ;
      RECT 36.386 2.665 36.465 2.946 ;
      RECT 36.3 2.665 36.386 2.938 ;
      RECT 36.285 2.697 36.3 2.933 ;
      RECT 36.21 2.707 36.285 2.929 ;
      RECT 36.19 2.717 36.21 2.924 ;
      RECT 36.165 2.717 36.19 2.921 ;
      RECT 36.155 2.707 36.165 2.92 ;
      RECT 36.145 2.68 36.155 2.919 ;
      RECT 36.105 2.675 36.145 2.917 ;
      RECT 36.06 2.675 36.105 2.913 ;
      RECT 36.035 2.675 36.06 2.908 ;
      RECT 35.985 2.675 36.035 2.895 ;
      RECT 35.945 2.68 35.955 2.88 ;
      RECT 35.955 2.675 35.985 2.885 ;
      RECT 37.94 2.455 38.2 2.715 ;
      RECT 37.935 2.477 38.2 2.673 ;
      RECT 37.175 2.305 37.395 2.67 ;
      RECT 37.157 2.392 37.395 2.669 ;
      RECT 37.14 2.397 37.395 2.666 ;
      RECT 37.14 2.397 37.415 2.665 ;
      RECT 37.11 2.407 37.415 2.663 ;
      RECT 37.105 2.422 37.415 2.659 ;
      RECT 37.105 2.422 37.42 2.658 ;
      RECT 37.1 2.48 37.42 2.656 ;
      RECT 37.1 2.48 37.43 2.653 ;
      RECT 37.095 2.545 37.43 2.648 ;
      RECT 37.175 2.305 37.435 2.565 ;
      RECT 35.92 2.135 36.18 2.395 ;
      RECT 35.92 2.178 36.266 2.369 ;
      RECT 35.92 2.178 36.31 2.368 ;
      RECT 35.92 2.178 36.33 2.366 ;
      RECT 35.92 2.178 36.43 2.365 ;
      RECT 35.92 2.178 36.45 2.363 ;
      RECT 35.92 2.178 36.46 2.358 ;
      RECT 36.33 2.145 36.52 2.355 ;
      RECT 36.33 2.147 36.525 2.353 ;
      RECT 36.32 2.152 36.53 2.345 ;
      RECT 36.266 2.176 36.53 2.345 ;
      RECT 36.31 2.17 36.32 2.367 ;
      RECT 36.32 2.15 36.525 2.353 ;
      RECT 35.275 3.21 35.48 3.44 ;
      RECT 35.215 3.16 35.27 3.42 ;
      RECT 35.275 3.16 35.475 3.44 ;
      RECT 36.245 3.475 36.25 3.502 ;
      RECT 36.235 3.385 36.245 3.507 ;
      RECT 36.23 3.307 36.235 3.513 ;
      RECT 36.22 3.297 36.23 3.52 ;
      RECT 36.215 3.287 36.22 3.526 ;
      RECT 36.205 3.282 36.215 3.528 ;
      RECT 36.19 3.274 36.205 3.536 ;
      RECT 36.175 3.265 36.19 3.548 ;
      RECT 36.165 3.257 36.175 3.558 ;
      RECT 36.13 3.175 36.165 3.576 ;
      RECT 36.095 3.175 36.13 3.595 ;
      RECT 36.08 3.175 36.095 3.603 ;
      RECT 36.025 3.175 36.08 3.603 ;
      RECT 35.991 3.175 36.025 3.594 ;
      RECT 35.905 3.175 35.991 3.57 ;
      RECT 35.895 3.235 35.905 3.552 ;
      RECT 35.855 3.237 35.895 3.543 ;
      RECT 35.85 3.239 35.855 3.533 ;
      RECT 35.83 3.241 35.85 3.528 ;
      RECT 35.82 3.244 35.83 3.523 ;
      RECT 35.81 3.245 35.82 3.518 ;
      RECT 35.786 3.246 35.81 3.51 ;
      RECT 35.7 3.251 35.786 3.488 ;
      RECT 35.645 3.25 35.7 3.461 ;
      RECT 35.63 3.243 35.645 3.448 ;
      RECT 35.595 3.238 35.63 3.444 ;
      RECT 35.54 3.23 35.595 3.443 ;
      RECT 35.48 3.217 35.54 3.441 ;
      RECT 35.27 3.16 35.275 3.428 ;
      RECT 35.345 2.53 35.53 2.74 ;
      RECT 35.335 2.535 35.545 2.733 ;
      RECT 35.375 2.44 35.635 2.7 ;
      RECT 35.33 2.597 35.635 2.623 ;
      RECT 34.675 2.39 34.68 3.19 ;
      RECT 34.62 2.44 34.65 3.19 ;
      RECT 34.61 2.44 34.615 2.75 ;
      RECT 34.595 2.44 34.6 2.745 ;
      RECT 34.14 2.485 34.155 2.7 ;
      RECT 34.07 2.485 34.155 2.695 ;
      RECT 35.335 2.065 35.405 2.275 ;
      RECT 35.405 2.072 35.415 2.27 ;
      RECT 35.301 2.065 35.335 2.282 ;
      RECT 35.215 2.065 35.301 2.306 ;
      RECT 35.205 2.07 35.215 2.325 ;
      RECT 35.2 2.082 35.205 2.328 ;
      RECT 35.185 2.097 35.2 2.332 ;
      RECT 35.18 2.115 35.185 2.336 ;
      RECT 35.14 2.125 35.18 2.345 ;
      RECT 35.125 2.132 35.14 2.357 ;
      RECT 35.11 2.137 35.125 2.362 ;
      RECT 35.095 2.14 35.11 2.367 ;
      RECT 35.085 2.142 35.095 2.371 ;
      RECT 35.05 2.149 35.085 2.379 ;
      RECT 35.015 2.157 35.05 2.393 ;
      RECT 35.005 2.163 35.015 2.402 ;
      RECT 35 2.165 35.005 2.404 ;
      RECT 34.98 2.168 35 2.41 ;
      RECT 34.95 2.175 34.98 2.421 ;
      RECT 34.94 2.181 34.95 2.428 ;
      RECT 34.915 2.184 34.94 2.435 ;
      RECT 34.905 2.188 34.915 2.443 ;
      RECT 34.9 2.189 34.905 2.465 ;
      RECT 34.895 2.19 34.9 2.48 ;
      RECT 34.89 2.191 34.895 2.495 ;
      RECT 34.885 2.192 34.89 2.51 ;
      RECT 34.88 2.193 34.885 2.54 ;
      RECT 34.87 2.195 34.88 2.573 ;
      RECT 34.855 2.199 34.87 2.62 ;
      RECT 34.845 2.202 34.855 2.665 ;
      RECT 34.84 2.205 34.845 2.693 ;
      RECT 34.83 2.207 34.84 2.72 ;
      RECT 34.825 2.21 34.83 2.755 ;
      RECT 34.795 2.215 34.825 2.813 ;
      RECT 34.79 2.22 34.795 2.898 ;
      RECT 34.785 2.222 34.79 2.933 ;
      RECT 34.78 2.224 34.785 3.015 ;
      RECT 34.775 2.226 34.78 3.103 ;
      RECT 34.765 2.228 34.775 3.185 ;
      RECT 34.75 2.242 34.765 3.19 ;
      RECT 34.715 2.287 34.75 3.19 ;
      RECT 34.705 2.327 34.715 3.19 ;
      RECT 34.69 2.355 34.705 3.19 ;
      RECT 34.685 2.372 34.69 3.19 ;
      RECT 34.68 2.38 34.685 3.19 ;
      RECT 34.67 2.395 34.675 3.19 ;
      RECT 34.665 2.402 34.67 3.19 ;
      RECT 34.655 2.422 34.665 3.19 ;
      RECT 34.65 2.435 34.655 3.19 ;
      RECT 34.615 2.44 34.62 2.775 ;
      RECT 34.6 2.83 34.62 3.19 ;
      RECT 34.6 2.44 34.61 2.748 ;
      RECT 34.595 2.87 34.6 3.19 ;
      RECT 34.545 2.44 34.595 2.743 ;
      RECT 34.59 2.907 34.595 3.19 ;
      RECT 34.58 2.93 34.59 3.19 ;
      RECT 34.575 2.975 34.58 3.19 ;
      RECT 34.565 2.985 34.575 3.183 ;
      RECT 34.491 2.44 34.545 2.737 ;
      RECT 34.405 2.44 34.491 2.73 ;
      RECT 34.356 2.487 34.405 2.723 ;
      RECT 34.27 2.495 34.356 2.716 ;
      RECT 34.255 2.492 34.27 2.711 ;
      RECT 34.241 2.485 34.255 2.71 ;
      RECT 34.155 2.485 34.241 2.705 ;
      RECT 34.06 2.49 34.07 2.69 ;
      RECT 33.65 1.92 33.665 2.32 ;
      RECT 33.845 1.92 33.85 2.18 ;
      RECT 33.59 1.92 33.635 2.18 ;
      RECT 34.045 3.225 34.05 3.43 ;
      RECT 34.04 3.215 34.045 3.435 ;
      RECT 34.035 3.202 34.04 3.44 ;
      RECT 34.03 3.182 34.035 3.44 ;
      RECT 34.005 3.135 34.03 3.44 ;
      RECT 33.97 3.05 34.005 3.44 ;
      RECT 33.965 2.987 33.97 3.44 ;
      RECT 33.96 2.972 33.965 3.44 ;
      RECT 33.945 2.932 33.96 3.44 ;
      RECT 33.94 2.907 33.945 3.44 ;
      RECT 33.93 2.89 33.94 3.44 ;
      RECT 33.895 2.812 33.93 3.44 ;
      RECT 33.89 2.755 33.895 3.44 ;
      RECT 33.885 2.742 33.89 3.44 ;
      RECT 33.875 2.72 33.885 3.44 ;
      RECT 33.865 2.685 33.875 3.44 ;
      RECT 33.855 2.655 33.865 3.44 ;
      RECT 33.845 2.57 33.855 3.083 ;
      RECT 33.852 3.215 33.855 3.44 ;
      RECT 33.85 3.225 33.852 3.44 ;
      RECT 33.84 3.235 33.85 3.435 ;
      RECT 33.835 1.92 33.845 2.315 ;
      RECT 33.84 2.447 33.845 3.058 ;
      RECT 33.835 2.345 33.84 3.041 ;
      RECT 33.825 1.92 33.835 3.017 ;
      RECT 33.82 1.92 33.825 2.988 ;
      RECT 33.815 1.92 33.82 2.978 ;
      RECT 33.795 1.92 33.815 2.94 ;
      RECT 33.79 1.92 33.795 2.898 ;
      RECT 33.785 1.92 33.79 2.878 ;
      RECT 33.755 1.92 33.785 2.828 ;
      RECT 33.745 1.92 33.755 2.775 ;
      RECT 33.74 1.92 33.745 2.748 ;
      RECT 33.735 1.92 33.74 2.733 ;
      RECT 33.725 1.92 33.735 2.71 ;
      RECT 33.715 1.92 33.725 2.685 ;
      RECT 33.71 1.92 33.715 2.625 ;
      RECT 33.7 1.92 33.71 2.563 ;
      RECT 33.695 1.92 33.7 2.483 ;
      RECT 33.69 1.92 33.695 2.448 ;
      RECT 33.685 1.92 33.69 2.423 ;
      RECT 33.68 1.92 33.685 2.408 ;
      RECT 33.675 1.92 33.68 2.378 ;
      RECT 33.67 1.92 33.675 2.355 ;
      RECT 33.665 1.92 33.67 2.328 ;
      RECT 33.635 1.92 33.65 2.315 ;
      RECT 32.79 3.455 32.975 3.665 ;
      RECT 32.78 3.46 32.99 3.658 ;
      RECT 32.78 3.46 33.01 3.63 ;
      RECT 32.78 3.46 33.025 3.609 ;
      RECT 32.78 3.46 33.04 3.607 ;
      RECT 32.78 3.46 33.05 3.606 ;
      RECT 32.78 3.46 33.08 3.603 ;
      RECT 33.43 3.305 33.69 3.565 ;
      RECT 33.39 3.352 33.69 3.548 ;
      RECT 33.381 3.36 33.39 3.551 ;
      RECT 32.975 3.453 33.69 3.548 ;
      RECT 33.295 3.378 33.381 3.558 ;
      RECT 32.99 3.45 33.69 3.548 ;
      RECT 33.236 3.4 33.295 3.57 ;
      RECT 33.01 3.446 33.69 3.548 ;
      RECT 33.15 3.412 33.236 3.581 ;
      RECT 33.025 3.442 33.69 3.548 ;
      RECT 33.095 3.425 33.15 3.593 ;
      RECT 33.04 3.44 33.69 3.548 ;
      RECT 33.08 3.431 33.095 3.599 ;
      RECT 33.05 3.436 33.69 3.548 ;
      RECT 33.195 2.96 33.455 3.22 ;
      RECT 33.195 2.98 33.565 3.19 ;
      RECT 33.195 2.985 33.575 3.185 ;
      RECT 33.386 2.399 33.465 2.63 ;
      RECT 33.3 2.402 33.515 2.625 ;
      RECT 33.295 2.402 33.515 2.62 ;
      RECT 33.295 2.407 33.525 2.618 ;
      RECT 33.27 2.407 33.525 2.615 ;
      RECT 33.27 2.415 33.535 2.613 ;
      RECT 33.15 2.35 33.41 2.61 ;
      RECT 33.15 2.397 33.46 2.61 ;
      RECT 32.405 2.97 32.41 3.23 ;
      RECT 32.235 2.74 32.24 3.23 ;
      RECT 32.12 2.98 32.125 3.205 ;
      RECT 32.83 2.075 32.835 2.285 ;
      RECT 32.835 2.08 32.85 2.28 ;
      RECT 32.77 2.075 32.83 2.293 ;
      RECT 32.755 2.075 32.77 2.303 ;
      RECT 32.705 2.075 32.755 2.32 ;
      RECT 32.685 2.075 32.705 2.343 ;
      RECT 32.67 2.075 32.685 2.355 ;
      RECT 32.65 2.075 32.67 2.365 ;
      RECT 32.64 2.08 32.65 2.374 ;
      RECT 32.635 2.09 32.64 2.379 ;
      RECT 32.63 2.102 32.635 2.383 ;
      RECT 32.62 2.125 32.63 2.388 ;
      RECT 32.615 2.14 32.62 2.392 ;
      RECT 32.61 2.157 32.615 2.395 ;
      RECT 32.605 2.165 32.61 2.398 ;
      RECT 32.595 2.17 32.605 2.402 ;
      RECT 32.59 2.177 32.595 2.407 ;
      RECT 32.58 2.182 32.59 2.411 ;
      RECT 32.555 2.194 32.58 2.422 ;
      RECT 32.535 2.211 32.555 2.438 ;
      RECT 32.51 2.228 32.535 2.46 ;
      RECT 32.475 2.251 32.51 2.518 ;
      RECT 32.455 2.273 32.475 2.58 ;
      RECT 32.45 2.283 32.455 2.615 ;
      RECT 32.44 2.29 32.45 2.653 ;
      RECT 32.435 2.297 32.44 2.673 ;
      RECT 32.43 2.308 32.435 2.71 ;
      RECT 32.425 2.316 32.43 2.775 ;
      RECT 32.415 2.327 32.425 2.828 ;
      RECT 32.41 2.345 32.415 2.898 ;
      RECT 32.405 2.355 32.41 2.935 ;
      RECT 32.4 2.365 32.405 3.23 ;
      RECT 32.395 2.377 32.4 3.23 ;
      RECT 32.39 2.387 32.395 3.23 ;
      RECT 32.38 2.397 32.39 3.23 ;
      RECT 32.37 2.42 32.38 3.23 ;
      RECT 32.355 2.455 32.37 3.23 ;
      RECT 32.315 2.517 32.355 3.23 ;
      RECT 32.31 2.57 32.315 3.23 ;
      RECT 32.285 2.605 32.31 3.23 ;
      RECT 32.27 2.65 32.285 3.23 ;
      RECT 32.265 2.672 32.27 3.23 ;
      RECT 32.255 2.685 32.265 3.23 ;
      RECT 32.245 2.71 32.255 3.23 ;
      RECT 32.24 2.732 32.245 3.23 ;
      RECT 32.215 2.77 32.235 3.23 ;
      RECT 32.175 2.827 32.215 3.23 ;
      RECT 32.17 2.877 32.175 3.23 ;
      RECT 32.165 2.895 32.17 3.23 ;
      RECT 32.16 2.907 32.165 3.23 ;
      RECT 32.15 2.925 32.16 3.23 ;
      RECT 32.14 2.945 32.15 3.205 ;
      RECT 32.135 2.962 32.14 3.205 ;
      RECT 32.125 2.975 32.135 3.205 ;
      RECT 32.095 2.985 32.12 3.205 ;
      RECT 32.085 2.992 32.095 3.205 ;
      RECT 32.07 3.002 32.085 3.2 ;
      RECT 31.1 2.365 31.39 2.595 ;
      RECT 31.16 0.885 31.33 2.595 ;
      RECT 31.13 0.885 31.48 1.235 ;
      RECT 31.1 0.885 31.48 1.115 ;
      RECT 31.1 7.765 31.39 7.995 ;
      RECT 31.16 6.285 31.33 7.995 ;
      RECT 31.1 6.285 31.39 6.515 ;
      RECT 30.69 2.735 31.02 2.965 ;
      RECT 30.69 2.765 31.19 2.935 ;
      RECT 30.69 2.395 30.88 2.965 ;
      RECT 30.11 2.365 30.4 2.595 ;
      RECT 30.11 2.395 30.88 2.565 ;
      RECT 30.17 0.885 30.34 2.595 ;
      RECT 30.11 0.885 30.4 1.115 ;
      RECT 30.11 7.765 30.4 7.995 ;
      RECT 30.17 6.285 30.34 7.995 ;
      RECT 30.11 6.285 30.4 6.515 ;
      RECT 30.11 6.325 30.96 6.485 ;
      RECT 30.79 5.915 30.96 6.485 ;
      RECT 30.11 6.32 30.5 6.485 ;
      RECT 30.73 5.915 31.02 6.145 ;
      RECT 30.73 5.945 31.19 6.115 ;
      RECT 29.74 2.735 30.03 2.965 ;
      RECT 29.74 2.765 30.2 2.935 ;
      RECT 29.8 1.655 29.965 2.965 ;
      RECT 28.315 1.625 28.605 1.855 ;
      RECT 28.315 1.655 29.965 1.825 ;
      RECT 28.375 0.885 28.545 1.855 ;
      RECT 28.315 0.885 28.605 1.115 ;
      RECT 28.315 7.765 28.605 7.995 ;
      RECT 28.375 7.025 28.545 7.995 ;
      RECT 28.375 7.12 29.965 7.29 ;
      RECT 29.795 5.915 29.965 7.29 ;
      RECT 28.315 7.025 28.605 7.255 ;
      RECT 29.74 5.915 30.03 6.145 ;
      RECT 29.74 5.945 30.2 6.115 ;
      RECT 28.745 1.965 29.095 2.315 ;
      RECT 28.575 2.025 29.095 2.195 ;
      RECT 28.77 6.655 29.095 6.98 ;
      RECT 28.745 6.655 29.095 6.885 ;
      RECT 28.575 6.685 29.095 6.855 ;
      RECT 27.97 2.365 28.29 2.685 ;
      RECT 27.94 2.365 28.29 2.595 ;
      RECT 26.41 2.395 28.29 2.565 ;
      RECT 26.41 1.34 26.58 2.565 ;
      RECT 26.31 1.34 26.66 1.69 ;
      RECT 27.97 6.28 28.29 6.605 ;
      RECT 27.94 6.285 28.29 6.515 ;
      RECT 27.77 6.315 28.29 6.485 ;
      RECT 26.915 2.705 27.265 3.055 ;
      RECT 26.915 2.765 27.405 2.935 ;
      RECT 26.92 5.855 27.27 6.205 ;
      RECT 26.92 5.945 27.405 6.115 ;
      RECT 24.605 2.465 24.79 2.675 ;
      RECT 24.595 2.47 24.805 2.668 ;
      RECT 24.595 2.47 24.891 2.645 ;
      RECT 24.595 2.47 24.95 2.62 ;
      RECT 24.595 2.47 25.005 2.6 ;
      RECT 24.595 2.47 25.015 2.588 ;
      RECT 24.595 2.47 25.21 2.527 ;
      RECT 24.595 2.47 25.24 2.51 ;
      RECT 24.595 2.47 25.26 2.5 ;
      RECT 25.14 2.235 25.4 2.495 ;
      RECT 25.125 2.325 25.14 2.542 ;
      RECT 24.66 2.457 25.4 2.495 ;
      RECT 25.111 2.336 25.125 2.548 ;
      RECT 24.7 2.45 25.4 2.495 ;
      RECT 25.025 2.376 25.111 2.567 ;
      RECT 24.95 2.437 25.4 2.495 ;
      RECT 25.02 2.412 25.025 2.584 ;
      RECT 25.005 2.422 25.4 2.495 ;
      RECT 25.015 2.417 25.02 2.586 ;
      RECT 25.31 2.922 25.315 3.014 ;
      RECT 25.305 2.9 25.31 3.031 ;
      RECT 25.3 2.89 25.305 3.043 ;
      RECT 25.29 2.881 25.3 3.053 ;
      RECT 25.285 2.876 25.29 3.061 ;
      RECT 25.28 2.735 25.285 3.064 ;
      RECT 25.246 2.735 25.28 3.075 ;
      RECT 25.16 2.735 25.246 3.11 ;
      RECT 25.08 2.735 25.16 3.158 ;
      RECT 25.051 2.735 25.08 3.182 ;
      RECT 24.965 2.735 25.051 3.188 ;
      RECT 24.96 2.919 24.965 3.193 ;
      RECT 24.925 2.93 24.96 3.196 ;
      RECT 24.9 2.945 24.925 3.2 ;
      RECT 24.886 2.954 24.9 3.202 ;
      RECT 24.8 2.981 24.886 3.208 ;
      RECT 24.735 3.022 24.8 3.217 ;
      RECT 24.72 3.042 24.735 3.222 ;
      RECT 24.69 3.052 24.72 3.225 ;
      RECT 24.685 3.062 24.69 3.228 ;
      RECT 24.655 3.067 24.685 3.23 ;
      RECT 24.635 3.072 24.655 3.234 ;
      RECT 24.55 3.075 24.635 3.241 ;
      RECT 24.535 3.072 24.55 3.247 ;
      RECT 24.525 3.069 24.535 3.249 ;
      RECT 24.505 3.066 24.525 3.251 ;
      RECT 24.485 3.062 24.505 3.252 ;
      RECT 24.47 3.058 24.485 3.254 ;
      RECT 24.46 3.055 24.47 3.255 ;
      RECT 24.42 3.049 24.46 3.253 ;
      RECT 24.41 3.044 24.42 3.251 ;
      RECT 24.395 3.041 24.41 3.247 ;
      RECT 24.37 3.036 24.395 3.24 ;
      RECT 24.32 3.027 24.37 3.228 ;
      RECT 24.25 3.013 24.32 3.21 ;
      RECT 24.192 2.998 24.25 3.192 ;
      RECT 24.106 2.981 24.192 3.172 ;
      RECT 24.02 2.96 24.106 3.147 ;
      RECT 23.97 2.945 24.02 3.128 ;
      RECT 23.966 2.939 23.97 3.12 ;
      RECT 23.88 2.929 23.966 3.107 ;
      RECT 23.845 2.914 23.88 3.09 ;
      RECT 23.83 2.907 23.845 3.083 ;
      RECT 23.77 2.895 23.83 3.071 ;
      RECT 23.75 2.882 23.77 3.059 ;
      RECT 23.71 2.873 23.75 3.051 ;
      RECT 23.705 2.865 23.71 3.044 ;
      RECT 23.625 2.855 23.705 3.03 ;
      RECT 23.61 2.842 23.625 3.015 ;
      RECT 23.605 2.84 23.61 3.013 ;
      RECT 23.526 2.828 23.605 3 ;
      RECT 23.44 2.803 23.526 2.975 ;
      RECT 23.425 2.772 23.44 2.96 ;
      RECT 23.41 2.747 23.425 2.956 ;
      RECT 23.395 2.74 23.41 2.952 ;
      RECT 23.22 2.745 23.225 2.948 ;
      RECT 23.215 2.75 23.22 2.943 ;
      RECT 23.225 2.74 23.395 2.95 ;
      RECT 23.94 2.5 24.045 2.76 ;
      RECT 24.755 2.025 24.76 2.25 ;
      RECT 24.885 2.025 24.94 2.235 ;
      RECT 24.94 2.03 24.95 2.228 ;
      RECT 24.846 2.025 24.885 2.238 ;
      RECT 24.76 2.025 24.846 2.245 ;
      RECT 24.74 2.03 24.755 2.251 ;
      RECT 24.73 2.07 24.74 2.253 ;
      RECT 24.7 2.08 24.73 2.255 ;
      RECT 24.695 2.085 24.7 2.257 ;
      RECT 24.67 2.09 24.695 2.259 ;
      RECT 24.655 2.095 24.67 2.261 ;
      RECT 24.64 2.097 24.655 2.263 ;
      RECT 24.635 2.102 24.64 2.265 ;
      RECT 24.585 2.11 24.635 2.268 ;
      RECT 24.56 2.119 24.585 2.273 ;
      RECT 24.55 2.126 24.56 2.278 ;
      RECT 24.545 2.129 24.55 2.282 ;
      RECT 24.525 2.132 24.545 2.291 ;
      RECT 24.495 2.14 24.525 2.311 ;
      RECT 24.466 2.153 24.495 2.333 ;
      RECT 24.38 2.187 24.466 2.377 ;
      RECT 24.375 2.213 24.38 2.415 ;
      RECT 24.37 2.217 24.375 2.424 ;
      RECT 24.335 2.23 24.37 2.457 ;
      RECT 24.325 2.244 24.335 2.495 ;
      RECT 24.32 2.248 24.325 2.508 ;
      RECT 24.315 2.252 24.32 2.513 ;
      RECT 24.305 2.26 24.315 2.525 ;
      RECT 24.3 2.267 24.305 2.54 ;
      RECT 24.275 2.28 24.3 2.565 ;
      RECT 24.235 2.309 24.275 2.62 ;
      RECT 24.22 2.334 24.235 2.675 ;
      RECT 24.21 2.345 24.22 2.698 ;
      RECT 24.205 2.352 24.21 2.71 ;
      RECT 24.2 2.356 24.205 2.718 ;
      RECT 24.145 2.384 24.2 2.76 ;
      RECT 24.125 2.42 24.145 2.76 ;
      RECT 24.11 2.435 24.125 2.76 ;
      RECT 24.055 2.467 24.11 2.76 ;
      RECT 24.045 2.497 24.055 2.76 ;
      RECT 23.655 2.112 23.84 2.35 ;
      RECT 23.64 2.114 23.85 2.345 ;
      RECT 23.525 2.06 23.785 2.32 ;
      RECT 23.52 2.097 23.785 2.274 ;
      RECT 23.515 2.107 23.785 2.271 ;
      RECT 23.51 2.147 23.85 2.265 ;
      RECT 23.505 2.18 23.85 2.255 ;
      RECT 23.515 2.122 23.865 2.193 ;
      RECT 23.812 3.22 23.825 3.75 ;
      RECT 23.726 3.22 23.825 3.749 ;
      RECT 23.726 3.22 23.83 3.748 ;
      RECT 23.64 3.22 23.83 3.746 ;
      RECT 23.635 3.22 23.83 3.743 ;
      RECT 23.635 3.22 23.84 3.741 ;
      RECT 23.63 3.512 23.84 3.738 ;
      RECT 23.63 3.522 23.845 3.735 ;
      RECT 23.63 3.59 23.85 3.731 ;
      RECT 23.62 3.595 23.85 3.73 ;
      RECT 23.62 3.687 23.855 3.727 ;
      RECT 23.605 3.22 23.865 3.48 ;
      RECT 22.835 2.21 22.88 3.745 ;
      RECT 23.035 2.21 23.065 2.425 ;
      RECT 21.41 1.95 21.53 2.16 ;
      RECT 21.07 1.9 21.33 2.16 ;
      RECT 21.07 1.945 21.365 2.15 ;
      RECT 23.075 2.226 23.08 2.28 ;
      RECT 23.07 2.219 23.075 2.413 ;
      RECT 23.065 2.213 23.07 2.42 ;
      RECT 23.02 2.21 23.035 2.433 ;
      RECT 23.015 2.21 23.02 2.455 ;
      RECT 23.01 2.21 23.015 2.503 ;
      RECT 23.005 2.21 23.01 2.523 ;
      RECT 22.995 2.21 23.005 2.63 ;
      RECT 22.99 2.21 22.995 2.693 ;
      RECT 22.985 2.21 22.99 2.75 ;
      RECT 22.98 2.21 22.985 2.758 ;
      RECT 22.965 2.21 22.98 2.865 ;
      RECT 22.955 2.21 22.965 3 ;
      RECT 22.945 2.21 22.955 3.11 ;
      RECT 22.935 2.21 22.945 3.167 ;
      RECT 22.93 2.21 22.935 3.207 ;
      RECT 22.925 2.21 22.93 3.243 ;
      RECT 22.915 2.21 22.925 3.283 ;
      RECT 22.91 2.21 22.915 3.325 ;
      RECT 22.89 2.21 22.91 3.39 ;
      RECT 22.895 3.535 22.9 3.715 ;
      RECT 22.89 3.517 22.895 3.723 ;
      RECT 22.885 2.21 22.89 3.453 ;
      RECT 22.885 3.497 22.89 3.73 ;
      RECT 22.88 2.21 22.885 3.74 ;
      RECT 22.825 2.21 22.835 2.51 ;
      RECT 22.83 2.757 22.835 3.745 ;
      RECT 22.825 2.822 22.83 3.745 ;
      RECT 22.82 2.211 22.825 2.5 ;
      RECT 22.815 2.887 22.825 3.745 ;
      RECT 22.81 2.212 22.82 2.49 ;
      RECT 22.8 3 22.815 3.745 ;
      RECT 22.805 2.213 22.81 2.48 ;
      RECT 22.785 2.214 22.805 2.458 ;
      RECT 22.79 3.097 22.8 3.745 ;
      RECT 22.785 3.172 22.79 3.745 ;
      RECT 22.775 2.213 22.785 2.435 ;
      RECT 22.78 3.215 22.785 3.745 ;
      RECT 22.775 3.242 22.78 3.745 ;
      RECT 22.765 2.211 22.775 2.423 ;
      RECT 22.77 3.285 22.775 3.745 ;
      RECT 22.765 3.312 22.77 3.745 ;
      RECT 22.755 2.21 22.765 2.41 ;
      RECT 22.76 3.327 22.765 3.745 ;
      RECT 22.72 3.385 22.76 3.745 ;
      RECT 22.75 2.209 22.755 2.395 ;
      RECT 22.745 2.207 22.75 2.388 ;
      RECT 22.735 2.204 22.745 2.378 ;
      RECT 22.73 2.201 22.735 2.363 ;
      RECT 22.715 2.197 22.73 2.356 ;
      RECT 22.71 3.44 22.72 3.745 ;
      RECT 22.71 2.194 22.715 2.351 ;
      RECT 22.695 2.19 22.71 2.345 ;
      RECT 22.705 3.457 22.71 3.745 ;
      RECT 22.695 3.52 22.705 3.745 ;
      RECT 22.615 2.175 22.695 2.325 ;
      RECT 22.69 3.527 22.695 3.74 ;
      RECT 22.685 3.535 22.69 3.73 ;
      RECT 22.605 2.161 22.615 2.309 ;
      RECT 22.59 2.157 22.605 2.307 ;
      RECT 22.58 2.152 22.59 2.303 ;
      RECT 22.555 2.145 22.58 2.295 ;
      RECT 22.55 2.14 22.555 2.29 ;
      RECT 22.54 2.14 22.55 2.288 ;
      RECT 22.53 2.138 22.54 2.286 ;
      RECT 22.5 2.13 22.53 2.28 ;
      RECT 22.485 2.122 22.5 2.273 ;
      RECT 22.465 2.117 22.485 2.266 ;
      RECT 22.46 2.113 22.465 2.261 ;
      RECT 22.43 2.106 22.46 2.255 ;
      RECT 22.405 2.097 22.43 2.245 ;
      RECT 22.375 2.09 22.405 2.237 ;
      RECT 22.35 2.08 22.375 2.228 ;
      RECT 22.335 2.072 22.35 2.222 ;
      RECT 22.31 2.067 22.335 2.217 ;
      RECT 22.3 2.063 22.31 2.212 ;
      RECT 22.28 2.058 22.3 2.207 ;
      RECT 22.245 2.053 22.28 2.2 ;
      RECT 22.185 2.048 22.245 2.193 ;
      RECT 22.172 2.044 22.185 2.191 ;
      RECT 22.086 2.039 22.172 2.188 ;
      RECT 22 2.029 22.086 2.184 ;
      RECT 21.959 2.022 22 2.181 ;
      RECT 21.873 2.015 21.959 2.178 ;
      RECT 21.787 2.005 21.873 2.174 ;
      RECT 21.701 1.995 21.787 2.169 ;
      RECT 21.615 1.985 21.701 2.165 ;
      RECT 21.605 1.97 21.615 2.163 ;
      RECT 21.595 1.955 21.605 2.163 ;
      RECT 21.53 1.95 21.595 2.162 ;
      RECT 21.365 1.947 21.41 2.155 ;
      RECT 22.61 2.852 22.615 3.043 ;
      RECT 22.605 2.847 22.61 3.05 ;
      RECT 22.591 2.845 22.605 3.056 ;
      RECT 22.505 2.845 22.591 3.058 ;
      RECT 22.501 2.845 22.505 3.061 ;
      RECT 22.415 2.845 22.501 3.079 ;
      RECT 22.405 2.85 22.415 3.098 ;
      RECT 22.395 2.905 22.405 3.102 ;
      RECT 22.37 2.92 22.395 3.109 ;
      RECT 22.33 2.94 22.37 3.122 ;
      RECT 22.325 2.952 22.33 3.132 ;
      RECT 22.31 2.958 22.325 3.137 ;
      RECT 22.305 2.963 22.31 3.141 ;
      RECT 22.285 2.97 22.305 3.146 ;
      RECT 22.215 2.995 22.285 3.163 ;
      RECT 22.175 3.023 22.215 3.183 ;
      RECT 22.17 3.033 22.175 3.191 ;
      RECT 22.15 3.04 22.17 3.193 ;
      RECT 22.145 3.047 22.15 3.196 ;
      RECT 22.115 3.055 22.145 3.199 ;
      RECT 22.11 3.06 22.115 3.203 ;
      RECT 22.036 3.064 22.11 3.211 ;
      RECT 21.95 3.073 22.036 3.227 ;
      RECT 21.946 3.078 21.95 3.236 ;
      RECT 21.86 3.083 21.946 3.246 ;
      RECT 21.82 3.091 21.86 3.258 ;
      RECT 21.77 3.097 21.82 3.265 ;
      RECT 21.685 3.106 21.77 3.28 ;
      RECT 21.61 3.117 21.685 3.298 ;
      RECT 21.575 3.124 21.61 3.308 ;
      RECT 21.5 3.132 21.575 3.313 ;
      RECT 21.445 3.141 21.5 3.313 ;
      RECT 21.42 3.146 21.445 3.311 ;
      RECT 21.41 3.149 21.42 3.309 ;
      RECT 21.375 3.151 21.41 3.307 ;
      RECT 21.345 3.153 21.375 3.303 ;
      RECT 21.3 3.152 21.345 3.299 ;
      RECT 21.28 3.147 21.3 3.296 ;
      RECT 21.23 3.132 21.28 3.293 ;
      RECT 21.22 3.117 21.23 3.288 ;
      RECT 21.17 3.102 21.22 3.278 ;
      RECT 21.12 3.077 21.17 3.258 ;
      RECT 21.11 3.062 21.12 3.24 ;
      RECT 21.105 3.06 21.11 3.234 ;
      RECT 21.085 3.055 21.105 3.229 ;
      RECT 21.08 3.047 21.085 3.223 ;
      RECT 21.065 3.041 21.08 3.216 ;
      RECT 21.06 3.036 21.065 3.208 ;
      RECT 21.04 3.031 21.06 3.2 ;
      RECT 21.025 3.024 21.04 3.193 ;
      RECT 21.01 3.018 21.025 3.184 ;
      RECT 21.005 3.012 21.01 3.177 ;
      RECT 20.96 2.987 21.005 3.163 ;
      RECT 20.945 2.957 20.96 3.145 ;
      RECT 20.93 2.94 20.945 3.136 ;
      RECT 20.905 2.92 20.93 3.124 ;
      RECT 20.865 2.89 20.905 3.104 ;
      RECT 20.855 2.86 20.865 3.089 ;
      RECT 20.84 2.85 20.855 3.082 ;
      RECT 20.785 2.815 20.84 3.061 ;
      RECT 20.77 2.778 20.785 3.04 ;
      RECT 20.76 2.765 20.77 3.032 ;
      RECT 20.71 2.735 20.76 3.014 ;
      RECT 20.695 2.665 20.71 2.995 ;
      RECT 20.65 2.665 20.695 2.978 ;
      RECT 20.625 2.665 20.65 2.96 ;
      RECT 20.615 2.665 20.625 2.953 ;
      RECT 20.536 2.665 20.615 2.946 ;
      RECT 20.45 2.665 20.536 2.938 ;
      RECT 20.435 2.697 20.45 2.933 ;
      RECT 20.36 2.707 20.435 2.929 ;
      RECT 20.34 2.717 20.36 2.924 ;
      RECT 20.315 2.717 20.34 2.921 ;
      RECT 20.305 2.707 20.315 2.92 ;
      RECT 20.295 2.68 20.305 2.919 ;
      RECT 20.255 2.675 20.295 2.917 ;
      RECT 20.21 2.675 20.255 2.913 ;
      RECT 20.185 2.675 20.21 2.908 ;
      RECT 20.135 2.675 20.185 2.895 ;
      RECT 20.095 2.68 20.105 2.88 ;
      RECT 20.105 2.675 20.135 2.885 ;
      RECT 22.09 2.455 22.35 2.715 ;
      RECT 22.085 2.477 22.35 2.673 ;
      RECT 21.325 2.305 21.545 2.67 ;
      RECT 21.307 2.392 21.545 2.669 ;
      RECT 21.29 2.397 21.545 2.666 ;
      RECT 21.29 2.397 21.565 2.665 ;
      RECT 21.26 2.407 21.565 2.663 ;
      RECT 21.255 2.422 21.565 2.659 ;
      RECT 21.255 2.422 21.57 2.658 ;
      RECT 21.25 2.48 21.57 2.656 ;
      RECT 21.25 2.48 21.58 2.653 ;
      RECT 21.245 2.545 21.58 2.648 ;
      RECT 21.325 2.305 21.585 2.565 ;
      RECT 20.07 2.135 20.33 2.395 ;
      RECT 20.07 2.178 20.416 2.369 ;
      RECT 20.07 2.178 20.46 2.368 ;
      RECT 20.07 2.178 20.48 2.366 ;
      RECT 20.07 2.178 20.58 2.365 ;
      RECT 20.07 2.178 20.6 2.363 ;
      RECT 20.07 2.178 20.61 2.358 ;
      RECT 20.48 2.145 20.67 2.355 ;
      RECT 20.48 2.147 20.675 2.353 ;
      RECT 20.47 2.152 20.68 2.345 ;
      RECT 20.416 2.176 20.68 2.345 ;
      RECT 20.46 2.17 20.47 2.367 ;
      RECT 20.47 2.15 20.675 2.353 ;
      RECT 19.425 3.21 19.63 3.44 ;
      RECT 19.365 3.16 19.42 3.42 ;
      RECT 19.425 3.16 19.625 3.44 ;
      RECT 20.395 3.475 20.4 3.502 ;
      RECT 20.385 3.385 20.395 3.507 ;
      RECT 20.38 3.307 20.385 3.513 ;
      RECT 20.37 3.297 20.38 3.52 ;
      RECT 20.365 3.287 20.37 3.526 ;
      RECT 20.355 3.282 20.365 3.528 ;
      RECT 20.34 3.274 20.355 3.536 ;
      RECT 20.325 3.265 20.34 3.548 ;
      RECT 20.315 3.257 20.325 3.558 ;
      RECT 20.28 3.175 20.315 3.576 ;
      RECT 20.245 3.175 20.28 3.595 ;
      RECT 20.23 3.175 20.245 3.603 ;
      RECT 20.175 3.175 20.23 3.603 ;
      RECT 20.141 3.175 20.175 3.594 ;
      RECT 20.055 3.175 20.141 3.57 ;
      RECT 20.045 3.235 20.055 3.552 ;
      RECT 20.005 3.237 20.045 3.543 ;
      RECT 20 3.239 20.005 3.533 ;
      RECT 19.98 3.241 20 3.528 ;
      RECT 19.97 3.244 19.98 3.523 ;
      RECT 19.96 3.245 19.97 3.518 ;
      RECT 19.936 3.246 19.96 3.51 ;
      RECT 19.85 3.251 19.936 3.488 ;
      RECT 19.795 3.25 19.85 3.461 ;
      RECT 19.78 3.243 19.795 3.448 ;
      RECT 19.745 3.238 19.78 3.444 ;
      RECT 19.69 3.23 19.745 3.443 ;
      RECT 19.63 3.217 19.69 3.441 ;
      RECT 19.42 3.16 19.425 3.428 ;
      RECT 19.495 2.53 19.68 2.74 ;
      RECT 19.485 2.535 19.695 2.733 ;
      RECT 19.525 2.44 19.785 2.7 ;
      RECT 19.48 2.597 19.785 2.623 ;
      RECT 18.825 2.39 18.83 3.19 ;
      RECT 18.77 2.44 18.8 3.19 ;
      RECT 18.76 2.44 18.765 2.75 ;
      RECT 18.745 2.44 18.75 2.745 ;
      RECT 18.29 2.485 18.305 2.7 ;
      RECT 18.22 2.485 18.305 2.695 ;
      RECT 19.485 2.065 19.555 2.275 ;
      RECT 19.555 2.072 19.565 2.27 ;
      RECT 19.451 2.065 19.485 2.282 ;
      RECT 19.365 2.065 19.451 2.306 ;
      RECT 19.355 2.07 19.365 2.325 ;
      RECT 19.35 2.082 19.355 2.328 ;
      RECT 19.335 2.097 19.35 2.332 ;
      RECT 19.33 2.115 19.335 2.336 ;
      RECT 19.29 2.125 19.33 2.345 ;
      RECT 19.275 2.132 19.29 2.357 ;
      RECT 19.26 2.137 19.275 2.362 ;
      RECT 19.245 2.14 19.26 2.367 ;
      RECT 19.235 2.142 19.245 2.371 ;
      RECT 19.2 2.149 19.235 2.379 ;
      RECT 19.165 2.157 19.2 2.393 ;
      RECT 19.155 2.163 19.165 2.402 ;
      RECT 19.15 2.165 19.155 2.404 ;
      RECT 19.13 2.168 19.15 2.41 ;
      RECT 19.1 2.175 19.13 2.421 ;
      RECT 19.09 2.181 19.1 2.428 ;
      RECT 19.065 2.184 19.09 2.435 ;
      RECT 19.055 2.188 19.065 2.443 ;
      RECT 19.05 2.189 19.055 2.465 ;
      RECT 19.045 2.19 19.05 2.48 ;
      RECT 19.04 2.191 19.045 2.495 ;
      RECT 19.035 2.192 19.04 2.51 ;
      RECT 19.03 2.193 19.035 2.54 ;
      RECT 19.02 2.195 19.03 2.573 ;
      RECT 19.005 2.199 19.02 2.62 ;
      RECT 18.995 2.202 19.005 2.665 ;
      RECT 18.99 2.205 18.995 2.693 ;
      RECT 18.98 2.207 18.99 2.72 ;
      RECT 18.975 2.21 18.98 2.755 ;
      RECT 18.945 2.215 18.975 2.813 ;
      RECT 18.94 2.22 18.945 2.898 ;
      RECT 18.935 2.222 18.94 2.933 ;
      RECT 18.93 2.224 18.935 3.015 ;
      RECT 18.925 2.226 18.93 3.103 ;
      RECT 18.915 2.228 18.925 3.185 ;
      RECT 18.9 2.242 18.915 3.19 ;
      RECT 18.865 2.287 18.9 3.19 ;
      RECT 18.855 2.327 18.865 3.19 ;
      RECT 18.84 2.355 18.855 3.19 ;
      RECT 18.835 2.372 18.84 3.19 ;
      RECT 18.83 2.38 18.835 3.19 ;
      RECT 18.82 2.395 18.825 3.19 ;
      RECT 18.815 2.402 18.82 3.19 ;
      RECT 18.805 2.422 18.815 3.19 ;
      RECT 18.8 2.435 18.805 3.19 ;
      RECT 18.765 2.44 18.77 2.775 ;
      RECT 18.75 2.83 18.77 3.19 ;
      RECT 18.75 2.44 18.76 2.748 ;
      RECT 18.745 2.87 18.75 3.19 ;
      RECT 18.695 2.44 18.745 2.743 ;
      RECT 18.74 2.907 18.745 3.19 ;
      RECT 18.73 2.93 18.74 3.19 ;
      RECT 18.725 2.975 18.73 3.19 ;
      RECT 18.715 2.985 18.725 3.183 ;
      RECT 18.641 2.44 18.695 2.737 ;
      RECT 18.555 2.44 18.641 2.73 ;
      RECT 18.506 2.487 18.555 2.723 ;
      RECT 18.42 2.495 18.506 2.716 ;
      RECT 18.405 2.492 18.42 2.711 ;
      RECT 18.391 2.485 18.405 2.71 ;
      RECT 18.305 2.485 18.391 2.705 ;
      RECT 18.21 2.49 18.22 2.69 ;
      RECT 17.8 1.92 17.815 2.32 ;
      RECT 17.995 1.92 18 2.18 ;
      RECT 17.74 1.92 17.785 2.18 ;
      RECT 18.195 3.225 18.2 3.43 ;
      RECT 18.19 3.215 18.195 3.435 ;
      RECT 18.185 3.202 18.19 3.44 ;
      RECT 18.18 3.182 18.185 3.44 ;
      RECT 18.155 3.135 18.18 3.44 ;
      RECT 18.12 3.05 18.155 3.44 ;
      RECT 18.115 2.987 18.12 3.44 ;
      RECT 18.11 2.972 18.115 3.44 ;
      RECT 18.095 2.932 18.11 3.44 ;
      RECT 18.09 2.907 18.095 3.44 ;
      RECT 18.08 2.89 18.09 3.44 ;
      RECT 18.045 2.812 18.08 3.44 ;
      RECT 18.04 2.755 18.045 3.44 ;
      RECT 18.035 2.742 18.04 3.44 ;
      RECT 18.025 2.72 18.035 3.44 ;
      RECT 18.015 2.685 18.025 3.44 ;
      RECT 18.005 2.655 18.015 3.44 ;
      RECT 17.995 2.57 18.005 3.083 ;
      RECT 18.002 3.215 18.005 3.44 ;
      RECT 18 3.225 18.002 3.44 ;
      RECT 17.99 3.235 18 3.435 ;
      RECT 17.985 1.92 17.995 2.315 ;
      RECT 17.99 2.447 17.995 3.058 ;
      RECT 17.985 2.345 17.99 3.041 ;
      RECT 17.975 1.92 17.985 3.017 ;
      RECT 17.97 1.92 17.975 2.988 ;
      RECT 17.965 1.92 17.97 2.978 ;
      RECT 17.945 1.92 17.965 2.94 ;
      RECT 17.94 1.92 17.945 2.898 ;
      RECT 17.935 1.92 17.94 2.878 ;
      RECT 17.905 1.92 17.935 2.828 ;
      RECT 17.895 1.92 17.905 2.775 ;
      RECT 17.89 1.92 17.895 2.748 ;
      RECT 17.885 1.92 17.89 2.733 ;
      RECT 17.875 1.92 17.885 2.71 ;
      RECT 17.865 1.92 17.875 2.685 ;
      RECT 17.86 1.92 17.865 2.625 ;
      RECT 17.85 1.92 17.86 2.563 ;
      RECT 17.845 1.92 17.85 2.483 ;
      RECT 17.84 1.92 17.845 2.448 ;
      RECT 17.835 1.92 17.84 2.423 ;
      RECT 17.83 1.92 17.835 2.408 ;
      RECT 17.825 1.92 17.83 2.378 ;
      RECT 17.82 1.92 17.825 2.355 ;
      RECT 17.815 1.92 17.82 2.328 ;
      RECT 17.785 1.92 17.8 2.315 ;
      RECT 16.94 3.455 17.125 3.665 ;
      RECT 16.93 3.46 17.14 3.658 ;
      RECT 16.93 3.46 17.16 3.63 ;
      RECT 16.93 3.46 17.175 3.609 ;
      RECT 16.93 3.46 17.19 3.607 ;
      RECT 16.93 3.46 17.2 3.606 ;
      RECT 16.93 3.46 17.23 3.603 ;
      RECT 17.58 3.305 17.84 3.565 ;
      RECT 17.54 3.352 17.84 3.548 ;
      RECT 17.531 3.36 17.54 3.551 ;
      RECT 17.125 3.453 17.84 3.548 ;
      RECT 17.445 3.378 17.531 3.558 ;
      RECT 17.14 3.45 17.84 3.548 ;
      RECT 17.386 3.4 17.445 3.57 ;
      RECT 17.16 3.446 17.84 3.548 ;
      RECT 17.3 3.412 17.386 3.581 ;
      RECT 17.175 3.442 17.84 3.548 ;
      RECT 17.245 3.425 17.3 3.593 ;
      RECT 17.19 3.44 17.84 3.548 ;
      RECT 17.23 3.431 17.245 3.599 ;
      RECT 17.2 3.436 17.84 3.548 ;
      RECT 17.345 2.96 17.605 3.22 ;
      RECT 17.345 2.98 17.715 3.19 ;
      RECT 17.345 2.985 17.725 3.185 ;
      RECT 17.536 2.399 17.615 2.63 ;
      RECT 17.45 2.402 17.665 2.625 ;
      RECT 17.445 2.402 17.665 2.62 ;
      RECT 17.445 2.407 17.675 2.618 ;
      RECT 17.42 2.407 17.675 2.615 ;
      RECT 17.42 2.415 17.685 2.613 ;
      RECT 17.3 2.35 17.56 2.61 ;
      RECT 17.3 2.397 17.61 2.61 ;
      RECT 16.555 2.97 16.56 3.23 ;
      RECT 16.385 2.74 16.39 3.23 ;
      RECT 16.27 2.98 16.275 3.205 ;
      RECT 16.98 2.075 16.985 2.285 ;
      RECT 16.985 2.08 17 2.28 ;
      RECT 16.92 2.075 16.98 2.293 ;
      RECT 16.905 2.075 16.92 2.303 ;
      RECT 16.855 2.075 16.905 2.32 ;
      RECT 16.835 2.075 16.855 2.343 ;
      RECT 16.82 2.075 16.835 2.355 ;
      RECT 16.8 2.075 16.82 2.365 ;
      RECT 16.79 2.08 16.8 2.374 ;
      RECT 16.785 2.09 16.79 2.379 ;
      RECT 16.78 2.102 16.785 2.383 ;
      RECT 16.77 2.125 16.78 2.388 ;
      RECT 16.765 2.14 16.77 2.392 ;
      RECT 16.76 2.157 16.765 2.395 ;
      RECT 16.755 2.165 16.76 2.398 ;
      RECT 16.745 2.17 16.755 2.402 ;
      RECT 16.74 2.177 16.745 2.407 ;
      RECT 16.73 2.182 16.74 2.411 ;
      RECT 16.705 2.194 16.73 2.422 ;
      RECT 16.685 2.211 16.705 2.438 ;
      RECT 16.66 2.228 16.685 2.46 ;
      RECT 16.625 2.251 16.66 2.518 ;
      RECT 16.605 2.273 16.625 2.58 ;
      RECT 16.6 2.283 16.605 2.615 ;
      RECT 16.59 2.29 16.6 2.653 ;
      RECT 16.585 2.297 16.59 2.673 ;
      RECT 16.58 2.308 16.585 2.71 ;
      RECT 16.575 2.316 16.58 2.775 ;
      RECT 16.565 2.327 16.575 2.828 ;
      RECT 16.56 2.345 16.565 2.898 ;
      RECT 16.555 2.355 16.56 2.935 ;
      RECT 16.55 2.365 16.555 3.23 ;
      RECT 16.545 2.377 16.55 3.23 ;
      RECT 16.54 2.387 16.545 3.23 ;
      RECT 16.53 2.397 16.54 3.23 ;
      RECT 16.52 2.42 16.53 3.23 ;
      RECT 16.505 2.455 16.52 3.23 ;
      RECT 16.465 2.517 16.505 3.23 ;
      RECT 16.46 2.57 16.465 3.23 ;
      RECT 16.435 2.605 16.46 3.23 ;
      RECT 16.42 2.65 16.435 3.23 ;
      RECT 16.415 2.672 16.42 3.23 ;
      RECT 16.405 2.685 16.415 3.23 ;
      RECT 16.395 2.71 16.405 3.23 ;
      RECT 16.39 2.732 16.395 3.23 ;
      RECT 16.365 2.77 16.385 3.23 ;
      RECT 16.325 2.827 16.365 3.23 ;
      RECT 16.32 2.877 16.325 3.23 ;
      RECT 16.315 2.895 16.32 3.23 ;
      RECT 16.31 2.907 16.315 3.23 ;
      RECT 16.3 2.925 16.31 3.23 ;
      RECT 16.29 2.945 16.3 3.205 ;
      RECT 16.285 2.962 16.29 3.205 ;
      RECT 16.275 2.975 16.285 3.205 ;
      RECT 16.245 2.985 16.27 3.205 ;
      RECT 16.235 2.992 16.245 3.205 ;
      RECT 16.22 3.002 16.235 3.2 ;
      RECT 15.25 2.365 15.54 2.595 ;
      RECT 15.31 0.885 15.48 2.595 ;
      RECT 15.28 0.885 15.63 1.235 ;
      RECT 15.25 0.885 15.63 1.115 ;
      RECT 15.25 7.765 15.54 7.995 ;
      RECT 15.31 6.285 15.48 7.995 ;
      RECT 15.25 6.285 15.54 6.515 ;
      RECT 14.84 2.735 15.17 2.965 ;
      RECT 14.84 2.765 15.34 2.935 ;
      RECT 14.84 2.395 15.03 2.965 ;
      RECT 14.26 2.365 14.55 2.595 ;
      RECT 14.26 2.395 15.03 2.565 ;
      RECT 14.32 0.885 14.49 2.595 ;
      RECT 14.26 0.885 14.55 1.115 ;
      RECT 14.26 7.765 14.55 7.995 ;
      RECT 14.32 6.285 14.49 7.995 ;
      RECT 14.26 6.285 14.55 6.515 ;
      RECT 14.26 6.325 15.11 6.485 ;
      RECT 14.94 5.915 15.11 6.485 ;
      RECT 14.26 6.32 14.65 6.485 ;
      RECT 14.88 5.915 15.17 6.145 ;
      RECT 14.88 5.945 15.34 6.115 ;
      RECT 13.89 2.735 14.18 2.965 ;
      RECT 13.89 2.765 14.35 2.935 ;
      RECT 13.95 1.655 14.115 2.965 ;
      RECT 12.465 1.625 12.755 1.855 ;
      RECT 12.465 1.655 14.115 1.825 ;
      RECT 12.525 0.885 12.695 1.855 ;
      RECT 12.465 0.885 12.755 1.115 ;
      RECT 12.465 7.765 12.755 7.995 ;
      RECT 12.525 7.025 12.695 7.995 ;
      RECT 12.525 7.12 14.115 7.29 ;
      RECT 13.945 5.915 14.115 7.29 ;
      RECT 12.465 7.025 12.755 7.255 ;
      RECT 13.89 5.915 14.18 6.145 ;
      RECT 13.89 5.945 14.35 6.115 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 12.725 2.025 13.245 2.195 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 12.895 6.655 13.245 6.885 ;
      RECT 12.725 6.685 13.245 6.855 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 12.09 2.365 12.44 2.595 ;
      RECT 10.56 2.395 12.44 2.565 ;
      RECT 10.56 1.34 10.73 2.565 ;
      RECT 10.46 1.34 10.81 1.69 ;
      RECT 12.12 6.28 12.44 6.605 ;
      RECT 12.09 6.285 12.44 6.515 ;
      RECT 11.92 6.315 12.44 6.485 ;
      RECT 11.065 2.705 11.415 3.055 ;
      RECT 11.065 2.765 11.555 2.935 ;
      RECT 11.07 5.855 11.42 6.205 ;
      RECT 11.07 5.945 11.555 6.115 ;
      RECT 8.755 2.465 8.94 2.675 ;
      RECT 8.745 2.47 8.955 2.668 ;
      RECT 8.745 2.47 9.041 2.645 ;
      RECT 8.745 2.47 9.1 2.62 ;
      RECT 8.745 2.47 9.155 2.6 ;
      RECT 8.745 2.47 9.165 2.588 ;
      RECT 8.745 2.47 9.36 2.527 ;
      RECT 8.745 2.47 9.39 2.51 ;
      RECT 8.745 2.47 9.41 2.5 ;
      RECT 9.29 2.235 9.55 2.495 ;
      RECT 9.275 2.325 9.29 2.542 ;
      RECT 8.81 2.457 9.55 2.495 ;
      RECT 9.261 2.336 9.275 2.548 ;
      RECT 8.85 2.45 9.55 2.495 ;
      RECT 9.175 2.376 9.261 2.567 ;
      RECT 9.1 2.437 9.55 2.495 ;
      RECT 9.17 2.412 9.175 2.584 ;
      RECT 9.155 2.422 9.55 2.495 ;
      RECT 9.165 2.417 9.17 2.586 ;
      RECT 9.46 2.922 9.465 3.014 ;
      RECT 9.455 2.9 9.46 3.031 ;
      RECT 9.45 2.89 9.455 3.043 ;
      RECT 9.44 2.881 9.45 3.053 ;
      RECT 9.435 2.876 9.44 3.061 ;
      RECT 9.43 2.735 9.435 3.064 ;
      RECT 9.396 2.735 9.43 3.075 ;
      RECT 9.31 2.735 9.396 3.11 ;
      RECT 9.23 2.735 9.31 3.158 ;
      RECT 9.201 2.735 9.23 3.182 ;
      RECT 9.115 2.735 9.201 3.188 ;
      RECT 9.11 2.919 9.115 3.193 ;
      RECT 9.075 2.93 9.11 3.196 ;
      RECT 9.05 2.945 9.075 3.2 ;
      RECT 9.036 2.954 9.05 3.202 ;
      RECT 8.95 2.981 9.036 3.208 ;
      RECT 8.885 3.022 8.95 3.217 ;
      RECT 8.87 3.042 8.885 3.222 ;
      RECT 8.84 3.052 8.87 3.225 ;
      RECT 8.835 3.062 8.84 3.228 ;
      RECT 8.805 3.067 8.835 3.23 ;
      RECT 8.785 3.072 8.805 3.234 ;
      RECT 8.7 3.075 8.785 3.241 ;
      RECT 8.685 3.072 8.7 3.247 ;
      RECT 8.675 3.069 8.685 3.249 ;
      RECT 8.655 3.066 8.675 3.251 ;
      RECT 8.635 3.062 8.655 3.252 ;
      RECT 8.62 3.058 8.635 3.254 ;
      RECT 8.61 3.055 8.62 3.255 ;
      RECT 8.57 3.049 8.61 3.253 ;
      RECT 8.56 3.044 8.57 3.251 ;
      RECT 8.545 3.041 8.56 3.247 ;
      RECT 8.52 3.036 8.545 3.24 ;
      RECT 8.47 3.027 8.52 3.228 ;
      RECT 8.4 3.013 8.47 3.21 ;
      RECT 8.342 2.998 8.4 3.192 ;
      RECT 8.256 2.981 8.342 3.172 ;
      RECT 8.17 2.96 8.256 3.147 ;
      RECT 8.12 2.945 8.17 3.128 ;
      RECT 8.116 2.939 8.12 3.12 ;
      RECT 8.03 2.929 8.116 3.107 ;
      RECT 7.995 2.914 8.03 3.09 ;
      RECT 7.98 2.907 7.995 3.083 ;
      RECT 7.92 2.895 7.98 3.071 ;
      RECT 7.9 2.882 7.92 3.059 ;
      RECT 7.86 2.873 7.9 3.051 ;
      RECT 7.855 2.865 7.86 3.044 ;
      RECT 7.775 2.855 7.855 3.03 ;
      RECT 7.76 2.842 7.775 3.015 ;
      RECT 7.755 2.84 7.76 3.013 ;
      RECT 7.676 2.828 7.755 3 ;
      RECT 7.59 2.803 7.676 2.975 ;
      RECT 7.575 2.772 7.59 2.96 ;
      RECT 7.56 2.747 7.575 2.956 ;
      RECT 7.545 2.74 7.56 2.952 ;
      RECT 7.37 2.745 7.375 2.948 ;
      RECT 7.365 2.75 7.37 2.943 ;
      RECT 7.375 2.74 7.545 2.95 ;
      RECT 8.09 2.5 8.195 2.76 ;
      RECT 8.905 2.025 8.91 2.25 ;
      RECT 9.035 2.025 9.09 2.235 ;
      RECT 9.09 2.03 9.1 2.228 ;
      RECT 8.996 2.025 9.035 2.238 ;
      RECT 8.91 2.025 8.996 2.245 ;
      RECT 8.89 2.03 8.905 2.251 ;
      RECT 8.88 2.07 8.89 2.253 ;
      RECT 8.85 2.08 8.88 2.255 ;
      RECT 8.845 2.085 8.85 2.257 ;
      RECT 8.82 2.09 8.845 2.259 ;
      RECT 8.805 2.095 8.82 2.261 ;
      RECT 8.79 2.097 8.805 2.263 ;
      RECT 8.785 2.102 8.79 2.265 ;
      RECT 8.735 2.11 8.785 2.268 ;
      RECT 8.71 2.119 8.735 2.273 ;
      RECT 8.7 2.126 8.71 2.278 ;
      RECT 8.695 2.129 8.7 2.282 ;
      RECT 8.675 2.132 8.695 2.291 ;
      RECT 8.645 2.14 8.675 2.311 ;
      RECT 8.616 2.153 8.645 2.333 ;
      RECT 8.53 2.187 8.616 2.377 ;
      RECT 8.525 2.213 8.53 2.415 ;
      RECT 8.52 2.217 8.525 2.424 ;
      RECT 8.485 2.23 8.52 2.457 ;
      RECT 8.475 2.244 8.485 2.495 ;
      RECT 8.47 2.248 8.475 2.508 ;
      RECT 8.465 2.252 8.47 2.513 ;
      RECT 8.455 2.26 8.465 2.525 ;
      RECT 8.45 2.267 8.455 2.54 ;
      RECT 8.425 2.28 8.45 2.565 ;
      RECT 8.385 2.309 8.425 2.62 ;
      RECT 8.37 2.334 8.385 2.675 ;
      RECT 8.36 2.345 8.37 2.698 ;
      RECT 8.355 2.352 8.36 2.71 ;
      RECT 8.35 2.356 8.355 2.718 ;
      RECT 8.295 2.384 8.35 2.76 ;
      RECT 8.275 2.42 8.295 2.76 ;
      RECT 8.26 2.435 8.275 2.76 ;
      RECT 8.205 2.467 8.26 2.76 ;
      RECT 8.195 2.497 8.205 2.76 ;
      RECT 7.805 2.112 7.99 2.35 ;
      RECT 7.79 2.114 8 2.345 ;
      RECT 7.675 2.06 7.935 2.32 ;
      RECT 7.67 2.097 7.935 2.274 ;
      RECT 7.665 2.107 7.935 2.271 ;
      RECT 7.66 2.147 8 2.265 ;
      RECT 7.655 2.18 8 2.255 ;
      RECT 7.665 2.122 8.015 2.193 ;
      RECT 7.962 3.22 7.975 3.75 ;
      RECT 7.876 3.22 7.975 3.749 ;
      RECT 7.876 3.22 7.98 3.748 ;
      RECT 7.79 3.22 7.98 3.746 ;
      RECT 7.785 3.22 7.98 3.743 ;
      RECT 7.785 3.22 7.99 3.741 ;
      RECT 7.78 3.512 7.99 3.738 ;
      RECT 7.78 3.522 7.995 3.735 ;
      RECT 7.78 3.59 8 3.731 ;
      RECT 7.77 3.595 8 3.73 ;
      RECT 7.77 3.687 8.005 3.727 ;
      RECT 7.755 3.22 8.015 3.48 ;
      RECT 6.985 2.21 7.03 3.745 ;
      RECT 7.185 2.21 7.215 2.425 ;
      RECT 5.56 1.95 5.68 2.16 ;
      RECT 5.22 1.9 5.48 2.16 ;
      RECT 5.22 1.945 5.515 2.15 ;
      RECT 7.225 2.226 7.23 2.28 ;
      RECT 7.22 2.219 7.225 2.413 ;
      RECT 7.215 2.213 7.22 2.42 ;
      RECT 7.17 2.21 7.185 2.433 ;
      RECT 7.165 2.21 7.17 2.455 ;
      RECT 7.16 2.21 7.165 2.503 ;
      RECT 7.155 2.21 7.16 2.523 ;
      RECT 7.145 2.21 7.155 2.63 ;
      RECT 7.14 2.21 7.145 2.693 ;
      RECT 7.135 2.21 7.14 2.75 ;
      RECT 7.13 2.21 7.135 2.758 ;
      RECT 7.115 2.21 7.13 2.865 ;
      RECT 7.105 2.21 7.115 3 ;
      RECT 7.095 2.21 7.105 3.11 ;
      RECT 7.085 2.21 7.095 3.167 ;
      RECT 7.08 2.21 7.085 3.207 ;
      RECT 7.075 2.21 7.08 3.243 ;
      RECT 7.065 2.21 7.075 3.283 ;
      RECT 7.06 2.21 7.065 3.325 ;
      RECT 7.04 2.21 7.06 3.39 ;
      RECT 7.045 3.535 7.05 3.715 ;
      RECT 7.04 3.517 7.045 3.723 ;
      RECT 7.035 2.21 7.04 3.453 ;
      RECT 7.035 3.497 7.04 3.73 ;
      RECT 7.03 2.21 7.035 3.74 ;
      RECT 6.975 2.21 6.985 2.51 ;
      RECT 6.98 2.757 6.985 3.745 ;
      RECT 6.975 2.822 6.98 3.745 ;
      RECT 6.97 2.211 6.975 2.5 ;
      RECT 6.965 2.887 6.975 3.745 ;
      RECT 6.96 2.212 6.97 2.49 ;
      RECT 6.95 3 6.965 3.745 ;
      RECT 6.955 2.213 6.96 2.48 ;
      RECT 6.935 2.214 6.955 2.458 ;
      RECT 6.94 3.097 6.95 3.745 ;
      RECT 6.935 3.172 6.94 3.745 ;
      RECT 6.925 2.213 6.935 2.435 ;
      RECT 6.93 3.215 6.935 3.745 ;
      RECT 6.925 3.242 6.93 3.745 ;
      RECT 6.915 2.211 6.925 2.423 ;
      RECT 6.92 3.285 6.925 3.745 ;
      RECT 6.915 3.312 6.92 3.745 ;
      RECT 6.905 2.21 6.915 2.41 ;
      RECT 6.91 3.327 6.915 3.745 ;
      RECT 6.87 3.385 6.91 3.745 ;
      RECT 6.9 2.209 6.905 2.395 ;
      RECT 6.895 2.207 6.9 2.388 ;
      RECT 6.885 2.204 6.895 2.378 ;
      RECT 6.88 2.201 6.885 2.363 ;
      RECT 6.865 2.197 6.88 2.356 ;
      RECT 6.86 3.44 6.87 3.745 ;
      RECT 6.86 2.194 6.865 2.351 ;
      RECT 6.845 2.19 6.86 2.345 ;
      RECT 6.855 3.457 6.86 3.745 ;
      RECT 6.845 3.52 6.855 3.745 ;
      RECT 6.765 2.175 6.845 2.325 ;
      RECT 6.84 3.527 6.845 3.74 ;
      RECT 6.835 3.535 6.84 3.73 ;
      RECT 6.755 2.161 6.765 2.309 ;
      RECT 6.74 2.157 6.755 2.307 ;
      RECT 6.73 2.152 6.74 2.303 ;
      RECT 6.705 2.145 6.73 2.295 ;
      RECT 6.7 2.14 6.705 2.29 ;
      RECT 6.69 2.14 6.7 2.288 ;
      RECT 6.68 2.138 6.69 2.286 ;
      RECT 6.65 2.13 6.68 2.28 ;
      RECT 6.635 2.122 6.65 2.273 ;
      RECT 6.615 2.117 6.635 2.266 ;
      RECT 6.61 2.113 6.615 2.261 ;
      RECT 6.58 2.106 6.61 2.255 ;
      RECT 6.555 2.097 6.58 2.245 ;
      RECT 6.525 2.09 6.555 2.237 ;
      RECT 6.5 2.08 6.525 2.228 ;
      RECT 6.485 2.072 6.5 2.222 ;
      RECT 6.46 2.067 6.485 2.217 ;
      RECT 6.45 2.063 6.46 2.212 ;
      RECT 6.43 2.058 6.45 2.207 ;
      RECT 6.395 2.053 6.43 2.2 ;
      RECT 6.335 2.048 6.395 2.193 ;
      RECT 6.322 2.044 6.335 2.191 ;
      RECT 6.236 2.039 6.322 2.188 ;
      RECT 6.15 2.029 6.236 2.184 ;
      RECT 6.109 2.022 6.15 2.181 ;
      RECT 6.023 2.015 6.109 2.178 ;
      RECT 5.937 2.005 6.023 2.174 ;
      RECT 5.851 1.995 5.937 2.169 ;
      RECT 5.765 1.985 5.851 2.165 ;
      RECT 5.755 1.97 5.765 2.163 ;
      RECT 5.745 1.955 5.755 2.163 ;
      RECT 5.68 1.95 5.745 2.162 ;
      RECT 5.515 1.947 5.56 2.155 ;
      RECT 6.76 2.852 6.765 3.043 ;
      RECT 6.755 2.847 6.76 3.05 ;
      RECT 6.741 2.845 6.755 3.056 ;
      RECT 6.655 2.845 6.741 3.058 ;
      RECT 6.651 2.845 6.655 3.061 ;
      RECT 6.565 2.845 6.651 3.079 ;
      RECT 6.555 2.85 6.565 3.098 ;
      RECT 6.545 2.905 6.555 3.102 ;
      RECT 6.52 2.92 6.545 3.109 ;
      RECT 6.48 2.94 6.52 3.122 ;
      RECT 6.475 2.952 6.48 3.132 ;
      RECT 6.46 2.958 6.475 3.137 ;
      RECT 6.455 2.963 6.46 3.141 ;
      RECT 6.435 2.97 6.455 3.146 ;
      RECT 6.365 2.995 6.435 3.163 ;
      RECT 6.325 3.023 6.365 3.183 ;
      RECT 6.32 3.033 6.325 3.191 ;
      RECT 6.3 3.04 6.32 3.193 ;
      RECT 6.295 3.047 6.3 3.196 ;
      RECT 6.265 3.055 6.295 3.199 ;
      RECT 6.26 3.06 6.265 3.203 ;
      RECT 6.186 3.064 6.26 3.211 ;
      RECT 6.1 3.073 6.186 3.227 ;
      RECT 6.096 3.078 6.1 3.236 ;
      RECT 6.01 3.083 6.096 3.246 ;
      RECT 5.97 3.091 6.01 3.258 ;
      RECT 5.92 3.097 5.97 3.265 ;
      RECT 5.835 3.106 5.92 3.28 ;
      RECT 5.76 3.117 5.835 3.298 ;
      RECT 5.725 3.124 5.76 3.308 ;
      RECT 5.65 3.132 5.725 3.313 ;
      RECT 5.595 3.141 5.65 3.313 ;
      RECT 5.57 3.146 5.595 3.311 ;
      RECT 5.56 3.149 5.57 3.309 ;
      RECT 5.525 3.151 5.56 3.307 ;
      RECT 5.495 3.153 5.525 3.303 ;
      RECT 5.45 3.152 5.495 3.299 ;
      RECT 5.43 3.147 5.45 3.296 ;
      RECT 5.38 3.132 5.43 3.293 ;
      RECT 5.37 3.117 5.38 3.288 ;
      RECT 5.32 3.102 5.37 3.278 ;
      RECT 5.27 3.077 5.32 3.258 ;
      RECT 5.26 3.062 5.27 3.24 ;
      RECT 5.255 3.06 5.26 3.234 ;
      RECT 5.235 3.055 5.255 3.229 ;
      RECT 5.23 3.047 5.235 3.223 ;
      RECT 5.215 3.041 5.23 3.216 ;
      RECT 5.21 3.036 5.215 3.208 ;
      RECT 5.19 3.031 5.21 3.2 ;
      RECT 5.175 3.024 5.19 3.193 ;
      RECT 5.16 3.018 5.175 3.184 ;
      RECT 5.155 3.012 5.16 3.177 ;
      RECT 5.11 2.987 5.155 3.163 ;
      RECT 5.095 2.957 5.11 3.145 ;
      RECT 5.08 2.94 5.095 3.136 ;
      RECT 5.055 2.92 5.08 3.124 ;
      RECT 5.015 2.89 5.055 3.104 ;
      RECT 5.005 2.86 5.015 3.089 ;
      RECT 4.99 2.85 5.005 3.082 ;
      RECT 4.935 2.815 4.99 3.061 ;
      RECT 4.92 2.778 4.935 3.04 ;
      RECT 4.91 2.765 4.92 3.032 ;
      RECT 4.86 2.735 4.91 3.014 ;
      RECT 4.845 2.665 4.86 2.995 ;
      RECT 4.8 2.665 4.845 2.978 ;
      RECT 4.775 2.665 4.8 2.96 ;
      RECT 4.765 2.665 4.775 2.953 ;
      RECT 4.686 2.665 4.765 2.946 ;
      RECT 4.6 2.665 4.686 2.938 ;
      RECT 4.585 2.697 4.6 2.933 ;
      RECT 4.51 2.707 4.585 2.929 ;
      RECT 4.49 2.717 4.51 2.924 ;
      RECT 4.465 2.717 4.49 2.921 ;
      RECT 4.455 2.707 4.465 2.92 ;
      RECT 4.445 2.68 4.455 2.919 ;
      RECT 4.405 2.675 4.445 2.917 ;
      RECT 4.36 2.675 4.405 2.913 ;
      RECT 4.335 2.675 4.36 2.908 ;
      RECT 4.285 2.675 4.335 2.895 ;
      RECT 4.245 2.68 4.255 2.88 ;
      RECT 4.255 2.675 4.285 2.885 ;
      RECT 6.24 2.455 6.5 2.715 ;
      RECT 6.235 2.477 6.5 2.673 ;
      RECT 5.475 2.305 5.695 2.67 ;
      RECT 5.457 2.392 5.695 2.669 ;
      RECT 5.44 2.397 5.695 2.666 ;
      RECT 5.44 2.397 5.715 2.665 ;
      RECT 5.41 2.407 5.715 2.663 ;
      RECT 5.405 2.422 5.715 2.659 ;
      RECT 5.405 2.422 5.72 2.658 ;
      RECT 5.4 2.48 5.72 2.656 ;
      RECT 5.4 2.48 5.73 2.653 ;
      RECT 5.395 2.545 5.73 2.648 ;
      RECT 5.475 2.305 5.735 2.565 ;
      RECT 4.22 2.135 4.48 2.395 ;
      RECT 4.22 2.178 4.566 2.369 ;
      RECT 4.22 2.178 4.61 2.368 ;
      RECT 4.22 2.178 4.63 2.366 ;
      RECT 4.22 2.178 4.73 2.365 ;
      RECT 4.22 2.178 4.75 2.363 ;
      RECT 4.22 2.178 4.76 2.358 ;
      RECT 4.63 2.145 4.82 2.355 ;
      RECT 4.63 2.147 4.825 2.353 ;
      RECT 4.62 2.152 4.83 2.345 ;
      RECT 4.566 2.176 4.83 2.345 ;
      RECT 4.61 2.17 4.62 2.367 ;
      RECT 4.62 2.15 4.825 2.353 ;
      RECT 3.575 3.21 3.78 3.44 ;
      RECT 3.515 3.16 3.57 3.42 ;
      RECT 3.575 3.16 3.775 3.44 ;
      RECT 4.545 3.475 4.55 3.502 ;
      RECT 4.535 3.385 4.545 3.507 ;
      RECT 4.53 3.307 4.535 3.513 ;
      RECT 4.52 3.297 4.53 3.52 ;
      RECT 4.515 3.287 4.52 3.526 ;
      RECT 4.505 3.282 4.515 3.528 ;
      RECT 4.49 3.274 4.505 3.536 ;
      RECT 4.475 3.265 4.49 3.548 ;
      RECT 4.465 3.257 4.475 3.558 ;
      RECT 4.43 3.175 4.465 3.576 ;
      RECT 4.395 3.175 4.43 3.595 ;
      RECT 4.38 3.175 4.395 3.603 ;
      RECT 4.325 3.175 4.38 3.603 ;
      RECT 4.291 3.175 4.325 3.594 ;
      RECT 4.205 3.175 4.291 3.57 ;
      RECT 4.195 3.235 4.205 3.552 ;
      RECT 4.155 3.237 4.195 3.543 ;
      RECT 4.15 3.239 4.155 3.533 ;
      RECT 4.13 3.241 4.15 3.528 ;
      RECT 4.12 3.244 4.13 3.523 ;
      RECT 4.11 3.245 4.12 3.518 ;
      RECT 4.086 3.246 4.11 3.51 ;
      RECT 4 3.251 4.086 3.488 ;
      RECT 3.945 3.25 4 3.461 ;
      RECT 3.93 3.243 3.945 3.448 ;
      RECT 3.895 3.238 3.93 3.444 ;
      RECT 3.84 3.23 3.895 3.443 ;
      RECT 3.78 3.217 3.84 3.441 ;
      RECT 3.57 3.16 3.575 3.428 ;
      RECT 3.645 2.53 3.83 2.74 ;
      RECT 3.635 2.535 3.845 2.733 ;
      RECT 3.675 2.44 3.935 2.7 ;
      RECT 3.63 2.597 3.935 2.623 ;
      RECT 2.975 2.39 2.98 3.19 ;
      RECT 2.92 2.44 2.95 3.19 ;
      RECT 2.91 2.44 2.915 2.75 ;
      RECT 2.895 2.44 2.9 2.745 ;
      RECT 2.44 2.485 2.455 2.7 ;
      RECT 2.37 2.485 2.455 2.695 ;
      RECT 3.635 2.065 3.705 2.275 ;
      RECT 3.705 2.072 3.715 2.27 ;
      RECT 3.601 2.065 3.635 2.282 ;
      RECT 3.515 2.065 3.601 2.306 ;
      RECT 3.505 2.07 3.515 2.325 ;
      RECT 3.5 2.082 3.505 2.328 ;
      RECT 3.485 2.097 3.5 2.332 ;
      RECT 3.48 2.115 3.485 2.336 ;
      RECT 3.44 2.125 3.48 2.345 ;
      RECT 3.425 2.132 3.44 2.357 ;
      RECT 3.41 2.137 3.425 2.362 ;
      RECT 3.395 2.14 3.41 2.367 ;
      RECT 3.385 2.142 3.395 2.371 ;
      RECT 3.35 2.149 3.385 2.379 ;
      RECT 3.315 2.157 3.35 2.393 ;
      RECT 3.305 2.163 3.315 2.402 ;
      RECT 3.3 2.165 3.305 2.404 ;
      RECT 3.28 2.168 3.3 2.41 ;
      RECT 3.25 2.175 3.28 2.421 ;
      RECT 3.24 2.181 3.25 2.428 ;
      RECT 3.215 2.184 3.24 2.435 ;
      RECT 3.205 2.188 3.215 2.443 ;
      RECT 3.2 2.189 3.205 2.465 ;
      RECT 3.195 2.19 3.2 2.48 ;
      RECT 3.19 2.191 3.195 2.495 ;
      RECT 3.185 2.192 3.19 2.51 ;
      RECT 3.18 2.193 3.185 2.54 ;
      RECT 3.17 2.195 3.18 2.573 ;
      RECT 3.155 2.199 3.17 2.62 ;
      RECT 3.145 2.202 3.155 2.665 ;
      RECT 3.14 2.205 3.145 2.693 ;
      RECT 3.13 2.207 3.14 2.72 ;
      RECT 3.125 2.21 3.13 2.755 ;
      RECT 3.095 2.215 3.125 2.813 ;
      RECT 3.09 2.22 3.095 2.898 ;
      RECT 3.085 2.222 3.09 2.933 ;
      RECT 3.08 2.224 3.085 3.015 ;
      RECT 3.075 2.226 3.08 3.103 ;
      RECT 3.065 2.228 3.075 3.185 ;
      RECT 3.05 2.242 3.065 3.19 ;
      RECT 3.015 2.287 3.05 3.19 ;
      RECT 3.005 2.327 3.015 3.19 ;
      RECT 2.99 2.355 3.005 3.19 ;
      RECT 2.985 2.372 2.99 3.19 ;
      RECT 2.98 2.38 2.985 3.19 ;
      RECT 2.97 2.395 2.975 3.19 ;
      RECT 2.965 2.402 2.97 3.19 ;
      RECT 2.955 2.422 2.965 3.19 ;
      RECT 2.95 2.435 2.955 3.19 ;
      RECT 2.915 2.44 2.92 2.775 ;
      RECT 2.9 2.83 2.92 3.19 ;
      RECT 2.9 2.44 2.91 2.748 ;
      RECT 2.895 2.87 2.9 3.19 ;
      RECT 2.845 2.44 2.895 2.743 ;
      RECT 2.89 2.907 2.895 3.19 ;
      RECT 2.88 2.93 2.89 3.19 ;
      RECT 2.875 2.975 2.88 3.19 ;
      RECT 2.865 2.985 2.875 3.183 ;
      RECT 2.791 2.44 2.845 2.737 ;
      RECT 2.705 2.44 2.791 2.73 ;
      RECT 2.656 2.487 2.705 2.723 ;
      RECT 2.57 2.495 2.656 2.716 ;
      RECT 2.555 2.492 2.57 2.711 ;
      RECT 2.541 2.485 2.555 2.71 ;
      RECT 2.455 2.485 2.541 2.705 ;
      RECT 2.36 2.49 2.37 2.69 ;
      RECT 1.95 1.92 1.965 2.32 ;
      RECT 2.145 1.92 2.15 2.18 ;
      RECT 1.89 1.92 1.935 2.18 ;
      RECT 2.345 3.225 2.35 3.43 ;
      RECT 2.34 3.215 2.345 3.435 ;
      RECT 2.335 3.202 2.34 3.44 ;
      RECT 2.33 3.182 2.335 3.44 ;
      RECT 2.305 3.135 2.33 3.44 ;
      RECT 2.27 3.05 2.305 3.44 ;
      RECT 2.265 2.987 2.27 3.44 ;
      RECT 2.26 2.972 2.265 3.44 ;
      RECT 2.245 2.932 2.26 3.44 ;
      RECT 2.24 2.907 2.245 3.44 ;
      RECT 2.23 2.89 2.24 3.44 ;
      RECT 2.195 2.812 2.23 3.44 ;
      RECT 2.19 2.755 2.195 3.44 ;
      RECT 2.185 2.742 2.19 3.44 ;
      RECT 2.175 2.72 2.185 3.44 ;
      RECT 2.165 2.685 2.175 3.44 ;
      RECT 2.155 2.655 2.165 3.44 ;
      RECT 2.145 2.57 2.155 3.083 ;
      RECT 2.152 3.215 2.155 3.44 ;
      RECT 2.15 3.225 2.152 3.44 ;
      RECT 2.14 3.235 2.15 3.435 ;
      RECT 2.135 1.92 2.145 2.315 ;
      RECT 2.14 2.447 2.145 3.058 ;
      RECT 2.135 2.345 2.14 3.041 ;
      RECT 2.125 1.92 2.135 3.017 ;
      RECT 2.12 1.92 2.125 2.988 ;
      RECT 2.115 1.92 2.12 2.978 ;
      RECT 2.095 1.92 2.115 2.94 ;
      RECT 2.09 1.92 2.095 2.898 ;
      RECT 2.085 1.92 2.09 2.878 ;
      RECT 2.055 1.92 2.085 2.828 ;
      RECT 2.045 1.92 2.055 2.775 ;
      RECT 2.04 1.92 2.045 2.748 ;
      RECT 2.035 1.92 2.04 2.733 ;
      RECT 2.025 1.92 2.035 2.71 ;
      RECT 2.015 1.92 2.025 2.685 ;
      RECT 2.01 1.92 2.015 2.625 ;
      RECT 2 1.92 2.01 2.563 ;
      RECT 1.995 1.92 2 2.483 ;
      RECT 1.99 1.92 1.995 2.448 ;
      RECT 1.985 1.92 1.99 2.423 ;
      RECT 1.98 1.92 1.985 2.408 ;
      RECT 1.975 1.92 1.98 2.378 ;
      RECT 1.97 1.92 1.975 2.355 ;
      RECT 1.965 1.92 1.97 2.328 ;
      RECT 1.935 1.92 1.95 2.315 ;
      RECT 1.09 3.455 1.275 3.665 ;
      RECT 1.08 3.46 1.29 3.658 ;
      RECT 1.08 3.46 1.31 3.63 ;
      RECT 1.08 3.46 1.325 3.609 ;
      RECT 1.08 3.46 1.34 3.607 ;
      RECT 1.08 3.46 1.35 3.606 ;
      RECT 1.08 3.46 1.38 3.603 ;
      RECT 1.73 3.305 1.99 3.565 ;
      RECT 1.69 3.352 1.99 3.548 ;
      RECT 1.681 3.36 1.69 3.551 ;
      RECT 1.275 3.453 1.99 3.548 ;
      RECT 1.595 3.378 1.681 3.558 ;
      RECT 1.29 3.45 1.99 3.548 ;
      RECT 1.536 3.4 1.595 3.57 ;
      RECT 1.31 3.446 1.99 3.548 ;
      RECT 1.45 3.412 1.536 3.581 ;
      RECT 1.325 3.442 1.99 3.548 ;
      RECT 1.395 3.425 1.45 3.593 ;
      RECT 1.34 3.44 1.99 3.548 ;
      RECT 1.38 3.431 1.395 3.599 ;
      RECT 1.35 3.436 1.99 3.548 ;
      RECT 1.495 2.96 1.755 3.22 ;
      RECT 1.495 2.98 1.865 3.19 ;
      RECT 1.495 2.985 1.875 3.185 ;
      RECT 1.686 2.399 1.765 2.63 ;
      RECT 1.6 2.402 1.815 2.625 ;
      RECT 1.595 2.402 1.815 2.62 ;
      RECT 1.595 2.407 1.825 2.618 ;
      RECT 1.57 2.407 1.825 2.615 ;
      RECT 1.57 2.415 1.835 2.613 ;
      RECT 1.45 2.35 1.71 2.61 ;
      RECT 1.45 2.397 1.76 2.61 ;
      RECT 0.705 2.97 0.71 3.23 ;
      RECT 0.535 2.74 0.54 3.23 ;
      RECT 0.42 2.98 0.425 3.205 ;
      RECT 1.13 2.075 1.135 2.285 ;
      RECT 1.135 2.08 1.15 2.28 ;
      RECT 1.07 2.075 1.13 2.293 ;
      RECT 1.055 2.075 1.07 2.303 ;
      RECT 1.005 2.075 1.055 2.32 ;
      RECT 0.985 2.075 1.005 2.343 ;
      RECT 0.97 2.075 0.985 2.355 ;
      RECT 0.95 2.075 0.97 2.365 ;
      RECT 0.94 2.08 0.95 2.374 ;
      RECT 0.935 2.09 0.94 2.379 ;
      RECT 0.93 2.102 0.935 2.383 ;
      RECT 0.92 2.125 0.93 2.388 ;
      RECT 0.915 2.14 0.92 2.392 ;
      RECT 0.91 2.157 0.915 2.395 ;
      RECT 0.905 2.165 0.91 2.398 ;
      RECT 0.895 2.17 0.905 2.402 ;
      RECT 0.89 2.177 0.895 2.407 ;
      RECT 0.88 2.182 0.89 2.411 ;
      RECT 0.855 2.194 0.88 2.422 ;
      RECT 0.835 2.211 0.855 2.438 ;
      RECT 0.81 2.228 0.835 2.46 ;
      RECT 0.775 2.251 0.81 2.518 ;
      RECT 0.755 2.273 0.775 2.58 ;
      RECT 0.75 2.283 0.755 2.615 ;
      RECT 0.74 2.29 0.75 2.653 ;
      RECT 0.735 2.297 0.74 2.673 ;
      RECT 0.73 2.308 0.735 2.71 ;
      RECT 0.725 2.316 0.73 2.775 ;
      RECT 0.715 2.327 0.725 2.828 ;
      RECT 0.71 2.345 0.715 2.898 ;
      RECT 0.705 2.355 0.71 2.935 ;
      RECT 0.7 2.365 0.705 3.23 ;
      RECT 0.695 2.377 0.7 3.23 ;
      RECT 0.69 2.387 0.695 3.23 ;
      RECT 0.68 2.397 0.69 3.23 ;
      RECT 0.67 2.42 0.68 3.23 ;
      RECT 0.655 2.455 0.67 3.23 ;
      RECT 0.615 2.517 0.655 3.23 ;
      RECT 0.61 2.57 0.615 3.23 ;
      RECT 0.585 2.605 0.61 3.23 ;
      RECT 0.57 2.65 0.585 3.23 ;
      RECT 0.565 2.672 0.57 3.23 ;
      RECT 0.555 2.685 0.565 3.23 ;
      RECT 0.545 2.71 0.555 3.23 ;
      RECT 0.54 2.732 0.545 3.23 ;
      RECT 0.515 2.77 0.535 3.23 ;
      RECT 0.475 2.827 0.515 3.23 ;
      RECT 0.47 2.877 0.475 3.23 ;
      RECT 0.465 2.895 0.47 3.23 ;
      RECT 0.46 2.907 0.465 3.23 ;
      RECT 0.45 2.925 0.46 3.23 ;
      RECT 0.44 2.945 0.45 3.205 ;
      RECT 0.435 2.962 0.44 3.205 ;
      RECT 0.425 2.975 0.435 3.205 ;
      RECT 0.395 2.985 0.42 3.205 ;
      RECT 0.385 2.992 0.395 3.205 ;
      RECT 0.37 3.002 0.385 3.2 ;
      RECT 0 8.575 79.25 8.88 ;
    LAYER mcon ;
      RECT 78.71 2.395 78.88 2.565 ;
      RECT 78.715 2.225 78.885 2.395 ;
      RECT 78.71 0.915 78.88 1.085 ;
      RECT 78.71 6.315 78.88 6.485 ;
      RECT 78.71 7.795 78.88 7.965 ;
      RECT 78.36 0.105 78.53 0.275 ;
      RECT 78.36 4.165 78.53 4.335 ;
      RECT 78.36 4.545 78.53 4.715 ;
      RECT 78.36 8.605 78.53 8.775 ;
      RECT 78.34 2.765 78.51 2.935 ;
      RECT 78.34 5.945 78.51 6.115 ;
      RECT 77.72 0.915 77.89 1.085 ;
      RECT 77.72 2.395 77.89 2.565 ;
      RECT 77.72 6.315 77.89 6.485 ;
      RECT 77.72 7.795 77.89 7.965 ;
      RECT 77.37 0.105 77.54 0.275 ;
      RECT 77.37 4.165 77.54 4.335 ;
      RECT 77.37 4.545 77.54 4.715 ;
      RECT 77.37 8.605 77.54 8.775 ;
      RECT 77.35 2.765 77.52 2.935 ;
      RECT 77.35 5.945 77.52 6.115 ;
      RECT 76.665 0.105 76.835 0.275 ;
      RECT 76.665 4.165 76.835 4.335 ;
      RECT 76.665 4.545 76.835 4.715 ;
      RECT 76.665 8.605 76.835 8.775 ;
      RECT 76.355 2.025 76.525 2.195 ;
      RECT 76.355 6.685 76.525 6.855 ;
      RECT 75.985 0.105 76.155 0.275 ;
      RECT 75.985 8.605 76.155 8.775 ;
      RECT 75.925 0.915 76.095 1.085 ;
      RECT 75.925 1.655 76.095 1.825 ;
      RECT 75.925 7.055 76.095 7.225 ;
      RECT 75.925 7.795 76.095 7.965 ;
      RECT 75.55 2.395 75.72 2.565 ;
      RECT 75.55 6.315 75.72 6.485 ;
      RECT 75.305 0.105 75.475 0.275 ;
      RECT 75.305 8.605 75.475 8.775 ;
      RECT 74.625 0.105 74.795 0.275 ;
      RECT 74.625 8.605 74.795 8.775 ;
      RECT 74.555 2.765 74.725 2.935 ;
      RECT 74.555 5.945 74.725 6.115 ;
      RECT 73 1.415 73.17 1.585 ;
      RECT 73 4.135 73.17 4.305 ;
      RECT 72.63 2.875 72.8 3.045 ;
      RECT 72.54 1.415 72.71 1.585 ;
      RECT 72.54 4.135 72.71 4.305 ;
      RECT 72.31 2.045 72.48 2.215 ;
      RECT 72.165 2.485 72.335 2.655 ;
      RECT 72.08 1.415 72.25 1.585 ;
      RECT 72.08 4.135 72.25 4.305 ;
      RECT 71.62 1.415 71.79 1.585 ;
      RECT 71.62 4.135 71.79 4.305 ;
      RECT 71.555 2.525 71.725 2.695 ;
      RECT 71.21 2.16 71.38 2.33 ;
      RECT 71.2 3.52 71.37 3.69 ;
      RECT 71.16 1.415 71.33 1.585 ;
      RECT 71.16 4.135 71.33 4.305 ;
      RECT 70.785 2.76 70.955 2.93 ;
      RECT 70.7 1.415 70.87 1.585 ;
      RECT 70.7 4.135 70.87 4.305 ;
      RECT 70.435 2.235 70.605 2.405 ;
      RECT 70.255 3.55 70.425 3.72 ;
      RECT 70.24 1.415 70.41 1.585 ;
      RECT 70.24 4.135 70.41 4.305 ;
      RECT 69.975 2.865 70.145 3.035 ;
      RECT 69.78 1.415 69.95 1.585 ;
      RECT 69.78 4.135 69.95 4.305 ;
      RECT 69.655 2.49 69.825 2.66 ;
      RECT 69.32 1.415 69.49 1.585 ;
      RECT 69.32 4.135 69.49 4.305 ;
      RECT 68.965 1.97 69.135 2.14 ;
      RECT 68.89 2.44 69.06 2.61 ;
      RECT 68.86 1.415 69.03 1.585 ;
      RECT 68.86 4.135 69.03 4.305 ;
      RECT 68.4 1.415 68.57 1.585 ;
      RECT 68.4 4.135 68.57 4.305 ;
      RECT 68.04 2.165 68.21 2.335 ;
      RECT 67.94 1.415 68.11 1.585 ;
      RECT 67.94 4.135 68.11 4.305 ;
      RECT 67.7 3.36 67.87 3.53 ;
      RECT 67.665 2.695 67.835 2.865 ;
      RECT 67.48 1.415 67.65 1.585 ;
      RECT 67.48 4.135 67.65 4.305 ;
      RECT 67.055 2.55 67.225 2.72 ;
      RECT 67.02 1.415 67.19 1.585 ;
      RECT 67.02 4.135 67.19 4.305 ;
      RECT 66.985 3.25 67.155 3.42 ;
      RECT 66.925 2.085 67.095 2.255 ;
      RECT 66.56 1.415 66.73 1.585 ;
      RECT 66.56 4.135 66.73 4.305 ;
      RECT 66.285 3 66.455 3.17 ;
      RECT 66.1 1.415 66.27 1.585 ;
      RECT 66.1 4.135 66.27 4.305 ;
      RECT 65.78 2.505 65.95 2.675 ;
      RECT 65.64 1.415 65.81 1.585 ;
      RECT 65.64 4.135 65.81 4.305 ;
      RECT 65.56 3.25 65.73 3.42 ;
      RECT 65.355 2.13 65.525 2.3 ;
      RECT 65.18 1.415 65.35 1.585 ;
      RECT 65.18 4.135 65.35 4.305 ;
      RECT 65.085 3 65.255 3.17 ;
      RECT 65.045 2.43 65.215 2.6 ;
      RECT 64.72 1.415 64.89 1.585 ;
      RECT 64.72 4.135 64.89 4.305 ;
      RECT 64.5 3.475 64.67 3.645 ;
      RECT 64.36 2.095 64.53 2.265 ;
      RECT 64.26 1.415 64.43 1.585 ;
      RECT 64.26 4.135 64.43 4.305 ;
      RECT 63.8 1.415 63.97 1.585 ;
      RECT 63.8 4.135 63.97 4.305 ;
      RECT 63.79 3.015 63.96 3.185 ;
      RECT 62.86 0.915 63.03 1.085 ;
      RECT 62.86 2.395 63.03 2.565 ;
      RECT 62.86 6.315 63.03 6.485 ;
      RECT 62.86 7.795 63.03 7.965 ;
      RECT 62.51 0.105 62.68 0.275 ;
      RECT 62.51 4.165 62.68 4.335 ;
      RECT 62.51 4.545 62.68 4.715 ;
      RECT 62.51 8.605 62.68 8.775 ;
      RECT 62.49 2.765 62.66 2.935 ;
      RECT 62.49 5.945 62.66 6.115 ;
      RECT 61.87 0.915 62.04 1.085 ;
      RECT 61.87 2.395 62.04 2.565 ;
      RECT 61.87 6.315 62.04 6.485 ;
      RECT 61.87 7.795 62.04 7.965 ;
      RECT 61.52 0.105 61.69 0.275 ;
      RECT 61.52 4.165 61.69 4.335 ;
      RECT 61.52 4.545 61.69 4.715 ;
      RECT 61.52 8.605 61.69 8.775 ;
      RECT 61.5 2.765 61.67 2.935 ;
      RECT 61.5 5.945 61.67 6.115 ;
      RECT 60.815 0.105 60.985 0.275 ;
      RECT 60.815 4.165 60.985 4.335 ;
      RECT 60.815 4.545 60.985 4.715 ;
      RECT 60.815 8.605 60.985 8.775 ;
      RECT 60.505 2.025 60.675 2.195 ;
      RECT 60.505 6.685 60.675 6.855 ;
      RECT 60.135 0.105 60.305 0.275 ;
      RECT 60.135 8.605 60.305 8.775 ;
      RECT 60.075 0.915 60.245 1.085 ;
      RECT 60.075 1.655 60.245 1.825 ;
      RECT 60.075 7.055 60.245 7.225 ;
      RECT 60.075 7.795 60.245 7.965 ;
      RECT 59.7 2.395 59.87 2.565 ;
      RECT 59.7 6.315 59.87 6.485 ;
      RECT 59.455 0.105 59.625 0.275 ;
      RECT 59.455 8.605 59.625 8.775 ;
      RECT 58.775 0.105 58.945 0.275 ;
      RECT 58.775 8.605 58.945 8.775 ;
      RECT 58.705 2.765 58.875 2.935 ;
      RECT 58.705 5.945 58.875 6.115 ;
      RECT 57.15 1.415 57.32 1.585 ;
      RECT 57.15 4.135 57.32 4.305 ;
      RECT 56.78 2.875 56.95 3.045 ;
      RECT 56.69 1.415 56.86 1.585 ;
      RECT 56.69 4.135 56.86 4.305 ;
      RECT 56.46 2.045 56.63 2.215 ;
      RECT 56.315 2.485 56.485 2.655 ;
      RECT 56.23 1.415 56.4 1.585 ;
      RECT 56.23 4.135 56.4 4.305 ;
      RECT 55.77 1.415 55.94 1.585 ;
      RECT 55.77 4.135 55.94 4.305 ;
      RECT 55.705 2.525 55.875 2.695 ;
      RECT 55.36 2.16 55.53 2.33 ;
      RECT 55.35 3.52 55.52 3.69 ;
      RECT 55.31 1.415 55.48 1.585 ;
      RECT 55.31 4.135 55.48 4.305 ;
      RECT 54.935 2.76 55.105 2.93 ;
      RECT 54.85 1.415 55.02 1.585 ;
      RECT 54.85 4.135 55.02 4.305 ;
      RECT 54.585 2.235 54.755 2.405 ;
      RECT 54.405 3.55 54.575 3.72 ;
      RECT 54.39 1.415 54.56 1.585 ;
      RECT 54.39 4.135 54.56 4.305 ;
      RECT 54.125 2.865 54.295 3.035 ;
      RECT 53.93 1.415 54.1 1.585 ;
      RECT 53.93 4.135 54.1 4.305 ;
      RECT 53.805 2.49 53.975 2.66 ;
      RECT 53.47 1.415 53.64 1.585 ;
      RECT 53.47 4.135 53.64 4.305 ;
      RECT 53.115 1.97 53.285 2.14 ;
      RECT 53.04 2.44 53.21 2.61 ;
      RECT 53.01 1.415 53.18 1.585 ;
      RECT 53.01 4.135 53.18 4.305 ;
      RECT 52.55 1.415 52.72 1.585 ;
      RECT 52.55 4.135 52.72 4.305 ;
      RECT 52.19 2.165 52.36 2.335 ;
      RECT 52.09 1.415 52.26 1.585 ;
      RECT 52.09 4.135 52.26 4.305 ;
      RECT 51.85 3.36 52.02 3.53 ;
      RECT 51.815 2.695 51.985 2.865 ;
      RECT 51.63 1.415 51.8 1.585 ;
      RECT 51.63 4.135 51.8 4.305 ;
      RECT 51.205 2.55 51.375 2.72 ;
      RECT 51.17 1.415 51.34 1.585 ;
      RECT 51.17 4.135 51.34 4.305 ;
      RECT 51.135 3.25 51.305 3.42 ;
      RECT 51.075 2.085 51.245 2.255 ;
      RECT 50.71 1.415 50.88 1.585 ;
      RECT 50.71 4.135 50.88 4.305 ;
      RECT 50.435 3 50.605 3.17 ;
      RECT 50.25 1.415 50.42 1.585 ;
      RECT 50.25 4.135 50.42 4.305 ;
      RECT 49.93 2.505 50.1 2.675 ;
      RECT 49.79 1.415 49.96 1.585 ;
      RECT 49.79 4.135 49.96 4.305 ;
      RECT 49.71 3.25 49.88 3.42 ;
      RECT 49.505 2.13 49.675 2.3 ;
      RECT 49.33 1.415 49.5 1.585 ;
      RECT 49.33 4.135 49.5 4.305 ;
      RECT 49.235 3 49.405 3.17 ;
      RECT 49.195 2.43 49.365 2.6 ;
      RECT 48.87 1.415 49.04 1.585 ;
      RECT 48.87 4.135 49.04 4.305 ;
      RECT 48.65 3.475 48.82 3.645 ;
      RECT 48.51 2.095 48.68 2.265 ;
      RECT 48.41 1.415 48.58 1.585 ;
      RECT 48.41 4.135 48.58 4.305 ;
      RECT 47.95 1.415 48.12 1.585 ;
      RECT 47.95 4.135 48.12 4.305 ;
      RECT 47.94 3.015 48.11 3.185 ;
      RECT 47.01 0.915 47.18 1.085 ;
      RECT 47.01 2.395 47.18 2.565 ;
      RECT 47.01 6.315 47.18 6.485 ;
      RECT 47.01 7.795 47.18 7.965 ;
      RECT 46.66 0.105 46.83 0.275 ;
      RECT 46.66 4.165 46.83 4.335 ;
      RECT 46.66 4.545 46.83 4.715 ;
      RECT 46.66 8.605 46.83 8.775 ;
      RECT 46.64 2.765 46.81 2.935 ;
      RECT 46.64 5.945 46.81 6.115 ;
      RECT 46.02 0.915 46.19 1.085 ;
      RECT 46.02 2.395 46.19 2.565 ;
      RECT 46.02 6.315 46.19 6.485 ;
      RECT 46.02 7.795 46.19 7.965 ;
      RECT 45.67 0.105 45.84 0.275 ;
      RECT 45.67 4.165 45.84 4.335 ;
      RECT 45.67 4.545 45.84 4.715 ;
      RECT 45.67 8.605 45.84 8.775 ;
      RECT 45.65 2.765 45.82 2.935 ;
      RECT 45.65 5.945 45.82 6.115 ;
      RECT 44.965 0.105 45.135 0.275 ;
      RECT 44.965 4.165 45.135 4.335 ;
      RECT 44.965 4.545 45.135 4.715 ;
      RECT 44.965 8.605 45.135 8.775 ;
      RECT 44.655 2.025 44.825 2.195 ;
      RECT 44.655 6.685 44.825 6.855 ;
      RECT 44.285 0.105 44.455 0.275 ;
      RECT 44.285 8.605 44.455 8.775 ;
      RECT 44.225 0.915 44.395 1.085 ;
      RECT 44.225 1.655 44.395 1.825 ;
      RECT 44.225 7.055 44.395 7.225 ;
      RECT 44.225 7.795 44.395 7.965 ;
      RECT 43.85 2.395 44.02 2.565 ;
      RECT 43.85 6.315 44.02 6.485 ;
      RECT 43.605 0.105 43.775 0.275 ;
      RECT 43.605 8.605 43.775 8.775 ;
      RECT 42.925 0.105 43.095 0.275 ;
      RECT 42.925 8.605 43.095 8.775 ;
      RECT 42.855 2.765 43.025 2.935 ;
      RECT 42.855 5.945 43.025 6.115 ;
      RECT 41.3 1.415 41.47 1.585 ;
      RECT 41.3 4.135 41.47 4.305 ;
      RECT 40.93 2.875 41.1 3.045 ;
      RECT 40.84 1.415 41.01 1.585 ;
      RECT 40.84 4.135 41.01 4.305 ;
      RECT 40.61 2.045 40.78 2.215 ;
      RECT 40.465 2.485 40.635 2.655 ;
      RECT 40.38 1.415 40.55 1.585 ;
      RECT 40.38 4.135 40.55 4.305 ;
      RECT 39.92 1.415 40.09 1.585 ;
      RECT 39.92 4.135 40.09 4.305 ;
      RECT 39.855 2.525 40.025 2.695 ;
      RECT 39.51 2.16 39.68 2.33 ;
      RECT 39.5 3.52 39.67 3.69 ;
      RECT 39.46 1.415 39.63 1.585 ;
      RECT 39.46 4.135 39.63 4.305 ;
      RECT 39.085 2.76 39.255 2.93 ;
      RECT 39 1.415 39.17 1.585 ;
      RECT 39 4.135 39.17 4.305 ;
      RECT 38.735 2.235 38.905 2.405 ;
      RECT 38.555 3.55 38.725 3.72 ;
      RECT 38.54 1.415 38.71 1.585 ;
      RECT 38.54 4.135 38.71 4.305 ;
      RECT 38.275 2.865 38.445 3.035 ;
      RECT 38.08 1.415 38.25 1.585 ;
      RECT 38.08 4.135 38.25 4.305 ;
      RECT 37.955 2.49 38.125 2.66 ;
      RECT 37.62 1.415 37.79 1.585 ;
      RECT 37.62 4.135 37.79 4.305 ;
      RECT 37.265 1.97 37.435 2.14 ;
      RECT 37.19 2.44 37.36 2.61 ;
      RECT 37.16 1.415 37.33 1.585 ;
      RECT 37.16 4.135 37.33 4.305 ;
      RECT 36.7 1.415 36.87 1.585 ;
      RECT 36.7 4.135 36.87 4.305 ;
      RECT 36.34 2.165 36.51 2.335 ;
      RECT 36.24 1.415 36.41 1.585 ;
      RECT 36.24 4.135 36.41 4.305 ;
      RECT 36 3.36 36.17 3.53 ;
      RECT 35.965 2.695 36.135 2.865 ;
      RECT 35.78 1.415 35.95 1.585 ;
      RECT 35.78 4.135 35.95 4.305 ;
      RECT 35.355 2.55 35.525 2.72 ;
      RECT 35.32 1.415 35.49 1.585 ;
      RECT 35.32 4.135 35.49 4.305 ;
      RECT 35.285 3.25 35.455 3.42 ;
      RECT 35.225 2.085 35.395 2.255 ;
      RECT 34.86 1.415 35.03 1.585 ;
      RECT 34.86 4.135 35.03 4.305 ;
      RECT 34.585 3 34.755 3.17 ;
      RECT 34.4 1.415 34.57 1.585 ;
      RECT 34.4 4.135 34.57 4.305 ;
      RECT 34.08 2.505 34.25 2.675 ;
      RECT 33.94 1.415 34.11 1.585 ;
      RECT 33.94 4.135 34.11 4.305 ;
      RECT 33.86 3.25 34.03 3.42 ;
      RECT 33.655 2.13 33.825 2.3 ;
      RECT 33.48 1.415 33.65 1.585 ;
      RECT 33.48 4.135 33.65 4.305 ;
      RECT 33.385 3 33.555 3.17 ;
      RECT 33.345 2.43 33.515 2.6 ;
      RECT 33.02 1.415 33.19 1.585 ;
      RECT 33.02 4.135 33.19 4.305 ;
      RECT 32.8 3.475 32.97 3.645 ;
      RECT 32.66 2.095 32.83 2.265 ;
      RECT 32.56 1.415 32.73 1.585 ;
      RECT 32.56 4.135 32.73 4.305 ;
      RECT 32.1 1.415 32.27 1.585 ;
      RECT 32.1 4.135 32.27 4.305 ;
      RECT 32.09 3.015 32.26 3.185 ;
      RECT 31.16 0.915 31.33 1.085 ;
      RECT 31.16 2.395 31.33 2.565 ;
      RECT 31.16 6.315 31.33 6.485 ;
      RECT 31.16 7.795 31.33 7.965 ;
      RECT 30.81 0.105 30.98 0.275 ;
      RECT 30.81 4.165 30.98 4.335 ;
      RECT 30.81 4.545 30.98 4.715 ;
      RECT 30.81 8.605 30.98 8.775 ;
      RECT 30.79 2.765 30.96 2.935 ;
      RECT 30.79 5.945 30.96 6.115 ;
      RECT 30.17 0.915 30.34 1.085 ;
      RECT 30.17 2.395 30.34 2.565 ;
      RECT 30.17 6.315 30.34 6.485 ;
      RECT 30.17 7.795 30.34 7.965 ;
      RECT 29.82 0.105 29.99 0.275 ;
      RECT 29.82 4.165 29.99 4.335 ;
      RECT 29.82 4.545 29.99 4.715 ;
      RECT 29.82 8.605 29.99 8.775 ;
      RECT 29.8 2.765 29.97 2.935 ;
      RECT 29.8 5.945 29.97 6.115 ;
      RECT 29.115 0.105 29.285 0.275 ;
      RECT 29.115 4.165 29.285 4.335 ;
      RECT 29.115 4.545 29.285 4.715 ;
      RECT 29.115 8.605 29.285 8.775 ;
      RECT 28.805 2.025 28.975 2.195 ;
      RECT 28.805 6.685 28.975 6.855 ;
      RECT 28.435 0.105 28.605 0.275 ;
      RECT 28.435 8.605 28.605 8.775 ;
      RECT 28.375 0.915 28.545 1.085 ;
      RECT 28.375 1.655 28.545 1.825 ;
      RECT 28.375 7.055 28.545 7.225 ;
      RECT 28.375 7.795 28.545 7.965 ;
      RECT 28 2.395 28.17 2.565 ;
      RECT 28 6.315 28.17 6.485 ;
      RECT 27.755 0.105 27.925 0.275 ;
      RECT 27.755 8.605 27.925 8.775 ;
      RECT 27.075 0.105 27.245 0.275 ;
      RECT 27.075 8.605 27.245 8.775 ;
      RECT 27.005 2.765 27.175 2.935 ;
      RECT 27.005 5.945 27.175 6.115 ;
      RECT 25.45 1.415 25.62 1.585 ;
      RECT 25.45 4.135 25.62 4.305 ;
      RECT 25.08 2.875 25.25 3.045 ;
      RECT 24.99 1.415 25.16 1.585 ;
      RECT 24.99 4.135 25.16 4.305 ;
      RECT 24.76 2.045 24.93 2.215 ;
      RECT 24.615 2.485 24.785 2.655 ;
      RECT 24.53 1.415 24.7 1.585 ;
      RECT 24.53 4.135 24.7 4.305 ;
      RECT 24.07 1.415 24.24 1.585 ;
      RECT 24.07 4.135 24.24 4.305 ;
      RECT 24.005 2.525 24.175 2.695 ;
      RECT 23.66 2.16 23.83 2.33 ;
      RECT 23.65 3.52 23.82 3.69 ;
      RECT 23.61 1.415 23.78 1.585 ;
      RECT 23.61 4.135 23.78 4.305 ;
      RECT 23.235 2.76 23.405 2.93 ;
      RECT 23.15 1.415 23.32 1.585 ;
      RECT 23.15 4.135 23.32 4.305 ;
      RECT 22.885 2.235 23.055 2.405 ;
      RECT 22.705 3.55 22.875 3.72 ;
      RECT 22.69 1.415 22.86 1.585 ;
      RECT 22.69 4.135 22.86 4.305 ;
      RECT 22.425 2.865 22.595 3.035 ;
      RECT 22.23 1.415 22.4 1.585 ;
      RECT 22.23 4.135 22.4 4.305 ;
      RECT 22.105 2.49 22.275 2.66 ;
      RECT 21.77 1.415 21.94 1.585 ;
      RECT 21.77 4.135 21.94 4.305 ;
      RECT 21.415 1.97 21.585 2.14 ;
      RECT 21.34 2.44 21.51 2.61 ;
      RECT 21.31 1.415 21.48 1.585 ;
      RECT 21.31 4.135 21.48 4.305 ;
      RECT 20.85 1.415 21.02 1.585 ;
      RECT 20.85 4.135 21.02 4.305 ;
      RECT 20.49 2.165 20.66 2.335 ;
      RECT 20.39 1.415 20.56 1.585 ;
      RECT 20.39 4.135 20.56 4.305 ;
      RECT 20.15 3.36 20.32 3.53 ;
      RECT 20.115 2.695 20.285 2.865 ;
      RECT 19.93 1.415 20.1 1.585 ;
      RECT 19.93 4.135 20.1 4.305 ;
      RECT 19.505 2.55 19.675 2.72 ;
      RECT 19.47 1.415 19.64 1.585 ;
      RECT 19.47 4.135 19.64 4.305 ;
      RECT 19.435 3.25 19.605 3.42 ;
      RECT 19.375 2.085 19.545 2.255 ;
      RECT 19.01 1.415 19.18 1.585 ;
      RECT 19.01 4.135 19.18 4.305 ;
      RECT 18.735 3 18.905 3.17 ;
      RECT 18.55 1.415 18.72 1.585 ;
      RECT 18.55 4.135 18.72 4.305 ;
      RECT 18.23 2.505 18.4 2.675 ;
      RECT 18.09 1.415 18.26 1.585 ;
      RECT 18.09 4.135 18.26 4.305 ;
      RECT 18.01 3.25 18.18 3.42 ;
      RECT 17.805 2.13 17.975 2.3 ;
      RECT 17.63 1.415 17.8 1.585 ;
      RECT 17.63 4.135 17.8 4.305 ;
      RECT 17.535 3 17.705 3.17 ;
      RECT 17.495 2.43 17.665 2.6 ;
      RECT 17.17 1.415 17.34 1.585 ;
      RECT 17.17 4.135 17.34 4.305 ;
      RECT 16.95 3.475 17.12 3.645 ;
      RECT 16.81 2.095 16.98 2.265 ;
      RECT 16.71 1.415 16.88 1.585 ;
      RECT 16.71 4.135 16.88 4.305 ;
      RECT 16.25 1.415 16.42 1.585 ;
      RECT 16.25 4.135 16.42 4.305 ;
      RECT 16.24 3.015 16.41 3.185 ;
      RECT 15.31 0.915 15.48 1.085 ;
      RECT 15.31 2.395 15.48 2.565 ;
      RECT 15.31 6.315 15.48 6.485 ;
      RECT 15.31 7.795 15.48 7.965 ;
      RECT 14.96 0.105 15.13 0.275 ;
      RECT 14.96 4.165 15.13 4.335 ;
      RECT 14.96 4.545 15.13 4.715 ;
      RECT 14.96 8.605 15.13 8.775 ;
      RECT 14.94 2.765 15.11 2.935 ;
      RECT 14.94 5.945 15.11 6.115 ;
      RECT 14.32 0.915 14.49 1.085 ;
      RECT 14.32 2.395 14.49 2.565 ;
      RECT 14.32 6.315 14.49 6.485 ;
      RECT 14.32 7.795 14.49 7.965 ;
      RECT 13.97 0.105 14.14 0.275 ;
      RECT 13.97 4.165 14.14 4.335 ;
      RECT 13.97 4.545 14.14 4.715 ;
      RECT 13.97 8.605 14.14 8.775 ;
      RECT 13.95 2.765 14.12 2.935 ;
      RECT 13.95 5.945 14.12 6.115 ;
      RECT 13.265 0.105 13.435 0.275 ;
      RECT 13.265 4.165 13.435 4.335 ;
      RECT 13.265 4.545 13.435 4.715 ;
      RECT 13.265 8.605 13.435 8.775 ;
      RECT 12.955 2.025 13.125 2.195 ;
      RECT 12.955 6.685 13.125 6.855 ;
      RECT 12.585 0.105 12.755 0.275 ;
      RECT 12.585 8.605 12.755 8.775 ;
      RECT 12.525 0.915 12.695 1.085 ;
      RECT 12.525 1.655 12.695 1.825 ;
      RECT 12.525 7.055 12.695 7.225 ;
      RECT 12.525 7.795 12.695 7.965 ;
      RECT 12.15 2.395 12.32 2.565 ;
      RECT 12.15 6.315 12.32 6.485 ;
      RECT 11.905 0.105 12.075 0.275 ;
      RECT 11.905 8.605 12.075 8.775 ;
      RECT 11.225 0.105 11.395 0.275 ;
      RECT 11.225 8.605 11.395 8.775 ;
      RECT 11.155 2.765 11.325 2.935 ;
      RECT 11.155 5.945 11.325 6.115 ;
      RECT 9.6 1.415 9.77 1.585 ;
      RECT 9.6 4.135 9.77 4.305 ;
      RECT 9.23 2.875 9.4 3.045 ;
      RECT 9.14 1.415 9.31 1.585 ;
      RECT 9.14 4.135 9.31 4.305 ;
      RECT 8.91 2.045 9.08 2.215 ;
      RECT 8.765 2.485 8.935 2.655 ;
      RECT 8.68 1.415 8.85 1.585 ;
      RECT 8.68 4.135 8.85 4.305 ;
      RECT 8.22 1.415 8.39 1.585 ;
      RECT 8.22 4.135 8.39 4.305 ;
      RECT 8.155 2.525 8.325 2.695 ;
      RECT 7.81 2.16 7.98 2.33 ;
      RECT 7.8 3.52 7.97 3.69 ;
      RECT 7.76 1.415 7.93 1.585 ;
      RECT 7.76 4.135 7.93 4.305 ;
      RECT 7.385 2.76 7.555 2.93 ;
      RECT 7.3 1.415 7.47 1.585 ;
      RECT 7.3 4.135 7.47 4.305 ;
      RECT 7.035 2.235 7.205 2.405 ;
      RECT 6.855 3.55 7.025 3.72 ;
      RECT 6.84 1.415 7.01 1.585 ;
      RECT 6.84 4.135 7.01 4.305 ;
      RECT 6.575 2.865 6.745 3.035 ;
      RECT 6.38 1.415 6.55 1.585 ;
      RECT 6.38 4.135 6.55 4.305 ;
      RECT 6.255 2.49 6.425 2.66 ;
      RECT 5.92 1.415 6.09 1.585 ;
      RECT 5.92 4.135 6.09 4.305 ;
      RECT 5.565 1.97 5.735 2.14 ;
      RECT 5.49 2.44 5.66 2.61 ;
      RECT 5.46 1.415 5.63 1.585 ;
      RECT 5.46 4.135 5.63 4.305 ;
      RECT 5 1.415 5.17 1.585 ;
      RECT 5 4.135 5.17 4.305 ;
      RECT 4.64 2.165 4.81 2.335 ;
      RECT 4.54 1.415 4.71 1.585 ;
      RECT 4.54 4.135 4.71 4.305 ;
      RECT 4.3 3.36 4.47 3.53 ;
      RECT 4.265 2.695 4.435 2.865 ;
      RECT 4.08 1.415 4.25 1.585 ;
      RECT 4.08 4.135 4.25 4.305 ;
      RECT 3.655 2.55 3.825 2.72 ;
      RECT 3.62 1.415 3.79 1.585 ;
      RECT 3.62 4.135 3.79 4.305 ;
      RECT 3.585 3.25 3.755 3.42 ;
      RECT 3.525 2.085 3.695 2.255 ;
      RECT 3.16 1.415 3.33 1.585 ;
      RECT 3.16 4.135 3.33 4.305 ;
      RECT 2.885 3 3.055 3.17 ;
      RECT 2.7 1.415 2.87 1.585 ;
      RECT 2.7 4.135 2.87 4.305 ;
      RECT 2.38 2.505 2.55 2.675 ;
      RECT 2.24 1.415 2.41 1.585 ;
      RECT 2.24 4.135 2.41 4.305 ;
      RECT 2.16 3.25 2.33 3.42 ;
      RECT 1.955 2.13 2.125 2.3 ;
      RECT 1.78 1.415 1.95 1.585 ;
      RECT 1.78 4.135 1.95 4.305 ;
      RECT 1.685 3 1.855 3.17 ;
      RECT 1.645 2.43 1.815 2.6 ;
      RECT 1.32 1.415 1.49 1.585 ;
      RECT 1.32 4.135 1.49 4.305 ;
      RECT 1.1 3.475 1.27 3.645 ;
      RECT 0.96 2.095 1.13 2.265 ;
      RECT 0.86 1.415 1.03 1.585 ;
      RECT 0.86 4.135 1.03 4.305 ;
      RECT 0.4 1.415 0.57 1.585 ;
      RECT 0.4 4.135 0.57 4.305 ;
      RECT 0.39 3.015 0.56 3.185 ;
    LAYER li ;
      RECT 71.785 0 71.955 2.085 ;
      RECT 69.825 0 69.995 2.085 ;
      RECT 67.385 0 67.555 2.085 ;
      RECT 66.425 0 66.595 2.085 ;
      RECT 65.905 0 66.075 2.085 ;
      RECT 64.945 0 65.115 2.085 ;
      RECT 63.985 0 64.155 2.085 ;
      RECT 55.935 0 56.105 2.085 ;
      RECT 53.975 0 54.145 2.085 ;
      RECT 51.535 0 51.705 2.085 ;
      RECT 50.575 0 50.745 2.085 ;
      RECT 50.055 0 50.225 2.085 ;
      RECT 49.095 0 49.265 2.085 ;
      RECT 48.135 0 48.305 2.085 ;
      RECT 40.085 0 40.255 2.085 ;
      RECT 38.125 0 38.295 2.085 ;
      RECT 35.685 0 35.855 2.085 ;
      RECT 34.725 0 34.895 2.085 ;
      RECT 34.205 0 34.375 2.085 ;
      RECT 33.245 0 33.415 2.085 ;
      RECT 32.285 0 32.455 2.085 ;
      RECT 24.235 0 24.405 2.085 ;
      RECT 22.275 0 22.445 2.085 ;
      RECT 19.835 0 20.005 2.085 ;
      RECT 18.875 0 19.045 2.085 ;
      RECT 18.355 0 18.525 2.085 ;
      RECT 17.395 0 17.565 2.085 ;
      RECT 16.435 0 16.605 2.085 ;
      RECT 8.385 0 8.555 2.085 ;
      RECT 6.425 0 6.595 2.085 ;
      RECT 3.985 0 4.155 2.085 ;
      RECT 3.025 0 3.195 2.085 ;
      RECT 2.505 0 2.675 2.085 ;
      RECT 1.545 0 1.715 2.085 ;
      RECT 0.585 0 0.755 2.085 ;
      RECT 63.77 0 73.37 1.59 ;
      RECT 47.92 0 57.52 1.59 ;
      RECT 32.07 0 41.67 1.59 ;
      RECT 16.22 0 25.82 1.59 ;
      RECT 0.37 0 9.97 1.59 ;
      RECT 63.655 1.415 73.485 1.585 ;
      RECT 63.77 0 73.485 1.585 ;
      RECT 47.805 1.415 57.635 1.585 ;
      RECT 47.92 0 57.635 1.585 ;
      RECT 31.955 1.415 41.785 1.585 ;
      RECT 32.07 0 41.785 1.585 ;
      RECT 16.105 1.415 25.935 1.585 ;
      RECT 16.22 0 25.935 1.585 ;
      RECT 0.255 1.415 10.085 1.585 ;
      RECT 0.37 0 10.085 1.585 ;
      RECT 78.28 0 78.45 0.935 ;
      RECT 77.29 0 77.46 0.935 ;
      RECT 74.545 0 74.715 0.935 ;
      RECT 62.43 0 62.6 0.935 ;
      RECT 61.44 0 61.61 0.935 ;
      RECT 58.695 0 58.865 0.935 ;
      RECT 46.58 0 46.75 0.935 ;
      RECT 45.59 0 45.76 0.935 ;
      RECT 42.845 0 43.015 0.935 ;
      RECT 30.73 0 30.9 0.935 ;
      RECT 29.74 0 29.91 0.935 ;
      RECT 26.995 0 27.165 0.935 ;
      RECT 14.88 0 15.05 0.935 ;
      RECT 13.89 0 14.06 0.935 ;
      RECT 11.145 0 11.315 0.935 ;
      RECT 0 0 79.25 0.305 ;
      RECT 78.28 3.405 78.45 5.475 ;
      RECT 77.29 3.405 77.46 5.475 ;
      RECT 74.545 3.405 74.715 5.475 ;
      RECT 62.43 3.405 62.6 5.475 ;
      RECT 61.44 3.405 61.61 5.475 ;
      RECT 58.695 3.405 58.865 5.475 ;
      RECT 46.58 3.405 46.75 5.475 ;
      RECT 45.59 3.405 45.76 5.475 ;
      RECT 42.845 3.405 43.015 5.475 ;
      RECT 30.73 3.405 30.9 5.475 ;
      RECT 29.74 3.405 29.91 5.475 ;
      RECT 26.995 3.405 27.165 5.475 ;
      RECT 14.88 3.405 15.05 5.475 ;
      RECT 13.89 3.405 14.06 5.475 ;
      RECT 11.145 3.405 11.315 5.475 ;
      RECT 63.19 4.135 63.69 4.75 ;
      RECT 0.005 4.305 79.25 4.745 ;
      RECT 0.255 4.135 79.25 4.745 ;
      RECT 72.745 3.635 72.915 4.745 ;
      RECT 71.785 3.635 71.955 4.745 ;
      RECT 69.345 3.635 69.515 4.745 ;
      RECT 68.345 3.635 68.515 4.745 ;
      RECT 67.385 3.635 67.555 4.745 ;
      RECT 64.945 3.635 65.115 4.745 ;
      RECT 56.895 3.635 57.065 4.745 ;
      RECT 55.935 3.635 56.105 4.745 ;
      RECT 53.495 3.635 53.665 4.745 ;
      RECT 52.495 3.635 52.665 4.745 ;
      RECT 51.535 3.635 51.705 4.745 ;
      RECT 49.095 3.635 49.265 4.745 ;
      RECT 47.34 4.13 47.84 4.745 ;
      RECT 41.045 3.635 41.215 4.745 ;
      RECT 40.085 3.635 40.255 4.745 ;
      RECT 37.645 3.635 37.815 4.745 ;
      RECT 36.645 3.635 36.815 4.745 ;
      RECT 35.685 3.635 35.855 4.745 ;
      RECT 33.245 3.635 33.415 4.745 ;
      RECT 25.195 3.635 25.365 4.745 ;
      RECT 24.235 3.635 24.405 4.745 ;
      RECT 21.795 3.635 21.965 4.745 ;
      RECT 20.795 3.635 20.965 4.745 ;
      RECT 19.835 3.635 20.005 4.745 ;
      RECT 17.395 3.635 17.565 4.745 ;
      RECT 9.345 3.635 9.515 4.745 ;
      RECT 8.385 3.635 8.555 4.745 ;
      RECT 5.945 3.635 6.115 4.745 ;
      RECT 4.945 3.635 5.115 4.745 ;
      RECT 3.985 3.635 4.155 4.745 ;
      RECT 1.545 3.635 1.715 4.745 ;
      RECT 0 8.575 79.25 8.88 ;
      RECT 78.28 7.945 78.45 8.88 ;
      RECT 77.29 7.945 77.46 8.88 ;
      RECT 74.545 7.945 74.715 8.88 ;
      RECT 62.43 7.945 62.6 8.88 ;
      RECT 61.44 7.945 61.61 8.88 ;
      RECT 58.695 7.945 58.865 8.88 ;
      RECT 46.58 7.945 46.75 8.88 ;
      RECT 45.59 7.945 45.76 8.88 ;
      RECT 42.845 7.945 43.015 8.88 ;
      RECT 30.73 7.945 30.9 8.88 ;
      RECT 29.74 7.945 29.91 8.88 ;
      RECT 26.995 7.945 27.165 8.88 ;
      RECT 14.88 7.945 15.05 8.88 ;
      RECT 13.89 7.945 14.06 8.88 ;
      RECT 11.145 7.945 11.315 8.88 ;
      RECT 78.71 2.395 78.88 3.865 ;
      RECT 78.715 2.16 78.885 2.525 ;
      RECT 78.34 1.74 78.51 2.935 ;
      RECT 78.34 1.74 78.805 1.91 ;
      RECT 78.34 6.97 78.805 7.14 ;
      RECT 78.34 5.945 78.51 7.14 ;
      RECT 77.35 1.74 77.52 2.935 ;
      RECT 77.35 1.74 77.815 1.91 ;
      RECT 77.35 6.97 77.815 7.14 ;
      RECT 77.35 5.945 77.52 7.14 ;
      RECT 75.495 2.635 75.665 3.865 ;
      RECT 75.55 0.855 75.72 2.805 ;
      RECT 75.495 0.575 75.665 1.025 ;
      RECT 75.495 7.855 75.665 8.305 ;
      RECT 75.55 6.075 75.72 8.025 ;
      RECT 75.495 5.015 75.665 6.245 ;
      RECT 74.975 0.575 75.145 3.865 ;
      RECT 74.975 2.075 75.38 2.405 ;
      RECT 74.975 1.235 75.38 1.565 ;
      RECT 74.975 5.015 75.145 8.305 ;
      RECT 74.975 7.315 75.38 7.645 ;
      RECT 74.975 6.475 75.38 6.805 ;
      RECT 72.31 1.975 73.04 2.215 ;
      RECT 72.852 1.77 73.04 2.215 ;
      RECT 72.68 1.782 73.055 2.209 ;
      RECT 72.595 1.797 73.075 2.194 ;
      RECT 72.595 1.812 73.08 2.184 ;
      RECT 72.55 1.832 73.095 2.176 ;
      RECT 72.527 1.867 73.11 2.13 ;
      RECT 72.441 1.89 73.115 2.09 ;
      RECT 72.441 1.908 73.125 2.06 ;
      RECT 72.31 1.977 73.13 2.023 ;
      RECT 72.355 1.92 73.125 2.06 ;
      RECT 72.441 1.872 73.11 2.13 ;
      RECT 72.527 1.841 73.095 2.176 ;
      RECT 72.55 1.822 73.08 2.184 ;
      RECT 72.595 1.795 73.055 2.209 ;
      RECT 72.68 1.777 73.04 2.215 ;
      RECT 72.766 1.771 73.04 2.215 ;
      RECT 72.852 1.766 72.985 2.215 ;
      RECT 72.938 1.761 72.985 2.215 ;
      RECT 72.63 2.659 72.8 3.045 ;
      RECT 72.625 2.659 72.8 3.04 ;
      RECT 72.6 2.659 72.8 3.005 ;
      RECT 72.6 2.687 72.81 2.995 ;
      RECT 72.58 2.687 72.81 2.955 ;
      RECT 72.575 2.687 72.81 2.928 ;
      RECT 72.575 2.705 72.815 2.92 ;
      RECT 72.52 2.705 72.815 2.855 ;
      RECT 72.52 2.722 72.825 2.838 ;
      RECT 72.51 2.722 72.825 2.778 ;
      RECT 72.51 2.739 72.83 2.775 ;
      RECT 72.505 2.575 72.675 2.753 ;
      RECT 72.505 2.609 72.761 2.753 ;
      RECT 72.5 3.375 72.505 3.388 ;
      RECT 72.495 3.27 72.5 3.393 ;
      RECT 72.47 3.13 72.495 3.408 ;
      RECT 72.435 3.081 72.47 3.44 ;
      RECT 72.43 3.049 72.435 3.46 ;
      RECT 72.425 3.04 72.43 3.46 ;
      RECT 72.345 3.005 72.425 3.46 ;
      RECT 72.282 2.975 72.345 3.46 ;
      RECT 72.196 2.963 72.282 3.46 ;
      RECT 72.11 2.949 72.196 3.46 ;
      RECT 72.03 2.936 72.11 3.446 ;
      RECT 71.995 2.928 72.03 3.426 ;
      RECT 71.985 2.925 71.995 3.417 ;
      RECT 71.955 2.92 71.985 3.404 ;
      RECT 71.905 2.895 71.955 3.38 ;
      RECT 71.891 2.869 71.905 3.362 ;
      RECT 71.805 2.829 71.891 3.338 ;
      RECT 71.76 2.777 71.805 3.307 ;
      RECT 71.75 2.752 71.76 3.294 ;
      RECT 71.745 2.533 71.75 2.555 ;
      RECT 71.74 2.735 71.75 3.29 ;
      RECT 71.74 2.531 71.745 2.645 ;
      RECT 71.73 2.527 71.74 3.286 ;
      RECT 71.686 2.525 71.73 3.274 ;
      RECT 71.6 2.525 71.686 3.245 ;
      RECT 71.57 2.525 71.6 3.218 ;
      RECT 71.555 2.525 71.57 3.206 ;
      RECT 71.515 2.537 71.555 3.191 ;
      RECT 71.495 2.556 71.515 3.17 ;
      RECT 71.485 2.566 71.495 3.154 ;
      RECT 71.475 2.572 71.485 3.143 ;
      RECT 71.455 2.582 71.475 3.126 ;
      RECT 71.45 2.591 71.455 3.113 ;
      RECT 71.445 2.595 71.45 3.063 ;
      RECT 71.435 2.601 71.445 2.98 ;
      RECT 71.43 2.605 71.435 2.894 ;
      RECT 71.425 2.625 71.43 2.831 ;
      RECT 71.42 2.648 71.425 2.778 ;
      RECT 71.415 2.666 71.42 2.723 ;
      RECT 72.025 2.485 72.195 2.745 ;
      RECT 72.195 2.45 72.24 2.731 ;
      RECT 72.156 2.452 72.245 2.714 ;
      RECT 72.045 2.469 72.331 2.685 ;
      RECT 72.045 2.484 72.335 2.657 ;
      RECT 72.045 2.465 72.245 2.714 ;
      RECT 72.07 2.453 72.195 2.745 ;
      RECT 72.156 2.451 72.24 2.731 ;
      RECT 71.21 1.84 71.38 2.33 ;
      RECT 71.21 1.84 71.415 2.31 ;
      RECT 71.345 1.76 71.455 2.27 ;
      RECT 71.326 1.764 71.475 2.24 ;
      RECT 71.24 1.772 71.495 2.223 ;
      RECT 71.24 1.778 71.5 2.213 ;
      RECT 71.24 1.787 71.52 2.201 ;
      RECT 71.215 1.812 71.55 2.179 ;
      RECT 71.215 1.832 71.555 2.159 ;
      RECT 71.21 1.845 71.565 2.139 ;
      RECT 71.21 1.912 71.57 2.12 ;
      RECT 71.21 2.045 71.575 2.107 ;
      RECT 71.205 1.85 71.565 1.94 ;
      RECT 71.215 1.807 71.52 2.201 ;
      RECT 71.326 1.762 71.455 2.27 ;
      RECT 71.2 3.515 71.5 3.77 ;
      RECT 71.285 3.481 71.5 3.77 ;
      RECT 71.285 3.484 71.505 3.63 ;
      RECT 71.22 3.505 71.505 3.63 ;
      RECT 71.255 3.495 71.5 3.77 ;
      RECT 71.25 3.5 71.505 3.63 ;
      RECT 71.285 3.479 71.486 3.77 ;
      RECT 71.371 3.47 71.486 3.77 ;
      RECT 71.371 3.464 71.4 3.77 ;
      RECT 70.86 3.105 70.87 3.595 ;
      RECT 70.52 3.04 70.53 3.34 ;
      RECT 71.035 3.212 71.04 3.431 ;
      RECT 71.025 3.192 71.035 3.448 ;
      RECT 71.015 3.172 71.025 3.478 ;
      RECT 71.01 3.162 71.015 3.493 ;
      RECT 71.005 3.158 71.01 3.498 ;
      RECT 70.99 3.15 71.005 3.505 ;
      RECT 70.95 3.13 70.99 3.53 ;
      RECT 70.925 3.112 70.95 3.563 ;
      RECT 70.92 3.11 70.925 3.576 ;
      RECT 70.9 3.107 70.92 3.58 ;
      RECT 70.87 3.105 70.9 3.59 ;
      RECT 70.8 3.107 70.86 3.591 ;
      RECT 70.78 3.107 70.8 3.585 ;
      RECT 70.755 3.105 70.78 3.582 ;
      RECT 70.72 3.1 70.755 3.578 ;
      RECT 70.7 3.094 70.72 3.565 ;
      RECT 70.69 3.091 70.7 3.553 ;
      RECT 70.67 3.088 70.69 3.538 ;
      RECT 70.65 3.084 70.67 3.52 ;
      RECT 70.645 3.081 70.65 3.51 ;
      RECT 70.64 3.08 70.645 3.508 ;
      RECT 70.63 3.077 70.64 3.5 ;
      RECT 70.62 3.071 70.63 3.483 ;
      RECT 70.61 3.065 70.62 3.465 ;
      RECT 70.6 3.059 70.61 3.453 ;
      RECT 70.59 3.053 70.6 3.433 ;
      RECT 70.585 3.049 70.59 3.418 ;
      RECT 70.58 3.047 70.585 3.41 ;
      RECT 70.575 3.045 70.58 3.403 ;
      RECT 70.57 3.043 70.575 3.393 ;
      RECT 70.565 3.041 70.57 3.387 ;
      RECT 70.555 3.04 70.565 3.377 ;
      RECT 70.545 3.04 70.555 3.368 ;
      RECT 70.53 3.04 70.545 3.353 ;
      RECT 70.49 3.04 70.52 3.337 ;
      RECT 70.47 3.042 70.49 3.332 ;
      RECT 70.465 3.047 70.47 3.33 ;
      RECT 70.435 3.055 70.465 3.328 ;
      RECT 70.405 3.07 70.435 3.327 ;
      RECT 70.36 3.092 70.405 3.332 ;
      RECT 70.355 3.107 70.36 3.336 ;
      RECT 70.34 3.112 70.355 3.338 ;
      RECT 70.335 3.116 70.34 3.34 ;
      RECT 70.275 3.139 70.335 3.349 ;
      RECT 70.255 3.165 70.275 3.362 ;
      RECT 70.245 3.172 70.255 3.366 ;
      RECT 70.23 3.179 70.245 3.369 ;
      RECT 70.21 3.189 70.23 3.372 ;
      RECT 70.205 3.197 70.21 3.375 ;
      RECT 70.16 3.202 70.205 3.382 ;
      RECT 70.15 3.205 70.16 3.389 ;
      RECT 70.14 3.205 70.15 3.393 ;
      RECT 70.105 3.207 70.14 3.405 ;
      RECT 70.085 3.21 70.105 3.418 ;
      RECT 70.045 3.213 70.085 3.429 ;
      RECT 70.03 3.215 70.045 3.442 ;
      RECT 70.02 3.215 70.03 3.447 ;
      RECT 69.995 3.216 70.02 3.455 ;
      RECT 69.985 3.218 69.995 3.46 ;
      RECT 69.98 3.219 69.985 3.463 ;
      RECT 69.955 3.217 69.98 3.466 ;
      RECT 69.94 3.215 69.955 3.467 ;
      RECT 69.92 3.212 69.94 3.469 ;
      RECT 69.9 3.207 69.92 3.469 ;
      RECT 69.84 3.202 69.9 3.466 ;
      RECT 69.805 3.177 69.84 3.462 ;
      RECT 69.795 3.154 69.805 3.46 ;
      RECT 69.765 3.131 69.795 3.46 ;
      RECT 69.755 3.11 69.765 3.46 ;
      RECT 69.73 3.092 69.755 3.458 ;
      RECT 69.715 3.07 69.73 3.455 ;
      RECT 69.7 3.052 69.715 3.453 ;
      RECT 69.68 3.042 69.7 3.451 ;
      RECT 69.665 3.037 69.68 3.45 ;
      RECT 69.65 3.035 69.665 3.449 ;
      RECT 69.62 3.036 69.65 3.447 ;
      RECT 69.6 3.039 69.62 3.445 ;
      RECT 69.543 3.043 69.6 3.445 ;
      RECT 69.457 3.052 69.543 3.445 ;
      RECT 69.371 3.063 69.457 3.445 ;
      RECT 69.285 3.074 69.371 3.445 ;
      RECT 69.265 3.081 69.285 3.453 ;
      RECT 69.255 3.084 69.265 3.46 ;
      RECT 69.19 3.089 69.255 3.478 ;
      RECT 69.16 3.096 69.19 3.503 ;
      RECT 69.15 3.099 69.16 3.51 ;
      RECT 69.105 3.103 69.15 3.515 ;
      RECT 69.075 3.108 69.105 3.52 ;
      RECT 69.074 3.11 69.075 3.52 ;
      RECT 68.988 3.116 69.074 3.52 ;
      RECT 68.902 3.127 68.988 3.52 ;
      RECT 68.816 3.139 68.902 3.52 ;
      RECT 68.73 3.15 68.816 3.52 ;
      RECT 68.715 3.157 68.73 3.515 ;
      RECT 68.71 3.159 68.715 3.509 ;
      RECT 68.69 3.17 68.71 3.504 ;
      RECT 68.68 3.188 68.69 3.498 ;
      RECT 68.675 3.2 68.68 3.298 ;
      RECT 70.97 1.953 70.99 2.04 ;
      RECT 70.965 1.888 70.97 2.072 ;
      RECT 70.955 1.855 70.965 2.077 ;
      RECT 70.95 1.835 70.955 2.083 ;
      RECT 70.92 1.835 70.95 2.1 ;
      RECT 70.871 1.835 70.92 2.136 ;
      RECT 70.785 1.835 70.871 2.194 ;
      RECT 70.756 1.845 70.785 2.243 ;
      RECT 70.67 1.887 70.756 2.296 ;
      RECT 70.65 1.925 70.67 2.343 ;
      RECT 70.625 1.942 70.65 2.363 ;
      RECT 70.615 1.956 70.625 2.383 ;
      RECT 70.61 1.962 70.615 2.393 ;
      RECT 70.605 1.966 70.61 2.4 ;
      RECT 70.555 1.986 70.605 2.405 ;
      RECT 70.49 2.03 70.555 2.405 ;
      RECT 70.465 2.08 70.49 2.405 ;
      RECT 70.455 2.11 70.465 2.405 ;
      RECT 70.45 2.137 70.455 2.405 ;
      RECT 70.445 2.155 70.45 2.405 ;
      RECT 70.435 2.197 70.445 2.405 ;
      RECT 70.785 2.755 70.955 2.93 ;
      RECT 70.725 2.583 70.785 2.918 ;
      RECT 70.715 2.576 70.725 2.901 ;
      RECT 70.67 2.755 70.955 2.881 ;
      RECT 70.651 2.755 70.955 2.859 ;
      RECT 70.565 2.755 70.955 2.824 ;
      RECT 70.545 2.575 70.715 2.78 ;
      RECT 70.545 2.722 70.95 2.78 ;
      RECT 70.545 2.67 70.925 2.78 ;
      RECT 70.545 2.625 70.89 2.78 ;
      RECT 70.545 2.607 70.855 2.78 ;
      RECT 70.545 2.597 70.85 2.78 ;
      RECT 70.265 3.555 70.455 3.78 ;
      RECT 70.255 3.556 70.46 3.775 ;
      RECT 70.255 3.558 70.47 3.755 ;
      RECT 70.255 3.562 70.475 3.74 ;
      RECT 70.255 3.549 70.425 3.775 ;
      RECT 70.255 3.552 70.45 3.775 ;
      RECT 70.265 3.548 70.425 3.78 ;
      RECT 70.351 3.546 70.425 3.78 ;
      RECT 69.975 2.797 70.145 3.035 ;
      RECT 69.975 2.797 70.231 2.949 ;
      RECT 69.975 2.797 70.235 2.859 ;
      RECT 70.025 2.57 70.245 2.838 ;
      RECT 70.02 2.587 70.25 2.811 ;
      RECT 69.985 2.745 70.25 2.811 ;
      RECT 70.005 2.595 70.145 3.035 ;
      RECT 69.995 2.677 70.255 2.794 ;
      RECT 69.99 2.725 70.255 2.794 ;
      RECT 69.995 2.635 70.25 2.811 ;
      RECT 70.02 2.572 70.245 2.838 ;
      RECT 69.585 2.547 69.755 2.745 ;
      RECT 69.585 2.547 69.8 2.72 ;
      RECT 69.655 2.49 69.825 2.678 ;
      RECT 69.63 2.505 69.825 2.678 ;
      RECT 69.245 2.551 69.275 2.745 ;
      RECT 69.24 2.523 69.245 2.745 ;
      RECT 69.21 2.497 69.24 2.747 ;
      RECT 69.185 2.455 69.21 2.75 ;
      RECT 69.175 2.427 69.185 2.752 ;
      RECT 69.14 2.407 69.175 2.754 ;
      RECT 69.075 2.392 69.14 2.76 ;
      RECT 69.025 2.39 69.075 2.766 ;
      RECT 69.002 2.392 69.025 2.771 ;
      RECT 68.916 2.403 69.002 2.777 ;
      RECT 68.83 2.421 68.916 2.787 ;
      RECT 68.815 2.432 68.83 2.793 ;
      RECT 68.745 2.455 68.815 2.799 ;
      RECT 68.69 2.487 68.745 2.807 ;
      RECT 68.65 2.51 68.69 2.813 ;
      RECT 68.636 2.523 68.65 2.816 ;
      RECT 68.55 2.545 68.636 2.822 ;
      RECT 68.535 2.57 68.55 2.828 ;
      RECT 68.495 2.585 68.535 2.832 ;
      RECT 68.445 2.6 68.495 2.837 ;
      RECT 68.42 2.607 68.445 2.841 ;
      RECT 68.36 2.602 68.42 2.845 ;
      RECT 68.345 2.593 68.36 2.849 ;
      RECT 68.275 2.583 68.345 2.845 ;
      RECT 68.25 2.575 68.27 2.835 ;
      RECT 68.191 2.575 68.25 2.813 ;
      RECT 68.105 2.575 68.191 2.77 ;
      RECT 68.27 2.575 68.275 2.84 ;
      RECT 68.965 1.806 69.135 2.14 ;
      RECT 68.935 1.806 69.135 2.135 ;
      RECT 68.875 1.773 68.935 2.123 ;
      RECT 68.875 1.829 69.145 2.118 ;
      RECT 68.85 1.829 69.145 2.112 ;
      RECT 68.845 1.77 68.875 2.109 ;
      RECT 68.83 1.776 68.965 2.107 ;
      RECT 68.825 1.784 69.05 2.095 ;
      RECT 68.825 1.836 69.16 2.048 ;
      RECT 68.81 1.792 69.05 2.043 ;
      RECT 68.81 1.862 69.17 1.984 ;
      RECT 68.78 1.812 69.135 1.945 ;
      RECT 68.78 1.902 69.18 1.941 ;
      RECT 68.83 1.781 69.05 2.107 ;
      RECT 68.17 2.111 68.225 2.375 ;
      RECT 68.17 2.111 68.29 2.374 ;
      RECT 68.17 2.111 68.315 2.373 ;
      RECT 68.17 2.111 68.38 2.372 ;
      RECT 68.315 2.077 68.395 2.371 ;
      RECT 68.13 2.121 68.54 2.37 ;
      RECT 68.17 2.118 68.54 2.37 ;
      RECT 68.13 2.126 68.545 2.363 ;
      RECT 68.115 2.128 68.545 2.362 ;
      RECT 68.115 2.135 68.55 2.358 ;
      RECT 68.095 2.134 68.545 2.354 ;
      RECT 68.095 2.142 68.555 2.353 ;
      RECT 68.09 2.139 68.55 2.349 ;
      RECT 68.09 2.152 68.565 2.348 ;
      RECT 68.075 2.142 68.555 2.347 ;
      RECT 68.04 2.155 68.565 2.34 ;
      RECT 68.225 2.11 68.535 2.37 ;
      RECT 68.225 2.095 68.485 2.37 ;
      RECT 68.29 2.082 68.42 2.37 ;
      RECT 67.835 3.171 67.85 3.564 ;
      RECT 67.8 3.176 67.85 3.563 ;
      RECT 67.835 3.175 67.895 3.562 ;
      RECT 67.78 3.186 67.895 3.561 ;
      RECT 67.795 3.182 67.895 3.561 ;
      RECT 67.76 3.192 67.97 3.558 ;
      RECT 67.76 3.211 68.015 3.556 ;
      RECT 67.76 3.218 68.02 3.553 ;
      RECT 67.745 3.195 67.97 3.55 ;
      RECT 67.725 3.2 67.97 3.543 ;
      RECT 67.72 3.204 67.97 3.539 ;
      RECT 67.72 3.221 68.03 3.538 ;
      RECT 67.7 3.215 68.015 3.534 ;
      RECT 67.7 3.224 68.035 3.528 ;
      RECT 67.695 3.23 68.035 3.3 ;
      RECT 67.76 3.19 67.895 3.558 ;
      RECT 67.635 2.553 67.835 2.865 ;
      RECT 67.71 2.531 67.835 2.865 ;
      RECT 67.65 2.55 67.84 2.85 ;
      RECT 67.62 2.561 67.84 2.848 ;
      RECT 67.635 2.556 67.845 2.814 ;
      RECT 67.62 2.66 67.85 2.781 ;
      RECT 67.65 2.532 67.835 2.865 ;
      RECT 67.71 2.51 67.81 2.865 ;
      RECT 67.735 2.507 67.81 2.865 ;
      RECT 67.735 2.502 67.755 2.865 ;
      RECT 67.14 2.57 67.315 2.745 ;
      RECT 67.135 2.57 67.315 2.743 ;
      RECT 67.11 2.57 67.315 2.738 ;
      RECT 67.055 2.55 67.225 2.728 ;
      RECT 67.055 2.557 67.29 2.728 ;
      RECT 67.14 3.237 67.155 3.42 ;
      RECT 67.13 3.215 67.14 3.42 ;
      RECT 67.115 3.195 67.13 3.42 ;
      RECT 67.105 3.17 67.115 3.42 ;
      RECT 67.075 3.135 67.105 3.42 ;
      RECT 67.04 3.075 67.075 3.42 ;
      RECT 67.035 3.037 67.04 3.42 ;
      RECT 66.985 2.988 67.035 3.42 ;
      RECT 66.975 2.938 66.985 3.408 ;
      RECT 66.96 2.917 66.975 3.368 ;
      RECT 66.94 2.885 66.96 3.318 ;
      RECT 66.915 2.841 66.94 3.258 ;
      RECT 66.91 2.813 66.915 3.213 ;
      RECT 66.905 2.804 66.91 3.199 ;
      RECT 66.9 2.797 66.905 3.186 ;
      RECT 66.895 2.792 66.9 3.175 ;
      RECT 66.89 2.777 66.895 3.165 ;
      RECT 66.885 2.755 66.89 3.152 ;
      RECT 66.875 2.715 66.885 3.127 ;
      RECT 66.85 2.645 66.875 3.083 ;
      RECT 66.845 2.585 66.85 3.048 ;
      RECT 66.83 2.565 66.845 3.015 ;
      RECT 66.825 2.565 66.83 2.99 ;
      RECT 66.795 2.565 66.825 2.945 ;
      RECT 66.75 2.565 66.795 2.885 ;
      RECT 66.675 2.565 66.75 2.833 ;
      RECT 66.67 2.565 66.675 2.798 ;
      RECT 66.665 2.565 66.67 2.788 ;
      RECT 66.66 2.565 66.665 2.768 ;
      RECT 66.925 1.785 67.095 2.255 ;
      RECT 66.87 1.778 67.065 2.239 ;
      RECT 66.87 1.792 67.1 2.238 ;
      RECT 66.855 1.793 67.1 2.219 ;
      RECT 66.85 1.811 67.1 2.205 ;
      RECT 66.855 1.794 67.105 2.203 ;
      RECT 66.84 1.825 67.105 2.188 ;
      RECT 66.855 1.8 67.11 2.173 ;
      RECT 66.835 1.84 67.11 2.17 ;
      RECT 66.85 1.812 67.115 2.155 ;
      RECT 66.85 1.824 67.12 2.135 ;
      RECT 66.835 1.84 67.125 2.118 ;
      RECT 66.835 1.85 67.13 1.973 ;
      RECT 66.83 1.85 67.13 1.93 ;
      RECT 66.83 1.865 67.135 1.908 ;
      RECT 66.925 1.775 67.065 2.255 ;
      RECT 66.925 1.773 67.035 2.255 ;
      RECT 67.011 1.77 67.035 2.255 ;
      RECT 66.67 3.437 66.675 3.483 ;
      RECT 66.66 3.285 66.67 3.507 ;
      RECT 66.655 3.13 66.66 3.532 ;
      RECT 66.64 3.092 66.655 3.543 ;
      RECT 66.635 3.075 66.64 3.55 ;
      RECT 66.625 3.063 66.635 3.557 ;
      RECT 66.62 3.054 66.625 3.559 ;
      RECT 66.615 3.052 66.62 3.563 ;
      RECT 66.57 3.043 66.615 3.578 ;
      RECT 66.565 3.035 66.57 3.592 ;
      RECT 66.56 3.032 66.565 3.596 ;
      RECT 66.545 3.027 66.56 3.604 ;
      RECT 66.49 3.017 66.545 3.615 ;
      RECT 66.455 3.005 66.49 3.616 ;
      RECT 66.446 3 66.455 3.61 ;
      RECT 66.36 3 66.446 3.6 ;
      RECT 66.33 3 66.36 3.578 ;
      RECT 66.32 3 66.325 3.558 ;
      RECT 66.315 3 66.32 3.52 ;
      RECT 66.31 3 66.315 3.478 ;
      RECT 66.305 3 66.31 3.438 ;
      RECT 66.3 3 66.305 3.368 ;
      RECT 66.29 3 66.3 3.29 ;
      RECT 66.285 3 66.29 3.19 ;
      RECT 66.325 3 66.33 3.56 ;
      RECT 65.82 3.082 65.91 3.56 ;
      RECT 65.805 3.085 65.925 3.558 ;
      RECT 65.82 3.084 65.925 3.558 ;
      RECT 65.785 3.091 65.95 3.548 ;
      RECT 65.805 3.085 65.95 3.548 ;
      RECT 65.77 3.097 65.95 3.536 ;
      RECT 65.805 3.088 66 3.529 ;
      RECT 65.756 3.105 66 3.527 ;
      RECT 65.785 3.095 66.01 3.515 ;
      RECT 65.756 3.116 66.04 3.506 ;
      RECT 65.67 3.14 66.04 3.5 ;
      RECT 65.67 3.153 66.08 3.483 ;
      RECT 65.665 3.175 66.08 3.476 ;
      RECT 65.635 3.19 66.08 3.466 ;
      RECT 65.63 3.201 66.08 3.456 ;
      RECT 65.6 3.214 66.08 3.447 ;
      RECT 65.585 3.232 66.08 3.436 ;
      RECT 65.56 3.245 66.08 3.426 ;
      RECT 65.82 3.081 65.83 3.56 ;
      RECT 65.866 2.505 65.905 2.75 ;
      RECT 65.78 2.505 65.915 2.748 ;
      RECT 65.665 2.53 65.915 2.745 ;
      RECT 65.665 2.53 65.92 2.743 ;
      RECT 65.665 2.53 65.935 2.738 ;
      RECT 65.771 2.505 65.95 2.718 ;
      RECT 65.685 2.513 65.95 2.718 ;
      RECT 65.355 1.865 65.525 2.3 ;
      RECT 65.345 1.899 65.525 2.283 ;
      RECT 65.425 1.835 65.595 2.27 ;
      RECT 65.33 1.91 65.595 2.248 ;
      RECT 65.425 1.845 65.6 2.238 ;
      RECT 65.355 1.897 65.63 2.223 ;
      RECT 65.315 1.923 65.63 2.208 ;
      RECT 65.315 1.965 65.64 2.188 ;
      RECT 65.31 1.99 65.645 2.17 ;
      RECT 65.31 2 65.65 2.155 ;
      RECT 65.305 1.937 65.63 2.153 ;
      RECT 65.305 2.01 65.655 2.138 ;
      RECT 65.3 1.947 65.63 2.135 ;
      RECT 65.295 2.031 65.66 2.118 ;
      RECT 65.295 2.063 65.665 2.098 ;
      RECT 65.29 1.977 65.64 2.09 ;
      RECT 65.295 1.962 65.63 2.118 ;
      RECT 65.31 1.932 65.63 2.17 ;
      RECT 65.155 2.519 65.38 2.775 ;
      RECT 65.155 2.552 65.4 2.765 ;
      RECT 65.12 2.552 65.4 2.763 ;
      RECT 65.12 2.565 65.405 2.753 ;
      RECT 65.12 2.585 65.415 2.745 ;
      RECT 65.12 2.682 65.42 2.738 ;
      RECT 65.1 2.43 65.23 2.728 ;
      RECT 65.055 2.585 65.415 2.67 ;
      RECT 65.045 2.43 65.23 2.615 ;
      RECT 65.045 2.462 65.316 2.615 ;
      RECT 65.01 2.992 65.03 3.17 ;
      RECT 64.975 2.945 65.01 3.17 ;
      RECT 64.96 2.885 64.975 3.17 ;
      RECT 64.935 2.832 64.96 3.17 ;
      RECT 64.92 2.785 64.935 3.17 ;
      RECT 64.9 2.762 64.92 3.17 ;
      RECT 64.875 2.727 64.9 3.17 ;
      RECT 64.865 2.573 64.875 3.17 ;
      RECT 64.835 2.568 64.865 3.161 ;
      RECT 64.83 2.565 64.835 3.151 ;
      RECT 64.815 2.565 64.83 3.125 ;
      RECT 64.81 2.565 64.815 3.088 ;
      RECT 64.785 2.565 64.81 3.04 ;
      RECT 64.765 2.565 64.785 2.965 ;
      RECT 64.755 2.565 64.765 2.925 ;
      RECT 64.75 2.565 64.755 2.9 ;
      RECT 64.745 2.565 64.75 2.883 ;
      RECT 64.74 2.565 64.745 2.865 ;
      RECT 64.735 2.566 64.74 2.855 ;
      RECT 64.725 2.568 64.735 2.823 ;
      RECT 64.715 2.57 64.725 2.79 ;
      RECT 64.705 2.573 64.715 2.763 ;
      RECT 65.03 3 65.255 3.17 ;
      RECT 64.36 1.812 64.53 2.265 ;
      RECT 64.36 1.812 64.62 2.231 ;
      RECT 64.36 1.812 64.65 2.215 ;
      RECT 64.36 1.812 64.68 2.188 ;
      RECT 64.616 1.79 64.695 2.17 ;
      RECT 64.395 1.797 64.7 2.155 ;
      RECT 64.395 1.805 64.71 2.118 ;
      RECT 64.355 1.832 64.71 2.09 ;
      RECT 64.34 1.845 64.71 2.055 ;
      RECT 64.36 1.82 64.73 2.045 ;
      RECT 64.335 1.885 64.73 2.015 ;
      RECT 64.335 1.915 64.735 1.998 ;
      RECT 64.33 1.945 64.735 1.985 ;
      RECT 64.395 1.794 64.695 2.17 ;
      RECT 64.53 1.791 64.616 2.249 ;
      RECT 64.481 1.792 64.695 2.17 ;
      RECT 64.625 3.452 64.67 3.645 ;
      RECT 64.615 3.422 64.625 3.645 ;
      RECT 64.61 3.407 64.615 3.645 ;
      RECT 64.57 3.317 64.61 3.645 ;
      RECT 64.565 3.23 64.57 3.645 ;
      RECT 64.555 3.2 64.565 3.645 ;
      RECT 64.55 3.16 64.555 3.645 ;
      RECT 64.54 3.122 64.55 3.645 ;
      RECT 64.535 3.087 64.54 3.645 ;
      RECT 64.515 3.04 64.535 3.645 ;
      RECT 64.5 2.965 64.515 3.645 ;
      RECT 64.495 2.92 64.5 3.64 ;
      RECT 64.49 2.9 64.495 3.613 ;
      RECT 64.485 2.88 64.49 3.598 ;
      RECT 64.48 2.855 64.485 3.578 ;
      RECT 64.475 2.833 64.48 3.563 ;
      RECT 64.47 2.811 64.475 3.545 ;
      RECT 64.465 2.79 64.47 3.535 ;
      RECT 64.455 2.762 64.465 3.505 ;
      RECT 64.445 2.725 64.455 3.473 ;
      RECT 64.435 2.685 64.445 3.44 ;
      RECT 64.425 2.663 64.435 3.41 ;
      RECT 64.395 2.615 64.425 3.342 ;
      RECT 64.38 2.575 64.395 3.269 ;
      RECT 64.37 2.575 64.38 3.235 ;
      RECT 64.365 2.575 64.37 3.21 ;
      RECT 64.36 2.575 64.365 3.195 ;
      RECT 64.355 2.575 64.36 3.173 ;
      RECT 64.35 2.575 64.355 3.16 ;
      RECT 64.335 2.575 64.35 3.125 ;
      RECT 64.315 2.575 64.335 3.065 ;
      RECT 64.305 2.575 64.315 3.015 ;
      RECT 64.285 2.575 64.305 2.963 ;
      RECT 64.265 2.575 64.285 2.92 ;
      RECT 64.255 2.575 64.265 2.908 ;
      RECT 64.225 2.575 64.255 2.895 ;
      RECT 64.195 2.596 64.225 2.875 ;
      RECT 64.185 2.624 64.195 2.855 ;
      RECT 64.17 2.641 64.185 2.823 ;
      RECT 64.165 2.655 64.17 2.79 ;
      RECT 64.16 2.663 64.165 2.763 ;
      RECT 64.155 2.671 64.16 2.725 ;
      RECT 64.16 3.195 64.165 3.53 ;
      RECT 64.125 3.182 64.16 3.529 ;
      RECT 64.055 3.122 64.125 3.528 ;
      RECT 63.975 3.065 64.055 3.527 ;
      RECT 63.84 3.025 63.975 3.526 ;
      RECT 63.84 3.212 64.175 3.515 ;
      RECT 63.8 3.212 64.175 3.505 ;
      RECT 63.8 3.23 64.18 3.5 ;
      RECT 63.8 3.32 64.185 3.49 ;
      RECT 63.795 3.015 63.96 3.47 ;
      RECT 63.79 3.015 63.96 3.213 ;
      RECT 63.79 3.172 64.155 3.213 ;
      RECT 63.79 3.16 64.15 3.213 ;
      RECT 62.49 1.74 62.66 2.935 ;
      RECT 62.49 1.74 62.955 1.91 ;
      RECT 62.49 6.97 62.955 7.14 ;
      RECT 62.49 5.945 62.66 7.14 ;
      RECT 61.5 1.74 61.67 2.935 ;
      RECT 61.5 1.74 61.965 1.91 ;
      RECT 61.5 6.97 61.965 7.14 ;
      RECT 61.5 5.945 61.67 7.14 ;
      RECT 59.645 2.635 59.815 3.865 ;
      RECT 59.7 0.855 59.87 2.805 ;
      RECT 59.645 0.575 59.815 1.025 ;
      RECT 59.645 7.855 59.815 8.305 ;
      RECT 59.7 6.075 59.87 8.025 ;
      RECT 59.645 5.015 59.815 6.245 ;
      RECT 59.125 0.575 59.295 3.865 ;
      RECT 59.125 2.075 59.53 2.405 ;
      RECT 59.125 1.235 59.53 1.565 ;
      RECT 59.125 5.015 59.295 8.305 ;
      RECT 59.125 7.315 59.53 7.645 ;
      RECT 59.125 6.475 59.53 6.805 ;
      RECT 56.46 1.975 57.19 2.215 ;
      RECT 57.002 1.77 57.19 2.215 ;
      RECT 56.83 1.782 57.205 2.209 ;
      RECT 56.745 1.797 57.225 2.194 ;
      RECT 56.745 1.812 57.23 2.184 ;
      RECT 56.7 1.832 57.245 2.176 ;
      RECT 56.677 1.867 57.26 2.13 ;
      RECT 56.591 1.89 57.265 2.09 ;
      RECT 56.591 1.908 57.275 2.06 ;
      RECT 56.46 1.977 57.28 2.023 ;
      RECT 56.505 1.92 57.275 2.06 ;
      RECT 56.591 1.872 57.26 2.13 ;
      RECT 56.677 1.841 57.245 2.176 ;
      RECT 56.7 1.822 57.23 2.184 ;
      RECT 56.745 1.795 57.205 2.209 ;
      RECT 56.83 1.777 57.19 2.215 ;
      RECT 56.916 1.771 57.19 2.215 ;
      RECT 57.002 1.766 57.135 2.215 ;
      RECT 57.088 1.761 57.135 2.215 ;
      RECT 56.78 2.659 56.95 3.045 ;
      RECT 56.775 2.659 56.95 3.04 ;
      RECT 56.75 2.659 56.95 3.005 ;
      RECT 56.75 2.687 56.96 2.995 ;
      RECT 56.73 2.687 56.96 2.955 ;
      RECT 56.725 2.687 56.96 2.928 ;
      RECT 56.725 2.705 56.965 2.92 ;
      RECT 56.67 2.705 56.965 2.855 ;
      RECT 56.67 2.722 56.975 2.838 ;
      RECT 56.66 2.722 56.975 2.778 ;
      RECT 56.66 2.739 56.98 2.775 ;
      RECT 56.655 2.575 56.825 2.753 ;
      RECT 56.655 2.609 56.911 2.753 ;
      RECT 56.65 3.375 56.655 3.388 ;
      RECT 56.645 3.27 56.65 3.393 ;
      RECT 56.62 3.13 56.645 3.408 ;
      RECT 56.585 3.081 56.62 3.44 ;
      RECT 56.58 3.049 56.585 3.46 ;
      RECT 56.575 3.04 56.58 3.46 ;
      RECT 56.495 3.005 56.575 3.46 ;
      RECT 56.432 2.975 56.495 3.46 ;
      RECT 56.346 2.963 56.432 3.46 ;
      RECT 56.26 2.949 56.346 3.46 ;
      RECT 56.18 2.936 56.26 3.446 ;
      RECT 56.145 2.928 56.18 3.426 ;
      RECT 56.135 2.925 56.145 3.417 ;
      RECT 56.105 2.92 56.135 3.404 ;
      RECT 56.055 2.895 56.105 3.38 ;
      RECT 56.041 2.869 56.055 3.362 ;
      RECT 55.955 2.829 56.041 3.338 ;
      RECT 55.91 2.777 55.955 3.307 ;
      RECT 55.9 2.752 55.91 3.294 ;
      RECT 55.895 2.533 55.9 2.555 ;
      RECT 55.89 2.735 55.9 3.29 ;
      RECT 55.89 2.531 55.895 2.645 ;
      RECT 55.88 2.527 55.89 3.286 ;
      RECT 55.836 2.525 55.88 3.274 ;
      RECT 55.75 2.525 55.836 3.245 ;
      RECT 55.72 2.525 55.75 3.218 ;
      RECT 55.705 2.525 55.72 3.206 ;
      RECT 55.665 2.537 55.705 3.191 ;
      RECT 55.645 2.556 55.665 3.17 ;
      RECT 55.635 2.566 55.645 3.154 ;
      RECT 55.625 2.572 55.635 3.143 ;
      RECT 55.605 2.582 55.625 3.126 ;
      RECT 55.6 2.591 55.605 3.113 ;
      RECT 55.595 2.595 55.6 3.063 ;
      RECT 55.585 2.601 55.595 2.98 ;
      RECT 55.58 2.605 55.585 2.894 ;
      RECT 55.575 2.625 55.58 2.831 ;
      RECT 55.57 2.648 55.575 2.778 ;
      RECT 55.565 2.666 55.57 2.723 ;
      RECT 56.175 2.485 56.345 2.745 ;
      RECT 56.345 2.45 56.39 2.731 ;
      RECT 56.306 2.452 56.395 2.714 ;
      RECT 56.195 2.469 56.481 2.685 ;
      RECT 56.195 2.484 56.485 2.657 ;
      RECT 56.195 2.465 56.395 2.714 ;
      RECT 56.22 2.453 56.345 2.745 ;
      RECT 56.306 2.451 56.39 2.731 ;
      RECT 55.36 1.84 55.53 2.33 ;
      RECT 55.36 1.84 55.565 2.31 ;
      RECT 55.495 1.76 55.605 2.27 ;
      RECT 55.476 1.764 55.625 2.24 ;
      RECT 55.39 1.772 55.645 2.223 ;
      RECT 55.39 1.778 55.65 2.213 ;
      RECT 55.39 1.787 55.67 2.201 ;
      RECT 55.365 1.812 55.7 2.179 ;
      RECT 55.365 1.832 55.705 2.159 ;
      RECT 55.36 1.845 55.715 2.139 ;
      RECT 55.36 1.912 55.72 2.12 ;
      RECT 55.36 2.045 55.725 2.107 ;
      RECT 55.355 1.85 55.715 1.94 ;
      RECT 55.365 1.807 55.67 2.201 ;
      RECT 55.476 1.762 55.605 2.27 ;
      RECT 55.35 3.515 55.65 3.77 ;
      RECT 55.435 3.481 55.65 3.77 ;
      RECT 55.435 3.484 55.655 3.63 ;
      RECT 55.37 3.505 55.655 3.63 ;
      RECT 55.405 3.495 55.65 3.77 ;
      RECT 55.4 3.5 55.655 3.63 ;
      RECT 55.435 3.479 55.636 3.77 ;
      RECT 55.521 3.47 55.636 3.77 ;
      RECT 55.521 3.464 55.55 3.77 ;
      RECT 55.01 3.105 55.02 3.595 ;
      RECT 54.67 3.04 54.68 3.34 ;
      RECT 55.185 3.212 55.19 3.431 ;
      RECT 55.175 3.192 55.185 3.448 ;
      RECT 55.165 3.172 55.175 3.478 ;
      RECT 55.16 3.162 55.165 3.493 ;
      RECT 55.155 3.158 55.16 3.498 ;
      RECT 55.14 3.15 55.155 3.505 ;
      RECT 55.1 3.13 55.14 3.53 ;
      RECT 55.075 3.112 55.1 3.563 ;
      RECT 55.07 3.11 55.075 3.576 ;
      RECT 55.05 3.107 55.07 3.58 ;
      RECT 55.02 3.105 55.05 3.59 ;
      RECT 54.95 3.107 55.01 3.591 ;
      RECT 54.93 3.107 54.95 3.585 ;
      RECT 54.905 3.105 54.93 3.582 ;
      RECT 54.87 3.1 54.905 3.578 ;
      RECT 54.85 3.094 54.87 3.565 ;
      RECT 54.84 3.091 54.85 3.553 ;
      RECT 54.82 3.088 54.84 3.538 ;
      RECT 54.8 3.084 54.82 3.52 ;
      RECT 54.795 3.081 54.8 3.51 ;
      RECT 54.79 3.08 54.795 3.508 ;
      RECT 54.78 3.077 54.79 3.5 ;
      RECT 54.77 3.071 54.78 3.483 ;
      RECT 54.76 3.065 54.77 3.465 ;
      RECT 54.75 3.059 54.76 3.453 ;
      RECT 54.74 3.053 54.75 3.433 ;
      RECT 54.735 3.049 54.74 3.418 ;
      RECT 54.73 3.047 54.735 3.41 ;
      RECT 54.725 3.045 54.73 3.403 ;
      RECT 54.72 3.043 54.725 3.393 ;
      RECT 54.715 3.041 54.72 3.387 ;
      RECT 54.705 3.04 54.715 3.377 ;
      RECT 54.695 3.04 54.705 3.368 ;
      RECT 54.68 3.04 54.695 3.353 ;
      RECT 54.64 3.04 54.67 3.337 ;
      RECT 54.62 3.042 54.64 3.332 ;
      RECT 54.615 3.047 54.62 3.33 ;
      RECT 54.585 3.055 54.615 3.328 ;
      RECT 54.555 3.07 54.585 3.327 ;
      RECT 54.51 3.092 54.555 3.332 ;
      RECT 54.505 3.107 54.51 3.336 ;
      RECT 54.49 3.112 54.505 3.338 ;
      RECT 54.485 3.116 54.49 3.34 ;
      RECT 54.425 3.139 54.485 3.349 ;
      RECT 54.405 3.165 54.425 3.362 ;
      RECT 54.395 3.172 54.405 3.366 ;
      RECT 54.38 3.179 54.395 3.369 ;
      RECT 54.36 3.189 54.38 3.372 ;
      RECT 54.355 3.197 54.36 3.375 ;
      RECT 54.31 3.202 54.355 3.382 ;
      RECT 54.3 3.205 54.31 3.389 ;
      RECT 54.29 3.205 54.3 3.393 ;
      RECT 54.255 3.207 54.29 3.405 ;
      RECT 54.235 3.21 54.255 3.418 ;
      RECT 54.195 3.213 54.235 3.429 ;
      RECT 54.18 3.215 54.195 3.442 ;
      RECT 54.17 3.215 54.18 3.447 ;
      RECT 54.145 3.216 54.17 3.455 ;
      RECT 54.135 3.218 54.145 3.46 ;
      RECT 54.13 3.219 54.135 3.463 ;
      RECT 54.105 3.217 54.13 3.466 ;
      RECT 54.09 3.215 54.105 3.467 ;
      RECT 54.07 3.212 54.09 3.469 ;
      RECT 54.05 3.207 54.07 3.469 ;
      RECT 53.99 3.202 54.05 3.466 ;
      RECT 53.955 3.177 53.99 3.462 ;
      RECT 53.945 3.154 53.955 3.46 ;
      RECT 53.915 3.131 53.945 3.46 ;
      RECT 53.905 3.11 53.915 3.46 ;
      RECT 53.88 3.092 53.905 3.458 ;
      RECT 53.865 3.07 53.88 3.455 ;
      RECT 53.85 3.052 53.865 3.453 ;
      RECT 53.83 3.042 53.85 3.451 ;
      RECT 53.815 3.037 53.83 3.45 ;
      RECT 53.8 3.035 53.815 3.449 ;
      RECT 53.77 3.036 53.8 3.447 ;
      RECT 53.75 3.039 53.77 3.445 ;
      RECT 53.693 3.043 53.75 3.445 ;
      RECT 53.607 3.052 53.693 3.445 ;
      RECT 53.521 3.063 53.607 3.445 ;
      RECT 53.435 3.074 53.521 3.445 ;
      RECT 53.415 3.081 53.435 3.453 ;
      RECT 53.405 3.084 53.415 3.46 ;
      RECT 53.34 3.089 53.405 3.478 ;
      RECT 53.31 3.096 53.34 3.503 ;
      RECT 53.3 3.099 53.31 3.51 ;
      RECT 53.255 3.103 53.3 3.515 ;
      RECT 53.225 3.108 53.255 3.52 ;
      RECT 53.224 3.11 53.225 3.52 ;
      RECT 53.138 3.116 53.224 3.52 ;
      RECT 53.052 3.127 53.138 3.52 ;
      RECT 52.966 3.139 53.052 3.52 ;
      RECT 52.88 3.15 52.966 3.52 ;
      RECT 52.865 3.157 52.88 3.515 ;
      RECT 52.86 3.159 52.865 3.509 ;
      RECT 52.84 3.17 52.86 3.504 ;
      RECT 52.83 3.188 52.84 3.498 ;
      RECT 52.825 3.2 52.83 3.298 ;
      RECT 55.12 1.953 55.14 2.04 ;
      RECT 55.115 1.888 55.12 2.072 ;
      RECT 55.105 1.855 55.115 2.077 ;
      RECT 55.1 1.835 55.105 2.083 ;
      RECT 55.07 1.835 55.1 2.1 ;
      RECT 55.021 1.835 55.07 2.136 ;
      RECT 54.935 1.835 55.021 2.194 ;
      RECT 54.906 1.845 54.935 2.243 ;
      RECT 54.82 1.887 54.906 2.296 ;
      RECT 54.8 1.925 54.82 2.343 ;
      RECT 54.775 1.942 54.8 2.363 ;
      RECT 54.765 1.956 54.775 2.383 ;
      RECT 54.76 1.962 54.765 2.393 ;
      RECT 54.755 1.966 54.76 2.4 ;
      RECT 54.705 1.986 54.755 2.405 ;
      RECT 54.64 2.03 54.705 2.405 ;
      RECT 54.615 2.08 54.64 2.405 ;
      RECT 54.605 2.11 54.615 2.405 ;
      RECT 54.6 2.137 54.605 2.405 ;
      RECT 54.595 2.155 54.6 2.405 ;
      RECT 54.585 2.197 54.595 2.405 ;
      RECT 54.935 2.755 55.105 2.93 ;
      RECT 54.875 2.583 54.935 2.918 ;
      RECT 54.865 2.576 54.875 2.901 ;
      RECT 54.82 2.755 55.105 2.881 ;
      RECT 54.801 2.755 55.105 2.859 ;
      RECT 54.715 2.755 55.105 2.824 ;
      RECT 54.695 2.575 54.865 2.78 ;
      RECT 54.695 2.722 55.1 2.78 ;
      RECT 54.695 2.67 55.075 2.78 ;
      RECT 54.695 2.625 55.04 2.78 ;
      RECT 54.695 2.607 55.005 2.78 ;
      RECT 54.695 2.597 55 2.78 ;
      RECT 54.415 3.555 54.605 3.78 ;
      RECT 54.405 3.556 54.61 3.775 ;
      RECT 54.405 3.558 54.62 3.755 ;
      RECT 54.405 3.562 54.625 3.74 ;
      RECT 54.405 3.549 54.575 3.775 ;
      RECT 54.405 3.552 54.6 3.775 ;
      RECT 54.415 3.548 54.575 3.78 ;
      RECT 54.501 3.546 54.575 3.78 ;
      RECT 54.125 2.797 54.295 3.035 ;
      RECT 54.125 2.797 54.381 2.949 ;
      RECT 54.125 2.797 54.385 2.859 ;
      RECT 54.175 2.57 54.395 2.838 ;
      RECT 54.17 2.587 54.4 2.811 ;
      RECT 54.135 2.745 54.4 2.811 ;
      RECT 54.155 2.595 54.295 3.035 ;
      RECT 54.145 2.677 54.405 2.794 ;
      RECT 54.14 2.725 54.405 2.794 ;
      RECT 54.145 2.635 54.4 2.811 ;
      RECT 54.17 2.572 54.395 2.838 ;
      RECT 53.735 2.547 53.905 2.745 ;
      RECT 53.735 2.547 53.95 2.72 ;
      RECT 53.805 2.49 53.975 2.678 ;
      RECT 53.78 2.505 53.975 2.678 ;
      RECT 53.395 2.551 53.425 2.745 ;
      RECT 53.39 2.523 53.395 2.745 ;
      RECT 53.36 2.497 53.39 2.747 ;
      RECT 53.335 2.455 53.36 2.75 ;
      RECT 53.325 2.427 53.335 2.752 ;
      RECT 53.29 2.407 53.325 2.754 ;
      RECT 53.225 2.392 53.29 2.76 ;
      RECT 53.175 2.39 53.225 2.766 ;
      RECT 53.152 2.392 53.175 2.771 ;
      RECT 53.066 2.403 53.152 2.777 ;
      RECT 52.98 2.421 53.066 2.787 ;
      RECT 52.965 2.432 52.98 2.793 ;
      RECT 52.895 2.455 52.965 2.799 ;
      RECT 52.84 2.487 52.895 2.807 ;
      RECT 52.8 2.51 52.84 2.813 ;
      RECT 52.786 2.523 52.8 2.816 ;
      RECT 52.7 2.545 52.786 2.822 ;
      RECT 52.685 2.57 52.7 2.828 ;
      RECT 52.645 2.585 52.685 2.832 ;
      RECT 52.595 2.6 52.645 2.837 ;
      RECT 52.57 2.607 52.595 2.841 ;
      RECT 52.51 2.602 52.57 2.845 ;
      RECT 52.495 2.593 52.51 2.849 ;
      RECT 52.425 2.583 52.495 2.845 ;
      RECT 52.4 2.575 52.42 2.835 ;
      RECT 52.341 2.575 52.4 2.813 ;
      RECT 52.255 2.575 52.341 2.77 ;
      RECT 52.42 2.575 52.425 2.84 ;
      RECT 53.115 1.806 53.285 2.14 ;
      RECT 53.085 1.806 53.285 2.135 ;
      RECT 53.025 1.773 53.085 2.123 ;
      RECT 53.025 1.829 53.295 2.118 ;
      RECT 53 1.829 53.295 2.112 ;
      RECT 52.995 1.77 53.025 2.109 ;
      RECT 52.98 1.776 53.115 2.107 ;
      RECT 52.975 1.784 53.2 2.095 ;
      RECT 52.975 1.836 53.31 2.048 ;
      RECT 52.96 1.792 53.2 2.043 ;
      RECT 52.96 1.862 53.32 1.984 ;
      RECT 52.93 1.812 53.285 1.945 ;
      RECT 52.93 1.902 53.33 1.941 ;
      RECT 52.98 1.781 53.2 2.107 ;
      RECT 52.32 2.111 52.375 2.375 ;
      RECT 52.32 2.111 52.44 2.374 ;
      RECT 52.32 2.111 52.465 2.373 ;
      RECT 52.32 2.111 52.53 2.372 ;
      RECT 52.465 2.077 52.545 2.371 ;
      RECT 52.28 2.121 52.69 2.37 ;
      RECT 52.32 2.118 52.69 2.37 ;
      RECT 52.28 2.126 52.695 2.363 ;
      RECT 52.265 2.128 52.695 2.362 ;
      RECT 52.265 2.135 52.7 2.358 ;
      RECT 52.245 2.134 52.695 2.354 ;
      RECT 52.245 2.142 52.705 2.353 ;
      RECT 52.24 2.139 52.7 2.349 ;
      RECT 52.24 2.152 52.715 2.348 ;
      RECT 52.225 2.142 52.705 2.347 ;
      RECT 52.19 2.155 52.715 2.34 ;
      RECT 52.375 2.11 52.685 2.37 ;
      RECT 52.375 2.095 52.635 2.37 ;
      RECT 52.44 2.082 52.57 2.37 ;
      RECT 51.985 3.171 52 3.564 ;
      RECT 51.95 3.176 52 3.563 ;
      RECT 51.985 3.175 52.045 3.562 ;
      RECT 51.93 3.186 52.045 3.561 ;
      RECT 51.945 3.182 52.045 3.561 ;
      RECT 51.91 3.192 52.12 3.558 ;
      RECT 51.91 3.211 52.165 3.556 ;
      RECT 51.91 3.218 52.17 3.553 ;
      RECT 51.895 3.195 52.12 3.55 ;
      RECT 51.875 3.2 52.12 3.543 ;
      RECT 51.87 3.204 52.12 3.539 ;
      RECT 51.87 3.221 52.18 3.538 ;
      RECT 51.85 3.215 52.165 3.534 ;
      RECT 51.85 3.224 52.185 3.528 ;
      RECT 51.845 3.23 52.185 3.3 ;
      RECT 51.91 3.19 52.045 3.558 ;
      RECT 51.785 2.553 51.985 2.865 ;
      RECT 51.86 2.531 51.985 2.865 ;
      RECT 51.8 2.55 51.99 2.85 ;
      RECT 51.77 2.561 51.99 2.848 ;
      RECT 51.785 2.556 51.995 2.814 ;
      RECT 51.77 2.66 52 2.781 ;
      RECT 51.8 2.532 51.985 2.865 ;
      RECT 51.86 2.51 51.96 2.865 ;
      RECT 51.885 2.507 51.96 2.865 ;
      RECT 51.885 2.502 51.905 2.865 ;
      RECT 51.29 2.57 51.465 2.745 ;
      RECT 51.285 2.57 51.465 2.743 ;
      RECT 51.26 2.57 51.465 2.738 ;
      RECT 51.205 2.55 51.375 2.728 ;
      RECT 51.205 2.557 51.44 2.728 ;
      RECT 51.29 3.237 51.305 3.42 ;
      RECT 51.28 3.215 51.29 3.42 ;
      RECT 51.265 3.195 51.28 3.42 ;
      RECT 51.255 3.17 51.265 3.42 ;
      RECT 51.225 3.135 51.255 3.42 ;
      RECT 51.19 3.075 51.225 3.42 ;
      RECT 51.185 3.037 51.19 3.42 ;
      RECT 51.135 2.988 51.185 3.42 ;
      RECT 51.125 2.938 51.135 3.408 ;
      RECT 51.11 2.917 51.125 3.368 ;
      RECT 51.09 2.885 51.11 3.318 ;
      RECT 51.065 2.841 51.09 3.258 ;
      RECT 51.06 2.813 51.065 3.213 ;
      RECT 51.055 2.804 51.06 3.199 ;
      RECT 51.05 2.797 51.055 3.186 ;
      RECT 51.045 2.792 51.05 3.175 ;
      RECT 51.04 2.777 51.045 3.165 ;
      RECT 51.035 2.755 51.04 3.152 ;
      RECT 51.025 2.715 51.035 3.127 ;
      RECT 51 2.645 51.025 3.083 ;
      RECT 50.995 2.585 51 3.048 ;
      RECT 50.98 2.565 50.995 3.015 ;
      RECT 50.975 2.565 50.98 2.99 ;
      RECT 50.945 2.565 50.975 2.945 ;
      RECT 50.9 2.565 50.945 2.885 ;
      RECT 50.825 2.565 50.9 2.833 ;
      RECT 50.82 2.565 50.825 2.798 ;
      RECT 50.815 2.565 50.82 2.788 ;
      RECT 50.81 2.565 50.815 2.768 ;
      RECT 51.075 1.785 51.245 2.255 ;
      RECT 51.02 1.778 51.215 2.239 ;
      RECT 51.02 1.792 51.25 2.238 ;
      RECT 51.005 1.793 51.25 2.219 ;
      RECT 51 1.811 51.25 2.205 ;
      RECT 51.005 1.794 51.255 2.203 ;
      RECT 50.99 1.825 51.255 2.188 ;
      RECT 51.005 1.8 51.26 2.173 ;
      RECT 50.985 1.84 51.26 2.17 ;
      RECT 51 1.812 51.265 2.155 ;
      RECT 51 1.824 51.27 2.135 ;
      RECT 50.985 1.84 51.275 2.118 ;
      RECT 50.985 1.85 51.28 1.973 ;
      RECT 50.98 1.85 51.28 1.93 ;
      RECT 50.98 1.865 51.285 1.908 ;
      RECT 51.075 1.775 51.215 2.255 ;
      RECT 51.075 1.773 51.185 2.255 ;
      RECT 51.161 1.77 51.185 2.255 ;
      RECT 50.82 3.437 50.825 3.483 ;
      RECT 50.81 3.285 50.82 3.507 ;
      RECT 50.805 3.13 50.81 3.532 ;
      RECT 50.79 3.092 50.805 3.543 ;
      RECT 50.785 3.075 50.79 3.55 ;
      RECT 50.775 3.063 50.785 3.557 ;
      RECT 50.77 3.054 50.775 3.559 ;
      RECT 50.765 3.052 50.77 3.563 ;
      RECT 50.72 3.043 50.765 3.578 ;
      RECT 50.715 3.035 50.72 3.592 ;
      RECT 50.71 3.032 50.715 3.596 ;
      RECT 50.695 3.027 50.71 3.604 ;
      RECT 50.64 3.017 50.695 3.615 ;
      RECT 50.605 3.005 50.64 3.616 ;
      RECT 50.596 3 50.605 3.61 ;
      RECT 50.51 3 50.596 3.6 ;
      RECT 50.48 3 50.51 3.578 ;
      RECT 50.47 3 50.475 3.558 ;
      RECT 50.465 3 50.47 3.52 ;
      RECT 50.46 3 50.465 3.478 ;
      RECT 50.455 3 50.46 3.438 ;
      RECT 50.45 3 50.455 3.368 ;
      RECT 50.44 3 50.45 3.29 ;
      RECT 50.435 3 50.44 3.19 ;
      RECT 50.475 3 50.48 3.56 ;
      RECT 49.97 3.082 50.06 3.56 ;
      RECT 49.955 3.085 50.075 3.558 ;
      RECT 49.97 3.084 50.075 3.558 ;
      RECT 49.935 3.091 50.1 3.548 ;
      RECT 49.955 3.085 50.1 3.548 ;
      RECT 49.92 3.097 50.1 3.536 ;
      RECT 49.955 3.088 50.15 3.529 ;
      RECT 49.906 3.105 50.15 3.527 ;
      RECT 49.935 3.095 50.16 3.515 ;
      RECT 49.906 3.116 50.19 3.506 ;
      RECT 49.82 3.14 50.19 3.5 ;
      RECT 49.82 3.153 50.23 3.483 ;
      RECT 49.815 3.175 50.23 3.476 ;
      RECT 49.785 3.19 50.23 3.466 ;
      RECT 49.78 3.201 50.23 3.456 ;
      RECT 49.75 3.214 50.23 3.447 ;
      RECT 49.735 3.232 50.23 3.436 ;
      RECT 49.71 3.245 50.23 3.426 ;
      RECT 49.97 3.081 49.98 3.56 ;
      RECT 50.016 2.505 50.055 2.75 ;
      RECT 49.93 2.505 50.065 2.748 ;
      RECT 49.815 2.53 50.065 2.745 ;
      RECT 49.815 2.53 50.07 2.743 ;
      RECT 49.815 2.53 50.085 2.738 ;
      RECT 49.921 2.505 50.1 2.718 ;
      RECT 49.835 2.513 50.1 2.718 ;
      RECT 49.505 1.865 49.675 2.3 ;
      RECT 49.495 1.899 49.675 2.283 ;
      RECT 49.575 1.835 49.745 2.27 ;
      RECT 49.48 1.91 49.745 2.248 ;
      RECT 49.575 1.845 49.75 2.238 ;
      RECT 49.505 1.897 49.78 2.223 ;
      RECT 49.465 1.923 49.78 2.208 ;
      RECT 49.465 1.965 49.79 2.188 ;
      RECT 49.46 1.99 49.795 2.17 ;
      RECT 49.46 2 49.8 2.155 ;
      RECT 49.455 1.937 49.78 2.153 ;
      RECT 49.455 2.01 49.805 2.138 ;
      RECT 49.45 1.947 49.78 2.135 ;
      RECT 49.445 2.031 49.81 2.118 ;
      RECT 49.445 2.063 49.815 2.098 ;
      RECT 49.44 1.977 49.79 2.09 ;
      RECT 49.445 1.962 49.78 2.118 ;
      RECT 49.46 1.932 49.78 2.17 ;
      RECT 49.305 2.519 49.53 2.775 ;
      RECT 49.305 2.552 49.55 2.765 ;
      RECT 49.27 2.552 49.55 2.763 ;
      RECT 49.27 2.565 49.555 2.753 ;
      RECT 49.27 2.585 49.565 2.745 ;
      RECT 49.27 2.682 49.57 2.738 ;
      RECT 49.25 2.43 49.38 2.728 ;
      RECT 49.205 2.585 49.565 2.67 ;
      RECT 49.195 2.43 49.38 2.615 ;
      RECT 49.195 2.462 49.466 2.615 ;
      RECT 49.16 2.992 49.18 3.17 ;
      RECT 49.125 2.945 49.16 3.17 ;
      RECT 49.11 2.885 49.125 3.17 ;
      RECT 49.085 2.832 49.11 3.17 ;
      RECT 49.07 2.785 49.085 3.17 ;
      RECT 49.05 2.762 49.07 3.17 ;
      RECT 49.025 2.727 49.05 3.17 ;
      RECT 49.015 2.573 49.025 3.17 ;
      RECT 48.985 2.568 49.015 3.161 ;
      RECT 48.98 2.565 48.985 3.151 ;
      RECT 48.965 2.565 48.98 3.125 ;
      RECT 48.96 2.565 48.965 3.088 ;
      RECT 48.935 2.565 48.96 3.04 ;
      RECT 48.915 2.565 48.935 2.965 ;
      RECT 48.905 2.565 48.915 2.925 ;
      RECT 48.9 2.565 48.905 2.9 ;
      RECT 48.895 2.565 48.9 2.883 ;
      RECT 48.89 2.565 48.895 2.865 ;
      RECT 48.885 2.566 48.89 2.855 ;
      RECT 48.875 2.568 48.885 2.823 ;
      RECT 48.865 2.57 48.875 2.79 ;
      RECT 48.855 2.573 48.865 2.763 ;
      RECT 49.18 3 49.405 3.17 ;
      RECT 48.51 1.812 48.68 2.265 ;
      RECT 48.51 1.812 48.77 2.231 ;
      RECT 48.51 1.812 48.8 2.215 ;
      RECT 48.51 1.812 48.83 2.188 ;
      RECT 48.766 1.79 48.845 2.17 ;
      RECT 48.545 1.797 48.85 2.155 ;
      RECT 48.545 1.805 48.86 2.118 ;
      RECT 48.505 1.832 48.86 2.09 ;
      RECT 48.49 1.845 48.86 2.055 ;
      RECT 48.51 1.82 48.88 2.045 ;
      RECT 48.485 1.885 48.88 2.015 ;
      RECT 48.485 1.915 48.885 1.998 ;
      RECT 48.48 1.945 48.885 1.985 ;
      RECT 48.545 1.794 48.845 2.17 ;
      RECT 48.68 1.791 48.766 2.249 ;
      RECT 48.631 1.792 48.845 2.17 ;
      RECT 48.775 3.452 48.82 3.645 ;
      RECT 48.765 3.422 48.775 3.645 ;
      RECT 48.76 3.407 48.765 3.645 ;
      RECT 48.72 3.317 48.76 3.645 ;
      RECT 48.715 3.23 48.72 3.645 ;
      RECT 48.705 3.2 48.715 3.645 ;
      RECT 48.7 3.16 48.705 3.645 ;
      RECT 48.69 3.122 48.7 3.645 ;
      RECT 48.685 3.087 48.69 3.645 ;
      RECT 48.665 3.04 48.685 3.645 ;
      RECT 48.65 2.965 48.665 3.645 ;
      RECT 48.645 2.92 48.65 3.64 ;
      RECT 48.64 2.9 48.645 3.613 ;
      RECT 48.635 2.88 48.64 3.598 ;
      RECT 48.63 2.855 48.635 3.578 ;
      RECT 48.625 2.833 48.63 3.563 ;
      RECT 48.62 2.811 48.625 3.545 ;
      RECT 48.615 2.79 48.62 3.535 ;
      RECT 48.605 2.762 48.615 3.505 ;
      RECT 48.595 2.725 48.605 3.473 ;
      RECT 48.585 2.685 48.595 3.44 ;
      RECT 48.575 2.663 48.585 3.41 ;
      RECT 48.545 2.615 48.575 3.342 ;
      RECT 48.53 2.575 48.545 3.269 ;
      RECT 48.52 2.575 48.53 3.235 ;
      RECT 48.515 2.575 48.52 3.21 ;
      RECT 48.51 2.575 48.515 3.195 ;
      RECT 48.505 2.575 48.51 3.173 ;
      RECT 48.5 2.575 48.505 3.16 ;
      RECT 48.485 2.575 48.5 3.125 ;
      RECT 48.465 2.575 48.485 3.065 ;
      RECT 48.455 2.575 48.465 3.015 ;
      RECT 48.435 2.575 48.455 2.963 ;
      RECT 48.415 2.575 48.435 2.92 ;
      RECT 48.405 2.575 48.415 2.908 ;
      RECT 48.375 2.575 48.405 2.895 ;
      RECT 48.345 2.596 48.375 2.875 ;
      RECT 48.335 2.624 48.345 2.855 ;
      RECT 48.32 2.641 48.335 2.823 ;
      RECT 48.315 2.655 48.32 2.79 ;
      RECT 48.31 2.663 48.315 2.763 ;
      RECT 48.305 2.671 48.31 2.725 ;
      RECT 48.31 3.195 48.315 3.53 ;
      RECT 48.275 3.182 48.31 3.529 ;
      RECT 48.205 3.122 48.275 3.528 ;
      RECT 48.125 3.065 48.205 3.527 ;
      RECT 47.99 3.025 48.125 3.526 ;
      RECT 47.99 3.212 48.325 3.515 ;
      RECT 47.95 3.212 48.325 3.505 ;
      RECT 47.95 3.23 48.33 3.5 ;
      RECT 47.95 3.32 48.335 3.49 ;
      RECT 47.945 3.015 48.11 3.47 ;
      RECT 47.94 3.015 48.11 3.213 ;
      RECT 47.94 3.172 48.305 3.213 ;
      RECT 47.94 3.16 48.3 3.213 ;
      RECT 46.64 1.74 46.81 2.935 ;
      RECT 46.64 1.74 47.105 1.91 ;
      RECT 46.64 6.97 47.105 7.14 ;
      RECT 46.64 5.945 46.81 7.14 ;
      RECT 45.65 1.74 45.82 2.935 ;
      RECT 45.65 1.74 46.115 1.91 ;
      RECT 45.65 6.97 46.115 7.14 ;
      RECT 45.65 5.945 45.82 7.14 ;
      RECT 43.795 2.635 43.965 3.865 ;
      RECT 43.85 0.855 44.02 2.805 ;
      RECT 43.795 0.575 43.965 1.025 ;
      RECT 43.795 7.855 43.965 8.305 ;
      RECT 43.85 6.075 44.02 8.025 ;
      RECT 43.795 5.015 43.965 6.245 ;
      RECT 43.275 0.575 43.445 3.865 ;
      RECT 43.275 2.075 43.68 2.405 ;
      RECT 43.275 1.235 43.68 1.565 ;
      RECT 43.275 5.015 43.445 8.305 ;
      RECT 43.275 7.315 43.68 7.645 ;
      RECT 43.275 6.475 43.68 6.805 ;
      RECT 40.61 1.975 41.34 2.215 ;
      RECT 41.152 1.77 41.34 2.215 ;
      RECT 40.98 1.782 41.355 2.209 ;
      RECT 40.895 1.797 41.375 2.194 ;
      RECT 40.895 1.812 41.38 2.184 ;
      RECT 40.85 1.832 41.395 2.176 ;
      RECT 40.827 1.867 41.41 2.13 ;
      RECT 40.741 1.89 41.415 2.09 ;
      RECT 40.741 1.908 41.425 2.06 ;
      RECT 40.61 1.977 41.43 2.023 ;
      RECT 40.655 1.92 41.425 2.06 ;
      RECT 40.741 1.872 41.41 2.13 ;
      RECT 40.827 1.841 41.395 2.176 ;
      RECT 40.85 1.822 41.38 2.184 ;
      RECT 40.895 1.795 41.355 2.209 ;
      RECT 40.98 1.777 41.34 2.215 ;
      RECT 41.066 1.771 41.34 2.215 ;
      RECT 41.152 1.766 41.285 2.215 ;
      RECT 41.238 1.761 41.285 2.215 ;
      RECT 40.93 2.659 41.1 3.045 ;
      RECT 40.925 2.659 41.1 3.04 ;
      RECT 40.9 2.659 41.1 3.005 ;
      RECT 40.9 2.687 41.11 2.995 ;
      RECT 40.88 2.687 41.11 2.955 ;
      RECT 40.875 2.687 41.11 2.928 ;
      RECT 40.875 2.705 41.115 2.92 ;
      RECT 40.82 2.705 41.115 2.855 ;
      RECT 40.82 2.722 41.125 2.838 ;
      RECT 40.81 2.722 41.125 2.778 ;
      RECT 40.81 2.739 41.13 2.775 ;
      RECT 40.805 2.575 40.975 2.753 ;
      RECT 40.805 2.609 41.061 2.753 ;
      RECT 40.8 3.375 40.805 3.388 ;
      RECT 40.795 3.27 40.8 3.393 ;
      RECT 40.77 3.13 40.795 3.408 ;
      RECT 40.735 3.081 40.77 3.44 ;
      RECT 40.73 3.049 40.735 3.46 ;
      RECT 40.725 3.04 40.73 3.46 ;
      RECT 40.645 3.005 40.725 3.46 ;
      RECT 40.582 2.975 40.645 3.46 ;
      RECT 40.496 2.963 40.582 3.46 ;
      RECT 40.41 2.949 40.496 3.46 ;
      RECT 40.33 2.936 40.41 3.446 ;
      RECT 40.295 2.928 40.33 3.426 ;
      RECT 40.285 2.925 40.295 3.417 ;
      RECT 40.255 2.92 40.285 3.404 ;
      RECT 40.205 2.895 40.255 3.38 ;
      RECT 40.191 2.869 40.205 3.362 ;
      RECT 40.105 2.829 40.191 3.338 ;
      RECT 40.06 2.777 40.105 3.307 ;
      RECT 40.05 2.752 40.06 3.294 ;
      RECT 40.045 2.533 40.05 2.555 ;
      RECT 40.04 2.735 40.05 3.29 ;
      RECT 40.04 2.531 40.045 2.645 ;
      RECT 40.03 2.527 40.04 3.286 ;
      RECT 39.986 2.525 40.03 3.274 ;
      RECT 39.9 2.525 39.986 3.245 ;
      RECT 39.87 2.525 39.9 3.218 ;
      RECT 39.855 2.525 39.87 3.206 ;
      RECT 39.815 2.537 39.855 3.191 ;
      RECT 39.795 2.556 39.815 3.17 ;
      RECT 39.785 2.566 39.795 3.154 ;
      RECT 39.775 2.572 39.785 3.143 ;
      RECT 39.755 2.582 39.775 3.126 ;
      RECT 39.75 2.591 39.755 3.113 ;
      RECT 39.745 2.595 39.75 3.063 ;
      RECT 39.735 2.601 39.745 2.98 ;
      RECT 39.73 2.605 39.735 2.894 ;
      RECT 39.725 2.625 39.73 2.831 ;
      RECT 39.72 2.648 39.725 2.778 ;
      RECT 39.715 2.666 39.72 2.723 ;
      RECT 40.325 2.485 40.495 2.745 ;
      RECT 40.495 2.45 40.54 2.731 ;
      RECT 40.456 2.452 40.545 2.714 ;
      RECT 40.345 2.469 40.631 2.685 ;
      RECT 40.345 2.484 40.635 2.657 ;
      RECT 40.345 2.465 40.545 2.714 ;
      RECT 40.37 2.453 40.495 2.745 ;
      RECT 40.456 2.451 40.54 2.731 ;
      RECT 39.51 1.84 39.68 2.33 ;
      RECT 39.51 1.84 39.715 2.31 ;
      RECT 39.645 1.76 39.755 2.27 ;
      RECT 39.626 1.764 39.775 2.24 ;
      RECT 39.54 1.772 39.795 2.223 ;
      RECT 39.54 1.778 39.8 2.213 ;
      RECT 39.54 1.787 39.82 2.201 ;
      RECT 39.515 1.812 39.85 2.179 ;
      RECT 39.515 1.832 39.855 2.159 ;
      RECT 39.51 1.845 39.865 2.139 ;
      RECT 39.51 1.912 39.87 2.12 ;
      RECT 39.51 2.045 39.875 2.107 ;
      RECT 39.505 1.85 39.865 1.94 ;
      RECT 39.515 1.807 39.82 2.201 ;
      RECT 39.626 1.762 39.755 2.27 ;
      RECT 39.5 3.515 39.8 3.77 ;
      RECT 39.585 3.481 39.8 3.77 ;
      RECT 39.585 3.484 39.805 3.63 ;
      RECT 39.52 3.505 39.805 3.63 ;
      RECT 39.555 3.495 39.8 3.77 ;
      RECT 39.55 3.5 39.805 3.63 ;
      RECT 39.585 3.479 39.786 3.77 ;
      RECT 39.671 3.47 39.786 3.77 ;
      RECT 39.671 3.464 39.7 3.77 ;
      RECT 39.16 3.105 39.17 3.595 ;
      RECT 38.82 3.04 38.83 3.34 ;
      RECT 39.335 3.212 39.34 3.431 ;
      RECT 39.325 3.192 39.335 3.448 ;
      RECT 39.315 3.172 39.325 3.478 ;
      RECT 39.31 3.162 39.315 3.493 ;
      RECT 39.305 3.158 39.31 3.498 ;
      RECT 39.29 3.15 39.305 3.505 ;
      RECT 39.25 3.13 39.29 3.53 ;
      RECT 39.225 3.112 39.25 3.563 ;
      RECT 39.22 3.11 39.225 3.576 ;
      RECT 39.2 3.107 39.22 3.58 ;
      RECT 39.17 3.105 39.2 3.59 ;
      RECT 39.1 3.107 39.16 3.591 ;
      RECT 39.08 3.107 39.1 3.585 ;
      RECT 39.055 3.105 39.08 3.582 ;
      RECT 39.02 3.1 39.055 3.578 ;
      RECT 39 3.094 39.02 3.565 ;
      RECT 38.99 3.091 39 3.553 ;
      RECT 38.97 3.088 38.99 3.538 ;
      RECT 38.95 3.084 38.97 3.52 ;
      RECT 38.945 3.081 38.95 3.51 ;
      RECT 38.94 3.08 38.945 3.508 ;
      RECT 38.93 3.077 38.94 3.5 ;
      RECT 38.92 3.071 38.93 3.483 ;
      RECT 38.91 3.065 38.92 3.465 ;
      RECT 38.9 3.059 38.91 3.453 ;
      RECT 38.89 3.053 38.9 3.433 ;
      RECT 38.885 3.049 38.89 3.418 ;
      RECT 38.88 3.047 38.885 3.41 ;
      RECT 38.875 3.045 38.88 3.403 ;
      RECT 38.87 3.043 38.875 3.393 ;
      RECT 38.865 3.041 38.87 3.387 ;
      RECT 38.855 3.04 38.865 3.377 ;
      RECT 38.845 3.04 38.855 3.368 ;
      RECT 38.83 3.04 38.845 3.353 ;
      RECT 38.79 3.04 38.82 3.337 ;
      RECT 38.77 3.042 38.79 3.332 ;
      RECT 38.765 3.047 38.77 3.33 ;
      RECT 38.735 3.055 38.765 3.328 ;
      RECT 38.705 3.07 38.735 3.327 ;
      RECT 38.66 3.092 38.705 3.332 ;
      RECT 38.655 3.107 38.66 3.336 ;
      RECT 38.64 3.112 38.655 3.338 ;
      RECT 38.635 3.116 38.64 3.34 ;
      RECT 38.575 3.139 38.635 3.349 ;
      RECT 38.555 3.165 38.575 3.362 ;
      RECT 38.545 3.172 38.555 3.366 ;
      RECT 38.53 3.179 38.545 3.369 ;
      RECT 38.51 3.189 38.53 3.372 ;
      RECT 38.505 3.197 38.51 3.375 ;
      RECT 38.46 3.202 38.505 3.382 ;
      RECT 38.45 3.205 38.46 3.389 ;
      RECT 38.44 3.205 38.45 3.393 ;
      RECT 38.405 3.207 38.44 3.405 ;
      RECT 38.385 3.21 38.405 3.418 ;
      RECT 38.345 3.213 38.385 3.429 ;
      RECT 38.33 3.215 38.345 3.442 ;
      RECT 38.32 3.215 38.33 3.447 ;
      RECT 38.295 3.216 38.32 3.455 ;
      RECT 38.285 3.218 38.295 3.46 ;
      RECT 38.28 3.219 38.285 3.463 ;
      RECT 38.255 3.217 38.28 3.466 ;
      RECT 38.24 3.215 38.255 3.467 ;
      RECT 38.22 3.212 38.24 3.469 ;
      RECT 38.2 3.207 38.22 3.469 ;
      RECT 38.14 3.202 38.2 3.466 ;
      RECT 38.105 3.177 38.14 3.462 ;
      RECT 38.095 3.154 38.105 3.46 ;
      RECT 38.065 3.131 38.095 3.46 ;
      RECT 38.055 3.11 38.065 3.46 ;
      RECT 38.03 3.092 38.055 3.458 ;
      RECT 38.015 3.07 38.03 3.455 ;
      RECT 38 3.052 38.015 3.453 ;
      RECT 37.98 3.042 38 3.451 ;
      RECT 37.965 3.037 37.98 3.45 ;
      RECT 37.95 3.035 37.965 3.449 ;
      RECT 37.92 3.036 37.95 3.447 ;
      RECT 37.9 3.039 37.92 3.445 ;
      RECT 37.843 3.043 37.9 3.445 ;
      RECT 37.757 3.052 37.843 3.445 ;
      RECT 37.671 3.063 37.757 3.445 ;
      RECT 37.585 3.074 37.671 3.445 ;
      RECT 37.565 3.081 37.585 3.453 ;
      RECT 37.555 3.084 37.565 3.46 ;
      RECT 37.49 3.089 37.555 3.478 ;
      RECT 37.46 3.096 37.49 3.503 ;
      RECT 37.45 3.099 37.46 3.51 ;
      RECT 37.405 3.103 37.45 3.515 ;
      RECT 37.375 3.108 37.405 3.52 ;
      RECT 37.374 3.11 37.375 3.52 ;
      RECT 37.288 3.116 37.374 3.52 ;
      RECT 37.202 3.127 37.288 3.52 ;
      RECT 37.116 3.139 37.202 3.52 ;
      RECT 37.03 3.15 37.116 3.52 ;
      RECT 37.015 3.157 37.03 3.515 ;
      RECT 37.01 3.159 37.015 3.509 ;
      RECT 36.99 3.17 37.01 3.504 ;
      RECT 36.98 3.188 36.99 3.498 ;
      RECT 36.975 3.2 36.98 3.298 ;
      RECT 39.27 1.953 39.29 2.04 ;
      RECT 39.265 1.888 39.27 2.072 ;
      RECT 39.255 1.855 39.265 2.077 ;
      RECT 39.25 1.835 39.255 2.083 ;
      RECT 39.22 1.835 39.25 2.1 ;
      RECT 39.171 1.835 39.22 2.136 ;
      RECT 39.085 1.835 39.171 2.194 ;
      RECT 39.056 1.845 39.085 2.243 ;
      RECT 38.97 1.887 39.056 2.296 ;
      RECT 38.95 1.925 38.97 2.343 ;
      RECT 38.925 1.942 38.95 2.363 ;
      RECT 38.915 1.956 38.925 2.383 ;
      RECT 38.91 1.962 38.915 2.393 ;
      RECT 38.905 1.966 38.91 2.4 ;
      RECT 38.855 1.986 38.905 2.405 ;
      RECT 38.79 2.03 38.855 2.405 ;
      RECT 38.765 2.08 38.79 2.405 ;
      RECT 38.755 2.11 38.765 2.405 ;
      RECT 38.75 2.137 38.755 2.405 ;
      RECT 38.745 2.155 38.75 2.405 ;
      RECT 38.735 2.197 38.745 2.405 ;
      RECT 39.085 2.755 39.255 2.93 ;
      RECT 39.025 2.583 39.085 2.918 ;
      RECT 39.015 2.576 39.025 2.901 ;
      RECT 38.97 2.755 39.255 2.881 ;
      RECT 38.951 2.755 39.255 2.859 ;
      RECT 38.865 2.755 39.255 2.824 ;
      RECT 38.845 2.575 39.015 2.78 ;
      RECT 38.845 2.722 39.25 2.78 ;
      RECT 38.845 2.67 39.225 2.78 ;
      RECT 38.845 2.625 39.19 2.78 ;
      RECT 38.845 2.607 39.155 2.78 ;
      RECT 38.845 2.597 39.15 2.78 ;
      RECT 38.565 3.555 38.755 3.78 ;
      RECT 38.555 3.556 38.76 3.775 ;
      RECT 38.555 3.558 38.77 3.755 ;
      RECT 38.555 3.562 38.775 3.74 ;
      RECT 38.555 3.549 38.725 3.775 ;
      RECT 38.555 3.552 38.75 3.775 ;
      RECT 38.565 3.548 38.725 3.78 ;
      RECT 38.651 3.546 38.725 3.78 ;
      RECT 38.275 2.797 38.445 3.035 ;
      RECT 38.275 2.797 38.531 2.949 ;
      RECT 38.275 2.797 38.535 2.859 ;
      RECT 38.325 2.57 38.545 2.838 ;
      RECT 38.32 2.587 38.55 2.811 ;
      RECT 38.285 2.745 38.55 2.811 ;
      RECT 38.305 2.595 38.445 3.035 ;
      RECT 38.295 2.677 38.555 2.794 ;
      RECT 38.29 2.725 38.555 2.794 ;
      RECT 38.295 2.635 38.55 2.811 ;
      RECT 38.32 2.572 38.545 2.838 ;
      RECT 37.885 2.547 38.055 2.745 ;
      RECT 37.885 2.547 38.1 2.72 ;
      RECT 37.955 2.49 38.125 2.678 ;
      RECT 37.93 2.505 38.125 2.678 ;
      RECT 37.545 2.551 37.575 2.745 ;
      RECT 37.54 2.523 37.545 2.745 ;
      RECT 37.51 2.497 37.54 2.747 ;
      RECT 37.485 2.455 37.51 2.75 ;
      RECT 37.475 2.427 37.485 2.752 ;
      RECT 37.44 2.407 37.475 2.754 ;
      RECT 37.375 2.392 37.44 2.76 ;
      RECT 37.325 2.39 37.375 2.766 ;
      RECT 37.302 2.392 37.325 2.771 ;
      RECT 37.216 2.403 37.302 2.777 ;
      RECT 37.13 2.421 37.216 2.787 ;
      RECT 37.115 2.432 37.13 2.793 ;
      RECT 37.045 2.455 37.115 2.799 ;
      RECT 36.99 2.487 37.045 2.807 ;
      RECT 36.95 2.51 36.99 2.813 ;
      RECT 36.936 2.523 36.95 2.816 ;
      RECT 36.85 2.545 36.936 2.822 ;
      RECT 36.835 2.57 36.85 2.828 ;
      RECT 36.795 2.585 36.835 2.832 ;
      RECT 36.745 2.6 36.795 2.837 ;
      RECT 36.72 2.607 36.745 2.841 ;
      RECT 36.66 2.602 36.72 2.845 ;
      RECT 36.645 2.593 36.66 2.849 ;
      RECT 36.575 2.583 36.645 2.845 ;
      RECT 36.55 2.575 36.57 2.835 ;
      RECT 36.491 2.575 36.55 2.813 ;
      RECT 36.405 2.575 36.491 2.77 ;
      RECT 36.57 2.575 36.575 2.84 ;
      RECT 37.265 1.806 37.435 2.14 ;
      RECT 37.235 1.806 37.435 2.135 ;
      RECT 37.175 1.773 37.235 2.123 ;
      RECT 37.175 1.829 37.445 2.118 ;
      RECT 37.15 1.829 37.445 2.112 ;
      RECT 37.145 1.77 37.175 2.109 ;
      RECT 37.13 1.776 37.265 2.107 ;
      RECT 37.125 1.784 37.35 2.095 ;
      RECT 37.125 1.836 37.46 2.048 ;
      RECT 37.11 1.792 37.35 2.043 ;
      RECT 37.11 1.862 37.47 1.984 ;
      RECT 37.08 1.812 37.435 1.945 ;
      RECT 37.08 1.902 37.48 1.941 ;
      RECT 37.13 1.781 37.35 2.107 ;
      RECT 36.47 2.111 36.525 2.375 ;
      RECT 36.47 2.111 36.59 2.374 ;
      RECT 36.47 2.111 36.615 2.373 ;
      RECT 36.47 2.111 36.68 2.372 ;
      RECT 36.615 2.077 36.695 2.371 ;
      RECT 36.43 2.121 36.84 2.37 ;
      RECT 36.47 2.118 36.84 2.37 ;
      RECT 36.43 2.126 36.845 2.363 ;
      RECT 36.415 2.128 36.845 2.362 ;
      RECT 36.415 2.135 36.85 2.358 ;
      RECT 36.395 2.134 36.845 2.354 ;
      RECT 36.395 2.142 36.855 2.353 ;
      RECT 36.39 2.139 36.85 2.349 ;
      RECT 36.39 2.152 36.865 2.348 ;
      RECT 36.375 2.142 36.855 2.347 ;
      RECT 36.34 2.155 36.865 2.34 ;
      RECT 36.525 2.11 36.835 2.37 ;
      RECT 36.525 2.095 36.785 2.37 ;
      RECT 36.59 2.082 36.72 2.37 ;
      RECT 36.135 3.171 36.15 3.564 ;
      RECT 36.1 3.176 36.15 3.563 ;
      RECT 36.135 3.175 36.195 3.562 ;
      RECT 36.08 3.186 36.195 3.561 ;
      RECT 36.095 3.182 36.195 3.561 ;
      RECT 36.06 3.192 36.27 3.558 ;
      RECT 36.06 3.211 36.315 3.556 ;
      RECT 36.06 3.218 36.32 3.553 ;
      RECT 36.045 3.195 36.27 3.55 ;
      RECT 36.025 3.2 36.27 3.543 ;
      RECT 36.02 3.204 36.27 3.539 ;
      RECT 36.02 3.221 36.33 3.538 ;
      RECT 36 3.215 36.315 3.534 ;
      RECT 36 3.224 36.335 3.528 ;
      RECT 35.995 3.23 36.335 3.3 ;
      RECT 36.06 3.19 36.195 3.558 ;
      RECT 35.935 2.553 36.135 2.865 ;
      RECT 36.01 2.531 36.135 2.865 ;
      RECT 35.95 2.55 36.14 2.85 ;
      RECT 35.92 2.561 36.14 2.848 ;
      RECT 35.935 2.556 36.145 2.814 ;
      RECT 35.92 2.66 36.15 2.781 ;
      RECT 35.95 2.532 36.135 2.865 ;
      RECT 36.01 2.51 36.11 2.865 ;
      RECT 36.035 2.507 36.11 2.865 ;
      RECT 36.035 2.502 36.055 2.865 ;
      RECT 35.44 2.57 35.615 2.745 ;
      RECT 35.435 2.57 35.615 2.743 ;
      RECT 35.41 2.57 35.615 2.738 ;
      RECT 35.355 2.55 35.525 2.728 ;
      RECT 35.355 2.557 35.59 2.728 ;
      RECT 35.44 3.237 35.455 3.42 ;
      RECT 35.43 3.215 35.44 3.42 ;
      RECT 35.415 3.195 35.43 3.42 ;
      RECT 35.405 3.17 35.415 3.42 ;
      RECT 35.375 3.135 35.405 3.42 ;
      RECT 35.34 3.075 35.375 3.42 ;
      RECT 35.335 3.037 35.34 3.42 ;
      RECT 35.285 2.988 35.335 3.42 ;
      RECT 35.275 2.938 35.285 3.408 ;
      RECT 35.26 2.917 35.275 3.368 ;
      RECT 35.24 2.885 35.26 3.318 ;
      RECT 35.215 2.841 35.24 3.258 ;
      RECT 35.21 2.813 35.215 3.213 ;
      RECT 35.205 2.804 35.21 3.199 ;
      RECT 35.2 2.797 35.205 3.186 ;
      RECT 35.195 2.792 35.2 3.175 ;
      RECT 35.19 2.777 35.195 3.165 ;
      RECT 35.185 2.755 35.19 3.152 ;
      RECT 35.175 2.715 35.185 3.127 ;
      RECT 35.15 2.645 35.175 3.083 ;
      RECT 35.145 2.585 35.15 3.048 ;
      RECT 35.13 2.565 35.145 3.015 ;
      RECT 35.125 2.565 35.13 2.99 ;
      RECT 35.095 2.565 35.125 2.945 ;
      RECT 35.05 2.565 35.095 2.885 ;
      RECT 34.975 2.565 35.05 2.833 ;
      RECT 34.97 2.565 34.975 2.798 ;
      RECT 34.965 2.565 34.97 2.788 ;
      RECT 34.96 2.565 34.965 2.768 ;
      RECT 35.225 1.785 35.395 2.255 ;
      RECT 35.17 1.778 35.365 2.239 ;
      RECT 35.17 1.792 35.4 2.238 ;
      RECT 35.155 1.793 35.4 2.219 ;
      RECT 35.15 1.811 35.4 2.205 ;
      RECT 35.155 1.794 35.405 2.203 ;
      RECT 35.14 1.825 35.405 2.188 ;
      RECT 35.155 1.8 35.41 2.173 ;
      RECT 35.135 1.84 35.41 2.17 ;
      RECT 35.15 1.812 35.415 2.155 ;
      RECT 35.15 1.824 35.42 2.135 ;
      RECT 35.135 1.84 35.425 2.118 ;
      RECT 35.135 1.85 35.43 1.973 ;
      RECT 35.13 1.85 35.43 1.93 ;
      RECT 35.13 1.865 35.435 1.908 ;
      RECT 35.225 1.775 35.365 2.255 ;
      RECT 35.225 1.773 35.335 2.255 ;
      RECT 35.311 1.77 35.335 2.255 ;
      RECT 34.97 3.437 34.975 3.483 ;
      RECT 34.96 3.285 34.97 3.507 ;
      RECT 34.955 3.13 34.96 3.532 ;
      RECT 34.94 3.092 34.955 3.543 ;
      RECT 34.935 3.075 34.94 3.55 ;
      RECT 34.925 3.063 34.935 3.557 ;
      RECT 34.92 3.054 34.925 3.559 ;
      RECT 34.915 3.052 34.92 3.563 ;
      RECT 34.87 3.043 34.915 3.578 ;
      RECT 34.865 3.035 34.87 3.592 ;
      RECT 34.86 3.032 34.865 3.596 ;
      RECT 34.845 3.027 34.86 3.604 ;
      RECT 34.79 3.017 34.845 3.615 ;
      RECT 34.755 3.005 34.79 3.616 ;
      RECT 34.746 3 34.755 3.61 ;
      RECT 34.66 3 34.746 3.6 ;
      RECT 34.63 3 34.66 3.578 ;
      RECT 34.62 3 34.625 3.558 ;
      RECT 34.615 3 34.62 3.52 ;
      RECT 34.61 3 34.615 3.478 ;
      RECT 34.605 3 34.61 3.438 ;
      RECT 34.6 3 34.605 3.368 ;
      RECT 34.59 3 34.6 3.29 ;
      RECT 34.585 3 34.59 3.19 ;
      RECT 34.625 3 34.63 3.56 ;
      RECT 34.12 3.082 34.21 3.56 ;
      RECT 34.105 3.085 34.225 3.558 ;
      RECT 34.12 3.084 34.225 3.558 ;
      RECT 34.085 3.091 34.25 3.548 ;
      RECT 34.105 3.085 34.25 3.548 ;
      RECT 34.07 3.097 34.25 3.536 ;
      RECT 34.105 3.088 34.3 3.529 ;
      RECT 34.056 3.105 34.3 3.527 ;
      RECT 34.085 3.095 34.31 3.515 ;
      RECT 34.056 3.116 34.34 3.506 ;
      RECT 33.97 3.14 34.34 3.5 ;
      RECT 33.97 3.153 34.38 3.483 ;
      RECT 33.965 3.175 34.38 3.476 ;
      RECT 33.935 3.19 34.38 3.466 ;
      RECT 33.93 3.201 34.38 3.456 ;
      RECT 33.9 3.214 34.38 3.447 ;
      RECT 33.885 3.232 34.38 3.436 ;
      RECT 33.86 3.245 34.38 3.426 ;
      RECT 34.12 3.081 34.13 3.56 ;
      RECT 34.166 2.505 34.205 2.75 ;
      RECT 34.08 2.505 34.215 2.748 ;
      RECT 33.965 2.53 34.215 2.745 ;
      RECT 33.965 2.53 34.22 2.743 ;
      RECT 33.965 2.53 34.235 2.738 ;
      RECT 34.071 2.505 34.25 2.718 ;
      RECT 33.985 2.513 34.25 2.718 ;
      RECT 33.655 1.865 33.825 2.3 ;
      RECT 33.645 1.899 33.825 2.283 ;
      RECT 33.725 1.835 33.895 2.27 ;
      RECT 33.63 1.91 33.895 2.248 ;
      RECT 33.725 1.845 33.9 2.238 ;
      RECT 33.655 1.897 33.93 2.223 ;
      RECT 33.615 1.923 33.93 2.208 ;
      RECT 33.615 1.965 33.94 2.188 ;
      RECT 33.61 1.99 33.945 2.17 ;
      RECT 33.61 2 33.95 2.155 ;
      RECT 33.605 1.937 33.93 2.153 ;
      RECT 33.605 2.01 33.955 2.138 ;
      RECT 33.6 1.947 33.93 2.135 ;
      RECT 33.595 2.031 33.96 2.118 ;
      RECT 33.595 2.063 33.965 2.098 ;
      RECT 33.59 1.977 33.94 2.09 ;
      RECT 33.595 1.962 33.93 2.118 ;
      RECT 33.61 1.932 33.93 2.17 ;
      RECT 33.455 2.519 33.68 2.775 ;
      RECT 33.455 2.552 33.7 2.765 ;
      RECT 33.42 2.552 33.7 2.763 ;
      RECT 33.42 2.565 33.705 2.753 ;
      RECT 33.42 2.585 33.715 2.745 ;
      RECT 33.42 2.682 33.72 2.738 ;
      RECT 33.4 2.43 33.53 2.728 ;
      RECT 33.355 2.585 33.715 2.67 ;
      RECT 33.345 2.43 33.53 2.615 ;
      RECT 33.345 2.462 33.616 2.615 ;
      RECT 33.31 2.992 33.33 3.17 ;
      RECT 33.275 2.945 33.31 3.17 ;
      RECT 33.26 2.885 33.275 3.17 ;
      RECT 33.235 2.832 33.26 3.17 ;
      RECT 33.22 2.785 33.235 3.17 ;
      RECT 33.2 2.762 33.22 3.17 ;
      RECT 33.175 2.727 33.2 3.17 ;
      RECT 33.165 2.573 33.175 3.17 ;
      RECT 33.135 2.568 33.165 3.161 ;
      RECT 33.13 2.565 33.135 3.151 ;
      RECT 33.115 2.565 33.13 3.125 ;
      RECT 33.11 2.565 33.115 3.088 ;
      RECT 33.085 2.565 33.11 3.04 ;
      RECT 33.065 2.565 33.085 2.965 ;
      RECT 33.055 2.565 33.065 2.925 ;
      RECT 33.05 2.565 33.055 2.9 ;
      RECT 33.045 2.565 33.05 2.883 ;
      RECT 33.04 2.565 33.045 2.865 ;
      RECT 33.035 2.566 33.04 2.855 ;
      RECT 33.025 2.568 33.035 2.823 ;
      RECT 33.015 2.57 33.025 2.79 ;
      RECT 33.005 2.573 33.015 2.763 ;
      RECT 33.33 3 33.555 3.17 ;
      RECT 32.66 1.812 32.83 2.265 ;
      RECT 32.66 1.812 32.92 2.231 ;
      RECT 32.66 1.812 32.95 2.215 ;
      RECT 32.66 1.812 32.98 2.188 ;
      RECT 32.916 1.79 32.995 2.17 ;
      RECT 32.695 1.797 33 2.155 ;
      RECT 32.695 1.805 33.01 2.118 ;
      RECT 32.655 1.832 33.01 2.09 ;
      RECT 32.64 1.845 33.01 2.055 ;
      RECT 32.66 1.82 33.03 2.045 ;
      RECT 32.635 1.885 33.03 2.015 ;
      RECT 32.635 1.915 33.035 1.998 ;
      RECT 32.63 1.945 33.035 1.985 ;
      RECT 32.695 1.794 32.995 2.17 ;
      RECT 32.83 1.791 32.916 2.249 ;
      RECT 32.781 1.792 32.995 2.17 ;
      RECT 32.925 3.452 32.97 3.645 ;
      RECT 32.915 3.422 32.925 3.645 ;
      RECT 32.91 3.407 32.915 3.645 ;
      RECT 32.87 3.317 32.91 3.645 ;
      RECT 32.865 3.23 32.87 3.645 ;
      RECT 32.855 3.2 32.865 3.645 ;
      RECT 32.85 3.16 32.855 3.645 ;
      RECT 32.84 3.122 32.85 3.645 ;
      RECT 32.835 3.087 32.84 3.645 ;
      RECT 32.815 3.04 32.835 3.645 ;
      RECT 32.8 2.965 32.815 3.645 ;
      RECT 32.795 2.92 32.8 3.64 ;
      RECT 32.79 2.9 32.795 3.613 ;
      RECT 32.785 2.88 32.79 3.598 ;
      RECT 32.78 2.855 32.785 3.578 ;
      RECT 32.775 2.833 32.78 3.563 ;
      RECT 32.77 2.811 32.775 3.545 ;
      RECT 32.765 2.79 32.77 3.535 ;
      RECT 32.755 2.762 32.765 3.505 ;
      RECT 32.745 2.725 32.755 3.473 ;
      RECT 32.735 2.685 32.745 3.44 ;
      RECT 32.725 2.663 32.735 3.41 ;
      RECT 32.695 2.615 32.725 3.342 ;
      RECT 32.68 2.575 32.695 3.269 ;
      RECT 32.67 2.575 32.68 3.235 ;
      RECT 32.665 2.575 32.67 3.21 ;
      RECT 32.66 2.575 32.665 3.195 ;
      RECT 32.655 2.575 32.66 3.173 ;
      RECT 32.65 2.575 32.655 3.16 ;
      RECT 32.635 2.575 32.65 3.125 ;
      RECT 32.615 2.575 32.635 3.065 ;
      RECT 32.605 2.575 32.615 3.015 ;
      RECT 32.585 2.575 32.605 2.963 ;
      RECT 32.565 2.575 32.585 2.92 ;
      RECT 32.555 2.575 32.565 2.908 ;
      RECT 32.525 2.575 32.555 2.895 ;
      RECT 32.495 2.596 32.525 2.875 ;
      RECT 32.485 2.624 32.495 2.855 ;
      RECT 32.47 2.641 32.485 2.823 ;
      RECT 32.465 2.655 32.47 2.79 ;
      RECT 32.46 2.663 32.465 2.763 ;
      RECT 32.455 2.671 32.46 2.725 ;
      RECT 32.46 3.195 32.465 3.53 ;
      RECT 32.425 3.182 32.46 3.529 ;
      RECT 32.355 3.122 32.425 3.528 ;
      RECT 32.275 3.065 32.355 3.527 ;
      RECT 32.14 3.025 32.275 3.526 ;
      RECT 32.14 3.212 32.475 3.515 ;
      RECT 32.1 3.212 32.475 3.505 ;
      RECT 32.1 3.23 32.48 3.5 ;
      RECT 32.1 3.32 32.485 3.49 ;
      RECT 32.095 3.015 32.26 3.47 ;
      RECT 32.09 3.015 32.26 3.213 ;
      RECT 32.09 3.172 32.455 3.213 ;
      RECT 32.09 3.16 32.45 3.213 ;
      RECT 30.79 1.74 30.96 2.935 ;
      RECT 30.79 1.74 31.255 1.91 ;
      RECT 30.79 6.97 31.255 7.14 ;
      RECT 30.79 5.945 30.96 7.14 ;
      RECT 29.8 1.74 29.97 2.935 ;
      RECT 29.8 1.74 30.265 1.91 ;
      RECT 29.8 6.97 30.265 7.14 ;
      RECT 29.8 5.945 29.97 7.14 ;
      RECT 27.945 2.635 28.115 3.865 ;
      RECT 28 0.855 28.17 2.805 ;
      RECT 27.945 0.575 28.115 1.025 ;
      RECT 27.945 7.855 28.115 8.305 ;
      RECT 28 6.075 28.17 8.025 ;
      RECT 27.945 5.015 28.115 6.245 ;
      RECT 27.425 0.575 27.595 3.865 ;
      RECT 27.425 2.075 27.83 2.405 ;
      RECT 27.425 1.235 27.83 1.565 ;
      RECT 27.425 5.015 27.595 8.305 ;
      RECT 27.425 7.315 27.83 7.645 ;
      RECT 27.425 6.475 27.83 6.805 ;
      RECT 24.76 1.975 25.49 2.215 ;
      RECT 25.302 1.77 25.49 2.215 ;
      RECT 25.13 1.782 25.505 2.209 ;
      RECT 25.045 1.797 25.525 2.194 ;
      RECT 25.045 1.812 25.53 2.184 ;
      RECT 25 1.832 25.545 2.176 ;
      RECT 24.977 1.867 25.56 2.13 ;
      RECT 24.891 1.89 25.565 2.09 ;
      RECT 24.891 1.908 25.575 2.06 ;
      RECT 24.76 1.977 25.58 2.023 ;
      RECT 24.805 1.92 25.575 2.06 ;
      RECT 24.891 1.872 25.56 2.13 ;
      RECT 24.977 1.841 25.545 2.176 ;
      RECT 25 1.822 25.53 2.184 ;
      RECT 25.045 1.795 25.505 2.209 ;
      RECT 25.13 1.777 25.49 2.215 ;
      RECT 25.216 1.771 25.49 2.215 ;
      RECT 25.302 1.766 25.435 2.215 ;
      RECT 25.388 1.761 25.435 2.215 ;
      RECT 25.08 2.659 25.25 3.045 ;
      RECT 25.075 2.659 25.25 3.04 ;
      RECT 25.05 2.659 25.25 3.005 ;
      RECT 25.05 2.687 25.26 2.995 ;
      RECT 25.03 2.687 25.26 2.955 ;
      RECT 25.025 2.687 25.26 2.928 ;
      RECT 25.025 2.705 25.265 2.92 ;
      RECT 24.97 2.705 25.265 2.855 ;
      RECT 24.97 2.722 25.275 2.838 ;
      RECT 24.96 2.722 25.275 2.778 ;
      RECT 24.96 2.739 25.28 2.775 ;
      RECT 24.955 2.575 25.125 2.753 ;
      RECT 24.955 2.609 25.211 2.753 ;
      RECT 24.95 3.375 24.955 3.388 ;
      RECT 24.945 3.27 24.95 3.393 ;
      RECT 24.92 3.13 24.945 3.408 ;
      RECT 24.885 3.081 24.92 3.44 ;
      RECT 24.88 3.049 24.885 3.46 ;
      RECT 24.875 3.04 24.88 3.46 ;
      RECT 24.795 3.005 24.875 3.46 ;
      RECT 24.732 2.975 24.795 3.46 ;
      RECT 24.646 2.963 24.732 3.46 ;
      RECT 24.56 2.949 24.646 3.46 ;
      RECT 24.48 2.936 24.56 3.446 ;
      RECT 24.445 2.928 24.48 3.426 ;
      RECT 24.435 2.925 24.445 3.417 ;
      RECT 24.405 2.92 24.435 3.404 ;
      RECT 24.355 2.895 24.405 3.38 ;
      RECT 24.341 2.869 24.355 3.362 ;
      RECT 24.255 2.829 24.341 3.338 ;
      RECT 24.21 2.777 24.255 3.307 ;
      RECT 24.2 2.752 24.21 3.294 ;
      RECT 24.195 2.533 24.2 2.555 ;
      RECT 24.19 2.735 24.2 3.29 ;
      RECT 24.19 2.531 24.195 2.645 ;
      RECT 24.18 2.527 24.19 3.286 ;
      RECT 24.136 2.525 24.18 3.274 ;
      RECT 24.05 2.525 24.136 3.245 ;
      RECT 24.02 2.525 24.05 3.218 ;
      RECT 24.005 2.525 24.02 3.206 ;
      RECT 23.965 2.537 24.005 3.191 ;
      RECT 23.945 2.556 23.965 3.17 ;
      RECT 23.935 2.566 23.945 3.154 ;
      RECT 23.925 2.572 23.935 3.143 ;
      RECT 23.905 2.582 23.925 3.126 ;
      RECT 23.9 2.591 23.905 3.113 ;
      RECT 23.895 2.595 23.9 3.063 ;
      RECT 23.885 2.601 23.895 2.98 ;
      RECT 23.88 2.605 23.885 2.894 ;
      RECT 23.875 2.625 23.88 2.831 ;
      RECT 23.87 2.648 23.875 2.778 ;
      RECT 23.865 2.666 23.87 2.723 ;
      RECT 24.475 2.485 24.645 2.745 ;
      RECT 24.645 2.45 24.69 2.731 ;
      RECT 24.606 2.452 24.695 2.714 ;
      RECT 24.495 2.469 24.781 2.685 ;
      RECT 24.495 2.484 24.785 2.657 ;
      RECT 24.495 2.465 24.695 2.714 ;
      RECT 24.52 2.453 24.645 2.745 ;
      RECT 24.606 2.451 24.69 2.731 ;
      RECT 23.66 1.84 23.83 2.33 ;
      RECT 23.66 1.84 23.865 2.31 ;
      RECT 23.795 1.76 23.905 2.27 ;
      RECT 23.776 1.764 23.925 2.24 ;
      RECT 23.69 1.772 23.945 2.223 ;
      RECT 23.69 1.778 23.95 2.213 ;
      RECT 23.69 1.787 23.97 2.201 ;
      RECT 23.665 1.812 24 2.179 ;
      RECT 23.665 1.832 24.005 2.159 ;
      RECT 23.66 1.845 24.015 2.139 ;
      RECT 23.66 1.912 24.02 2.12 ;
      RECT 23.66 2.045 24.025 2.107 ;
      RECT 23.655 1.85 24.015 1.94 ;
      RECT 23.665 1.807 23.97 2.201 ;
      RECT 23.776 1.762 23.905 2.27 ;
      RECT 23.65 3.515 23.95 3.77 ;
      RECT 23.735 3.481 23.95 3.77 ;
      RECT 23.735 3.484 23.955 3.63 ;
      RECT 23.67 3.505 23.955 3.63 ;
      RECT 23.705 3.495 23.95 3.77 ;
      RECT 23.7 3.5 23.955 3.63 ;
      RECT 23.735 3.479 23.936 3.77 ;
      RECT 23.821 3.47 23.936 3.77 ;
      RECT 23.821 3.464 23.85 3.77 ;
      RECT 23.31 3.105 23.32 3.595 ;
      RECT 22.97 3.04 22.98 3.34 ;
      RECT 23.485 3.212 23.49 3.431 ;
      RECT 23.475 3.192 23.485 3.448 ;
      RECT 23.465 3.172 23.475 3.478 ;
      RECT 23.46 3.162 23.465 3.493 ;
      RECT 23.455 3.158 23.46 3.498 ;
      RECT 23.44 3.15 23.455 3.505 ;
      RECT 23.4 3.13 23.44 3.53 ;
      RECT 23.375 3.112 23.4 3.563 ;
      RECT 23.37 3.11 23.375 3.576 ;
      RECT 23.35 3.107 23.37 3.58 ;
      RECT 23.32 3.105 23.35 3.59 ;
      RECT 23.25 3.107 23.31 3.591 ;
      RECT 23.23 3.107 23.25 3.585 ;
      RECT 23.205 3.105 23.23 3.582 ;
      RECT 23.17 3.1 23.205 3.578 ;
      RECT 23.15 3.094 23.17 3.565 ;
      RECT 23.14 3.091 23.15 3.553 ;
      RECT 23.12 3.088 23.14 3.538 ;
      RECT 23.1 3.084 23.12 3.52 ;
      RECT 23.095 3.081 23.1 3.51 ;
      RECT 23.09 3.08 23.095 3.508 ;
      RECT 23.08 3.077 23.09 3.5 ;
      RECT 23.07 3.071 23.08 3.483 ;
      RECT 23.06 3.065 23.07 3.465 ;
      RECT 23.05 3.059 23.06 3.453 ;
      RECT 23.04 3.053 23.05 3.433 ;
      RECT 23.035 3.049 23.04 3.418 ;
      RECT 23.03 3.047 23.035 3.41 ;
      RECT 23.025 3.045 23.03 3.403 ;
      RECT 23.02 3.043 23.025 3.393 ;
      RECT 23.015 3.041 23.02 3.387 ;
      RECT 23.005 3.04 23.015 3.377 ;
      RECT 22.995 3.04 23.005 3.368 ;
      RECT 22.98 3.04 22.995 3.353 ;
      RECT 22.94 3.04 22.97 3.337 ;
      RECT 22.92 3.042 22.94 3.332 ;
      RECT 22.915 3.047 22.92 3.33 ;
      RECT 22.885 3.055 22.915 3.328 ;
      RECT 22.855 3.07 22.885 3.327 ;
      RECT 22.81 3.092 22.855 3.332 ;
      RECT 22.805 3.107 22.81 3.336 ;
      RECT 22.79 3.112 22.805 3.338 ;
      RECT 22.785 3.116 22.79 3.34 ;
      RECT 22.725 3.139 22.785 3.349 ;
      RECT 22.705 3.165 22.725 3.362 ;
      RECT 22.695 3.172 22.705 3.366 ;
      RECT 22.68 3.179 22.695 3.369 ;
      RECT 22.66 3.189 22.68 3.372 ;
      RECT 22.655 3.197 22.66 3.375 ;
      RECT 22.61 3.202 22.655 3.382 ;
      RECT 22.6 3.205 22.61 3.389 ;
      RECT 22.59 3.205 22.6 3.393 ;
      RECT 22.555 3.207 22.59 3.405 ;
      RECT 22.535 3.21 22.555 3.418 ;
      RECT 22.495 3.213 22.535 3.429 ;
      RECT 22.48 3.215 22.495 3.442 ;
      RECT 22.47 3.215 22.48 3.447 ;
      RECT 22.445 3.216 22.47 3.455 ;
      RECT 22.435 3.218 22.445 3.46 ;
      RECT 22.43 3.219 22.435 3.463 ;
      RECT 22.405 3.217 22.43 3.466 ;
      RECT 22.39 3.215 22.405 3.467 ;
      RECT 22.37 3.212 22.39 3.469 ;
      RECT 22.35 3.207 22.37 3.469 ;
      RECT 22.29 3.202 22.35 3.466 ;
      RECT 22.255 3.177 22.29 3.462 ;
      RECT 22.245 3.154 22.255 3.46 ;
      RECT 22.215 3.131 22.245 3.46 ;
      RECT 22.205 3.11 22.215 3.46 ;
      RECT 22.18 3.092 22.205 3.458 ;
      RECT 22.165 3.07 22.18 3.455 ;
      RECT 22.15 3.052 22.165 3.453 ;
      RECT 22.13 3.042 22.15 3.451 ;
      RECT 22.115 3.037 22.13 3.45 ;
      RECT 22.1 3.035 22.115 3.449 ;
      RECT 22.07 3.036 22.1 3.447 ;
      RECT 22.05 3.039 22.07 3.445 ;
      RECT 21.993 3.043 22.05 3.445 ;
      RECT 21.907 3.052 21.993 3.445 ;
      RECT 21.821 3.063 21.907 3.445 ;
      RECT 21.735 3.074 21.821 3.445 ;
      RECT 21.715 3.081 21.735 3.453 ;
      RECT 21.705 3.084 21.715 3.46 ;
      RECT 21.64 3.089 21.705 3.478 ;
      RECT 21.61 3.096 21.64 3.503 ;
      RECT 21.6 3.099 21.61 3.51 ;
      RECT 21.555 3.103 21.6 3.515 ;
      RECT 21.525 3.108 21.555 3.52 ;
      RECT 21.524 3.11 21.525 3.52 ;
      RECT 21.438 3.116 21.524 3.52 ;
      RECT 21.352 3.127 21.438 3.52 ;
      RECT 21.266 3.139 21.352 3.52 ;
      RECT 21.18 3.15 21.266 3.52 ;
      RECT 21.165 3.157 21.18 3.515 ;
      RECT 21.16 3.159 21.165 3.509 ;
      RECT 21.14 3.17 21.16 3.504 ;
      RECT 21.13 3.188 21.14 3.498 ;
      RECT 21.125 3.2 21.13 3.298 ;
      RECT 23.42 1.953 23.44 2.04 ;
      RECT 23.415 1.888 23.42 2.072 ;
      RECT 23.405 1.855 23.415 2.077 ;
      RECT 23.4 1.835 23.405 2.083 ;
      RECT 23.37 1.835 23.4 2.1 ;
      RECT 23.321 1.835 23.37 2.136 ;
      RECT 23.235 1.835 23.321 2.194 ;
      RECT 23.206 1.845 23.235 2.243 ;
      RECT 23.12 1.887 23.206 2.296 ;
      RECT 23.1 1.925 23.12 2.343 ;
      RECT 23.075 1.942 23.1 2.363 ;
      RECT 23.065 1.956 23.075 2.383 ;
      RECT 23.06 1.962 23.065 2.393 ;
      RECT 23.055 1.966 23.06 2.4 ;
      RECT 23.005 1.986 23.055 2.405 ;
      RECT 22.94 2.03 23.005 2.405 ;
      RECT 22.915 2.08 22.94 2.405 ;
      RECT 22.905 2.11 22.915 2.405 ;
      RECT 22.9 2.137 22.905 2.405 ;
      RECT 22.895 2.155 22.9 2.405 ;
      RECT 22.885 2.197 22.895 2.405 ;
      RECT 23.235 2.755 23.405 2.93 ;
      RECT 23.175 2.583 23.235 2.918 ;
      RECT 23.165 2.576 23.175 2.901 ;
      RECT 23.12 2.755 23.405 2.881 ;
      RECT 23.101 2.755 23.405 2.859 ;
      RECT 23.015 2.755 23.405 2.824 ;
      RECT 22.995 2.575 23.165 2.78 ;
      RECT 22.995 2.722 23.4 2.78 ;
      RECT 22.995 2.67 23.375 2.78 ;
      RECT 22.995 2.625 23.34 2.78 ;
      RECT 22.995 2.607 23.305 2.78 ;
      RECT 22.995 2.597 23.3 2.78 ;
      RECT 22.715 3.555 22.905 3.78 ;
      RECT 22.705 3.556 22.91 3.775 ;
      RECT 22.705 3.558 22.92 3.755 ;
      RECT 22.705 3.562 22.925 3.74 ;
      RECT 22.705 3.549 22.875 3.775 ;
      RECT 22.705 3.552 22.9 3.775 ;
      RECT 22.715 3.548 22.875 3.78 ;
      RECT 22.801 3.546 22.875 3.78 ;
      RECT 22.425 2.797 22.595 3.035 ;
      RECT 22.425 2.797 22.681 2.949 ;
      RECT 22.425 2.797 22.685 2.859 ;
      RECT 22.475 2.57 22.695 2.838 ;
      RECT 22.47 2.587 22.7 2.811 ;
      RECT 22.435 2.745 22.7 2.811 ;
      RECT 22.455 2.595 22.595 3.035 ;
      RECT 22.445 2.677 22.705 2.794 ;
      RECT 22.44 2.725 22.705 2.794 ;
      RECT 22.445 2.635 22.7 2.811 ;
      RECT 22.47 2.572 22.695 2.838 ;
      RECT 22.035 2.547 22.205 2.745 ;
      RECT 22.035 2.547 22.25 2.72 ;
      RECT 22.105 2.49 22.275 2.678 ;
      RECT 22.08 2.505 22.275 2.678 ;
      RECT 21.695 2.551 21.725 2.745 ;
      RECT 21.69 2.523 21.695 2.745 ;
      RECT 21.66 2.497 21.69 2.747 ;
      RECT 21.635 2.455 21.66 2.75 ;
      RECT 21.625 2.427 21.635 2.752 ;
      RECT 21.59 2.407 21.625 2.754 ;
      RECT 21.525 2.392 21.59 2.76 ;
      RECT 21.475 2.39 21.525 2.766 ;
      RECT 21.452 2.392 21.475 2.771 ;
      RECT 21.366 2.403 21.452 2.777 ;
      RECT 21.28 2.421 21.366 2.787 ;
      RECT 21.265 2.432 21.28 2.793 ;
      RECT 21.195 2.455 21.265 2.799 ;
      RECT 21.14 2.487 21.195 2.807 ;
      RECT 21.1 2.51 21.14 2.813 ;
      RECT 21.086 2.523 21.1 2.816 ;
      RECT 21 2.545 21.086 2.822 ;
      RECT 20.985 2.57 21 2.828 ;
      RECT 20.945 2.585 20.985 2.832 ;
      RECT 20.895 2.6 20.945 2.837 ;
      RECT 20.87 2.607 20.895 2.841 ;
      RECT 20.81 2.602 20.87 2.845 ;
      RECT 20.795 2.593 20.81 2.849 ;
      RECT 20.725 2.583 20.795 2.845 ;
      RECT 20.7 2.575 20.72 2.835 ;
      RECT 20.641 2.575 20.7 2.813 ;
      RECT 20.555 2.575 20.641 2.77 ;
      RECT 20.72 2.575 20.725 2.84 ;
      RECT 21.415 1.806 21.585 2.14 ;
      RECT 21.385 1.806 21.585 2.135 ;
      RECT 21.325 1.773 21.385 2.123 ;
      RECT 21.325 1.829 21.595 2.118 ;
      RECT 21.3 1.829 21.595 2.112 ;
      RECT 21.295 1.77 21.325 2.109 ;
      RECT 21.28 1.776 21.415 2.107 ;
      RECT 21.275 1.784 21.5 2.095 ;
      RECT 21.275 1.836 21.61 2.048 ;
      RECT 21.26 1.792 21.5 2.043 ;
      RECT 21.26 1.862 21.62 1.984 ;
      RECT 21.23 1.812 21.585 1.945 ;
      RECT 21.23 1.902 21.63 1.941 ;
      RECT 21.28 1.781 21.5 2.107 ;
      RECT 20.62 2.111 20.675 2.375 ;
      RECT 20.62 2.111 20.74 2.374 ;
      RECT 20.62 2.111 20.765 2.373 ;
      RECT 20.62 2.111 20.83 2.372 ;
      RECT 20.765 2.077 20.845 2.371 ;
      RECT 20.58 2.121 20.99 2.37 ;
      RECT 20.62 2.118 20.99 2.37 ;
      RECT 20.58 2.126 20.995 2.363 ;
      RECT 20.565 2.128 20.995 2.362 ;
      RECT 20.565 2.135 21 2.358 ;
      RECT 20.545 2.134 20.995 2.354 ;
      RECT 20.545 2.142 21.005 2.353 ;
      RECT 20.54 2.139 21 2.349 ;
      RECT 20.54 2.152 21.015 2.348 ;
      RECT 20.525 2.142 21.005 2.347 ;
      RECT 20.49 2.155 21.015 2.34 ;
      RECT 20.675 2.11 20.985 2.37 ;
      RECT 20.675 2.095 20.935 2.37 ;
      RECT 20.74 2.082 20.87 2.37 ;
      RECT 20.285 3.171 20.3 3.564 ;
      RECT 20.25 3.176 20.3 3.563 ;
      RECT 20.285 3.175 20.345 3.562 ;
      RECT 20.23 3.186 20.345 3.561 ;
      RECT 20.245 3.182 20.345 3.561 ;
      RECT 20.21 3.192 20.42 3.558 ;
      RECT 20.21 3.211 20.465 3.556 ;
      RECT 20.21 3.218 20.47 3.553 ;
      RECT 20.195 3.195 20.42 3.55 ;
      RECT 20.175 3.2 20.42 3.543 ;
      RECT 20.17 3.204 20.42 3.539 ;
      RECT 20.17 3.221 20.48 3.538 ;
      RECT 20.15 3.215 20.465 3.534 ;
      RECT 20.15 3.224 20.485 3.528 ;
      RECT 20.145 3.23 20.485 3.3 ;
      RECT 20.21 3.19 20.345 3.558 ;
      RECT 20.085 2.553 20.285 2.865 ;
      RECT 20.16 2.531 20.285 2.865 ;
      RECT 20.1 2.55 20.29 2.85 ;
      RECT 20.07 2.561 20.29 2.848 ;
      RECT 20.085 2.556 20.295 2.814 ;
      RECT 20.07 2.66 20.3 2.781 ;
      RECT 20.1 2.532 20.285 2.865 ;
      RECT 20.16 2.51 20.26 2.865 ;
      RECT 20.185 2.507 20.26 2.865 ;
      RECT 20.185 2.502 20.205 2.865 ;
      RECT 19.59 2.57 19.765 2.745 ;
      RECT 19.585 2.57 19.765 2.743 ;
      RECT 19.56 2.57 19.765 2.738 ;
      RECT 19.505 2.55 19.675 2.728 ;
      RECT 19.505 2.557 19.74 2.728 ;
      RECT 19.59 3.237 19.605 3.42 ;
      RECT 19.58 3.215 19.59 3.42 ;
      RECT 19.565 3.195 19.58 3.42 ;
      RECT 19.555 3.17 19.565 3.42 ;
      RECT 19.525 3.135 19.555 3.42 ;
      RECT 19.49 3.075 19.525 3.42 ;
      RECT 19.485 3.037 19.49 3.42 ;
      RECT 19.435 2.988 19.485 3.42 ;
      RECT 19.425 2.938 19.435 3.408 ;
      RECT 19.41 2.917 19.425 3.368 ;
      RECT 19.39 2.885 19.41 3.318 ;
      RECT 19.365 2.841 19.39 3.258 ;
      RECT 19.36 2.813 19.365 3.213 ;
      RECT 19.355 2.804 19.36 3.199 ;
      RECT 19.35 2.797 19.355 3.186 ;
      RECT 19.345 2.792 19.35 3.175 ;
      RECT 19.34 2.777 19.345 3.165 ;
      RECT 19.335 2.755 19.34 3.152 ;
      RECT 19.325 2.715 19.335 3.127 ;
      RECT 19.3 2.645 19.325 3.083 ;
      RECT 19.295 2.585 19.3 3.048 ;
      RECT 19.28 2.565 19.295 3.015 ;
      RECT 19.275 2.565 19.28 2.99 ;
      RECT 19.245 2.565 19.275 2.945 ;
      RECT 19.2 2.565 19.245 2.885 ;
      RECT 19.125 2.565 19.2 2.833 ;
      RECT 19.12 2.565 19.125 2.798 ;
      RECT 19.115 2.565 19.12 2.788 ;
      RECT 19.11 2.565 19.115 2.768 ;
      RECT 19.375 1.785 19.545 2.255 ;
      RECT 19.32 1.778 19.515 2.239 ;
      RECT 19.32 1.792 19.55 2.238 ;
      RECT 19.305 1.793 19.55 2.219 ;
      RECT 19.3 1.811 19.55 2.205 ;
      RECT 19.305 1.794 19.555 2.203 ;
      RECT 19.29 1.825 19.555 2.188 ;
      RECT 19.305 1.8 19.56 2.173 ;
      RECT 19.285 1.84 19.56 2.17 ;
      RECT 19.3 1.812 19.565 2.155 ;
      RECT 19.3 1.824 19.57 2.135 ;
      RECT 19.285 1.84 19.575 2.118 ;
      RECT 19.285 1.85 19.58 1.973 ;
      RECT 19.28 1.85 19.58 1.93 ;
      RECT 19.28 1.865 19.585 1.908 ;
      RECT 19.375 1.775 19.515 2.255 ;
      RECT 19.375 1.773 19.485 2.255 ;
      RECT 19.461 1.77 19.485 2.255 ;
      RECT 19.12 3.437 19.125 3.483 ;
      RECT 19.11 3.285 19.12 3.507 ;
      RECT 19.105 3.13 19.11 3.532 ;
      RECT 19.09 3.092 19.105 3.543 ;
      RECT 19.085 3.075 19.09 3.55 ;
      RECT 19.075 3.063 19.085 3.557 ;
      RECT 19.07 3.054 19.075 3.559 ;
      RECT 19.065 3.052 19.07 3.563 ;
      RECT 19.02 3.043 19.065 3.578 ;
      RECT 19.015 3.035 19.02 3.592 ;
      RECT 19.01 3.032 19.015 3.596 ;
      RECT 18.995 3.027 19.01 3.604 ;
      RECT 18.94 3.017 18.995 3.615 ;
      RECT 18.905 3.005 18.94 3.616 ;
      RECT 18.896 3 18.905 3.61 ;
      RECT 18.81 3 18.896 3.6 ;
      RECT 18.78 3 18.81 3.578 ;
      RECT 18.77 3 18.775 3.558 ;
      RECT 18.765 3 18.77 3.52 ;
      RECT 18.76 3 18.765 3.478 ;
      RECT 18.755 3 18.76 3.438 ;
      RECT 18.75 3 18.755 3.368 ;
      RECT 18.74 3 18.75 3.29 ;
      RECT 18.735 3 18.74 3.19 ;
      RECT 18.775 3 18.78 3.56 ;
      RECT 18.27 3.082 18.36 3.56 ;
      RECT 18.255 3.085 18.375 3.558 ;
      RECT 18.27 3.084 18.375 3.558 ;
      RECT 18.235 3.091 18.4 3.548 ;
      RECT 18.255 3.085 18.4 3.548 ;
      RECT 18.22 3.097 18.4 3.536 ;
      RECT 18.255 3.088 18.45 3.529 ;
      RECT 18.206 3.105 18.45 3.527 ;
      RECT 18.235 3.095 18.46 3.515 ;
      RECT 18.206 3.116 18.49 3.506 ;
      RECT 18.12 3.14 18.49 3.5 ;
      RECT 18.12 3.153 18.53 3.483 ;
      RECT 18.115 3.175 18.53 3.476 ;
      RECT 18.085 3.19 18.53 3.466 ;
      RECT 18.08 3.201 18.53 3.456 ;
      RECT 18.05 3.214 18.53 3.447 ;
      RECT 18.035 3.232 18.53 3.436 ;
      RECT 18.01 3.245 18.53 3.426 ;
      RECT 18.27 3.081 18.28 3.56 ;
      RECT 18.316 2.505 18.355 2.75 ;
      RECT 18.23 2.505 18.365 2.748 ;
      RECT 18.115 2.53 18.365 2.745 ;
      RECT 18.115 2.53 18.37 2.743 ;
      RECT 18.115 2.53 18.385 2.738 ;
      RECT 18.221 2.505 18.4 2.718 ;
      RECT 18.135 2.513 18.4 2.718 ;
      RECT 17.805 1.865 17.975 2.3 ;
      RECT 17.795 1.899 17.975 2.283 ;
      RECT 17.875 1.835 18.045 2.27 ;
      RECT 17.78 1.91 18.045 2.248 ;
      RECT 17.875 1.845 18.05 2.238 ;
      RECT 17.805 1.897 18.08 2.223 ;
      RECT 17.765 1.923 18.08 2.208 ;
      RECT 17.765 1.965 18.09 2.188 ;
      RECT 17.76 1.99 18.095 2.17 ;
      RECT 17.76 2 18.1 2.155 ;
      RECT 17.755 1.937 18.08 2.153 ;
      RECT 17.755 2.01 18.105 2.138 ;
      RECT 17.75 1.947 18.08 2.135 ;
      RECT 17.745 2.031 18.11 2.118 ;
      RECT 17.745 2.063 18.115 2.098 ;
      RECT 17.74 1.977 18.09 2.09 ;
      RECT 17.745 1.962 18.08 2.118 ;
      RECT 17.76 1.932 18.08 2.17 ;
      RECT 17.605 2.519 17.83 2.775 ;
      RECT 17.605 2.552 17.85 2.765 ;
      RECT 17.57 2.552 17.85 2.763 ;
      RECT 17.57 2.565 17.855 2.753 ;
      RECT 17.57 2.585 17.865 2.745 ;
      RECT 17.57 2.682 17.87 2.738 ;
      RECT 17.55 2.43 17.68 2.728 ;
      RECT 17.505 2.585 17.865 2.67 ;
      RECT 17.495 2.43 17.68 2.615 ;
      RECT 17.495 2.462 17.766 2.615 ;
      RECT 17.46 2.992 17.48 3.17 ;
      RECT 17.425 2.945 17.46 3.17 ;
      RECT 17.41 2.885 17.425 3.17 ;
      RECT 17.385 2.832 17.41 3.17 ;
      RECT 17.37 2.785 17.385 3.17 ;
      RECT 17.35 2.762 17.37 3.17 ;
      RECT 17.325 2.727 17.35 3.17 ;
      RECT 17.315 2.573 17.325 3.17 ;
      RECT 17.285 2.568 17.315 3.161 ;
      RECT 17.28 2.565 17.285 3.151 ;
      RECT 17.265 2.565 17.28 3.125 ;
      RECT 17.26 2.565 17.265 3.088 ;
      RECT 17.235 2.565 17.26 3.04 ;
      RECT 17.215 2.565 17.235 2.965 ;
      RECT 17.205 2.565 17.215 2.925 ;
      RECT 17.2 2.565 17.205 2.9 ;
      RECT 17.195 2.565 17.2 2.883 ;
      RECT 17.19 2.565 17.195 2.865 ;
      RECT 17.185 2.566 17.19 2.855 ;
      RECT 17.175 2.568 17.185 2.823 ;
      RECT 17.165 2.57 17.175 2.79 ;
      RECT 17.155 2.573 17.165 2.763 ;
      RECT 17.48 3 17.705 3.17 ;
      RECT 16.81 1.812 16.98 2.265 ;
      RECT 16.81 1.812 17.07 2.231 ;
      RECT 16.81 1.812 17.1 2.215 ;
      RECT 16.81 1.812 17.13 2.188 ;
      RECT 17.066 1.79 17.145 2.17 ;
      RECT 16.845 1.797 17.15 2.155 ;
      RECT 16.845 1.805 17.16 2.118 ;
      RECT 16.805 1.832 17.16 2.09 ;
      RECT 16.79 1.845 17.16 2.055 ;
      RECT 16.81 1.82 17.18 2.045 ;
      RECT 16.785 1.885 17.18 2.015 ;
      RECT 16.785 1.915 17.185 1.998 ;
      RECT 16.78 1.945 17.185 1.985 ;
      RECT 16.845 1.794 17.145 2.17 ;
      RECT 16.98 1.791 17.066 2.249 ;
      RECT 16.931 1.792 17.145 2.17 ;
      RECT 17.075 3.452 17.12 3.645 ;
      RECT 17.065 3.422 17.075 3.645 ;
      RECT 17.06 3.407 17.065 3.645 ;
      RECT 17.02 3.317 17.06 3.645 ;
      RECT 17.015 3.23 17.02 3.645 ;
      RECT 17.005 3.2 17.015 3.645 ;
      RECT 17 3.16 17.005 3.645 ;
      RECT 16.99 3.122 17 3.645 ;
      RECT 16.985 3.087 16.99 3.645 ;
      RECT 16.965 3.04 16.985 3.645 ;
      RECT 16.95 2.965 16.965 3.645 ;
      RECT 16.945 2.92 16.95 3.64 ;
      RECT 16.94 2.9 16.945 3.613 ;
      RECT 16.935 2.88 16.94 3.598 ;
      RECT 16.93 2.855 16.935 3.578 ;
      RECT 16.925 2.833 16.93 3.563 ;
      RECT 16.92 2.811 16.925 3.545 ;
      RECT 16.915 2.79 16.92 3.535 ;
      RECT 16.905 2.762 16.915 3.505 ;
      RECT 16.895 2.725 16.905 3.473 ;
      RECT 16.885 2.685 16.895 3.44 ;
      RECT 16.875 2.663 16.885 3.41 ;
      RECT 16.845 2.615 16.875 3.342 ;
      RECT 16.83 2.575 16.845 3.269 ;
      RECT 16.82 2.575 16.83 3.235 ;
      RECT 16.815 2.575 16.82 3.21 ;
      RECT 16.81 2.575 16.815 3.195 ;
      RECT 16.805 2.575 16.81 3.173 ;
      RECT 16.8 2.575 16.805 3.16 ;
      RECT 16.785 2.575 16.8 3.125 ;
      RECT 16.765 2.575 16.785 3.065 ;
      RECT 16.755 2.575 16.765 3.015 ;
      RECT 16.735 2.575 16.755 2.963 ;
      RECT 16.715 2.575 16.735 2.92 ;
      RECT 16.705 2.575 16.715 2.908 ;
      RECT 16.675 2.575 16.705 2.895 ;
      RECT 16.645 2.596 16.675 2.875 ;
      RECT 16.635 2.624 16.645 2.855 ;
      RECT 16.62 2.641 16.635 2.823 ;
      RECT 16.615 2.655 16.62 2.79 ;
      RECT 16.61 2.663 16.615 2.763 ;
      RECT 16.605 2.671 16.61 2.725 ;
      RECT 16.61 3.195 16.615 3.53 ;
      RECT 16.575 3.182 16.61 3.529 ;
      RECT 16.505 3.122 16.575 3.528 ;
      RECT 16.425 3.065 16.505 3.527 ;
      RECT 16.29 3.025 16.425 3.526 ;
      RECT 16.29 3.212 16.625 3.515 ;
      RECT 16.25 3.212 16.625 3.505 ;
      RECT 16.25 3.23 16.63 3.5 ;
      RECT 16.25 3.32 16.635 3.49 ;
      RECT 16.245 3.015 16.41 3.47 ;
      RECT 16.24 3.015 16.41 3.213 ;
      RECT 16.24 3.172 16.605 3.213 ;
      RECT 16.24 3.16 16.6 3.213 ;
      RECT 14.94 1.74 15.11 2.935 ;
      RECT 14.94 1.74 15.405 1.91 ;
      RECT 14.94 6.97 15.405 7.14 ;
      RECT 14.94 5.945 15.11 7.14 ;
      RECT 13.95 1.74 14.12 2.935 ;
      RECT 13.95 1.74 14.415 1.91 ;
      RECT 13.95 6.97 14.415 7.14 ;
      RECT 13.95 5.945 14.12 7.14 ;
      RECT 12.095 2.635 12.265 3.865 ;
      RECT 12.15 0.855 12.32 2.805 ;
      RECT 12.095 0.575 12.265 1.025 ;
      RECT 12.095 7.855 12.265 8.305 ;
      RECT 12.15 6.075 12.32 8.025 ;
      RECT 12.095 5.015 12.265 6.245 ;
      RECT 11.575 0.575 11.745 3.865 ;
      RECT 11.575 2.075 11.98 2.405 ;
      RECT 11.575 1.235 11.98 1.565 ;
      RECT 11.575 5.015 11.745 8.305 ;
      RECT 11.575 7.315 11.98 7.645 ;
      RECT 11.575 6.475 11.98 6.805 ;
      RECT 8.91 1.975 9.64 2.215 ;
      RECT 9.452 1.77 9.64 2.215 ;
      RECT 9.28 1.782 9.655 2.209 ;
      RECT 9.195 1.797 9.675 2.194 ;
      RECT 9.195 1.812 9.68 2.184 ;
      RECT 9.15 1.832 9.695 2.176 ;
      RECT 9.127 1.867 9.71 2.13 ;
      RECT 9.041 1.89 9.715 2.09 ;
      RECT 9.041 1.908 9.725 2.06 ;
      RECT 8.91 1.977 9.73 2.023 ;
      RECT 8.955 1.92 9.725 2.06 ;
      RECT 9.041 1.872 9.71 2.13 ;
      RECT 9.127 1.841 9.695 2.176 ;
      RECT 9.15 1.822 9.68 2.184 ;
      RECT 9.195 1.795 9.655 2.209 ;
      RECT 9.28 1.777 9.64 2.215 ;
      RECT 9.366 1.771 9.64 2.215 ;
      RECT 9.452 1.766 9.585 2.215 ;
      RECT 9.538 1.761 9.585 2.215 ;
      RECT 9.23 2.659 9.4 3.045 ;
      RECT 9.225 2.659 9.4 3.04 ;
      RECT 9.2 2.659 9.4 3.005 ;
      RECT 9.2 2.687 9.41 2.995 ;
      RECT 9.18 2.687 9.41 2.955 ;
      RECT 9.175 2.687 9.41 2.928 ;
      RECT 9.175 2.705 9.415 2.92 ;
      RECT 9.12 2.705 9.415 2.855 ;
      RECT 9.12 2.722 9.425 2.838 ;
      RECT 9.11 2.722 9.425 2.778 ;
      RECT 9.11 2.739 9.43 2.775 ;
      RECT 9.105 2.575 9.275 2.753 ;
      RECT 9.105 2.609 9.361 2.753 ;
      RECT 9.1 3.375 9.105 3.388 ;
      RECT 9.095 3.27 9.1 3.393 ;
      RECT 9.07 3.13 9.095 3.408 ;
      RECT 9.035 3.081 9.07 3.44 ;
      RECT 9.03 3.049 9.035 3.46 ;
      RECT 9.025 3.04 9.03 3.46 ;
      RECT 8.945 3.005 9.025 3.46 ;
      RECT 8.882 2.975 8.945 3.46 ;
      RECT 8.796 2.963 8.882 3.46 ;
      RECT 8.71 2.949 8.796 3.46 ;
      RECT 8.63 2.936 8.71 3.446 ;
      RECT 8.595 2.928 8.63 3.426 ;
      RECT 8.585 2.925 8.595 3.417 ;
      RECT 8.555 2.92 8.585 3.404 ;
      RECT 8.505 2.895 8.555 3.38 ;
      RECT 8.491 2.869 8.505 3.362 ;
      RECT 8.405 2.829 8.491 3.338 ;
      RECT 8.36 2.777 8.405 3.307 ;
      RECT 8.35 2.752 8.36 3.294 ;
      RECT 8.345 2.533 8.35 2.555 ;
      RECT 8.34 2.735 8.35 3.29 ;
      RECT 8.34 2.531 8.345 2.645 ;
      RECT 8.33 2.527 8.34 3.286 ;
      RECT 8.286 2.525 8.33 3.274 ;
      RECT 8.2 2.525 8.286 3.245 ;
      RECT 8.17 2.525 8.2 3.218 ;
      RECT 8.155 2.525 8.17 3.206 ;
      RECT 8.115 2.537 8.155 3.191 ;
      RECT 8.095 2.556 8.115 3.17 ;
      RECT 8.085 2.566 8.095 3.154 ;
      RECT 8.075 2.572 8.085 3.143 ;
      RECT 8.055 2.582 8.075 3.126 ;
      RECT 8.05 2.591 8.055 3.113 ;
      RECT 8.045 2.595 8.05 3.063 ;
      RECT 8.035 2.601 8.045 2.98 ;
      RECT 8.03 2.605 8.035 2.894 ;
      RECT 8.025 2.625 8.03 2.831 ;
      RECT 8.02 2.648 8.025 2.778 ;
      RECT 8.015 2.666 8.02 2.723 ;
      RECT 8.625 2.485 8.795 2.745 ;
      RECT 8.795 2.45 8.84 2.731 ;
      RECT 8.756 2.452 8.845 2.714 ;
      RECT 8.645 2.469 8.931 2.685 ;
      RECT 8.645 2.484 8.935 2.657 ;
      RECT 8.645 2.465 8.845 2.714 ;
      RECT 8.67 2.453 8.795 2.745 ;
      RECT 8.756 2.451 8.84 2.731 ;
      RECT 7.81 1.84 7.98 2.33 ;
      RECT 7.81 1.84 8.015 2.31 ;
      RECT 7.945 1.76 8.055 2.27 ;
      RECT 7.926 1.764 8.075 2.24 ;
      RECT 7.84 1.772 8.095 2.223 ;
      RECT 7.84 1.778 8.1 2.213 ;
      RECT 7.84 1.787 8.12 2.201 ;
      RECT 7.815 1.812 8.15 2.179 ;
      RECT 7.815 1.832 8.155 2.159 ;
      RECT 7.81 1.845 8.165 2.139 ;
      RECT 7.81 1.912 8.17 2.12 ;
      RECT 7.81 2.045 8.175 2.107 ;
      RECT 7.805 1.85 8.165 1.94 ;
      RECT 7.815 1.807 8.12 2.201 ;
      RECT 7.926 1.762 8.055 2.27 ;
      RECT 7.8 3.515 8.1 3.77 ;
      RECT 7.885 3.481 8.1 3.77 ;
      RECT 7.885 3.484 8.105 3.63 ;
      RECT 7.82 3.505 8.105 3.63 ;
      RECT 7.855 3.495 8.1 3.77 ;
      RECT 7.85 3.5 8.105 3.63 ;
      RECT 7.885 3.479 8.086 3.77 ;
      RECT 7.971 3.47 8.086 3.77 ;
      RECT 7.971 3.464 8 3.77 ;
      RECT 7.46 3.105 7.47 3.595 ;
      RECT 7.12 3.04 7.13 3.34 ;
      RECT 7.635 3.212 7.64 3.431 ;
      RECT 7.625 3.192 7.635 3.448 ;
      RECT 7.615 3.172 7.625 3.478 ;
      RECT 7.61 3.162 7.615 3.493 ;
      RECT 7.605 3.158 7.61 3.498 ;
      RECT 7.59 3.15 7.605 3.505 ;
      RECT 7.55 3.13 7.59 3.53 ;
      RECT 7.525 3.112 7.55 3.563 ;
      RECT 7.52 3.11 7.525 3.576 ;
      RECT 7.5 3.107 7.52 3.58 ;
      RECT 7.47 3.105 7.5 3.59 ;
      RECT 7.4 3.107 7.46 3.591 ;
      RECT 7.38 3.107 7.4 3.585 ;
      RECT 7.355 3.105 7.38 3.582 ;
      RECT 7.32 3.1 7.355 3.578 ;
      RECT 7.3 3.094 7.32 3.565 ;
      RECT 7.29 3.091 7.3 3.553 ;
      RECT 7.27 3.088 7.29 3.538 ;
      RECT 7.25 3.084 7.27 3.52 ;
      RECT 7.245 3.081 7.25 3.51 ;
      RECT 7.24 3.08 7.245 3.508 ;
      RECT 7.23 3.077 7.24 3.5 ;
      RECT 7.22 3.071 7.23 3.483 ;
      RECT 7.21 3.065 7.22 3.465 ;
      RECT 7.2 3.059 7.21 3.453 ;
      RECT 7.19 3.053 7.2 3.433 ;
      RECT 7.185 3.049 7.19 3.418 ;
      RECT 7.18 3.047 7.185 3.41 ;
      RECT 7.175 3.045 7.18 3.403 ;
      RECT 7.17 3.043 7.175 3.393 ;
      RECT 7.165 3.041 7.17 3.387 ;
      RECT 7.155 3.04 7.165 3.377 ;
      RECT 7.145 3.04 7.155 3.368 ;
      RECT 7.13 3.04 7.145 3.353 ;
      RECT 7.09 3.04 7.12 3.337 ;
      RECT 7.07 3.042 7.09 3.332 ;
      RECT 7.065 3.047 7.07 3.33 ;
      RECT 7.035 3.055 7.065 3.328 ;
      RECT 7.005 3.07 7.035 3.327 ;
      RECT 6.96 3.092 7.005 3.332 ;
      RECT 6.955 3.107 6.96 3.336 ;
      RECT 6.94 3.112 6.955 3.338 ;
      RECT 6.935 3.116 6.94 3.34 ;
      RECT 6.875 3.139 6.935 3.349 ;
      RECT 6.855 3.165 6.875 3.362 ;
      RECT 6.845 3.172 6.855 3.366 ;
      RECT 6.83 3.179 6.845 3.369 ;
      RECT 6.81 3.189 6.83 3.372 ;
      RECT 6.805 3.197 6.81 3.375 ;
      RECT 6.76 3.202 6.805 3.382 ;
      RECT 6.75 3.205 6.76 3.389 ;
      RECT 6.74 3.205 6.75 3.393 ;
      RECT 6.705 3.207 6.74 3.405 ;
      RECT 6.685 3.21 6.705 3.418 ;
      RECT 6.645 3.213 6.685 3.429 ;
      RECT 6.63 3.215 6.645 3.442 ;
      RECT 6.62 3.215 6.63 3.447 ;
      RECT 6.595 3.216 6.62 3.455 ;
      RECT 6.585 3.218 6.595 3.46 ;
      RECT 6.58 3.219 6.585 3.463 ;
      RECT 6.555 3.217 6.58 3.466 ;
      RECT 6.54 3.215 6.555 3.467 ;
      RECT 6.52 3.212 6.54 3.469 ;
      RECT 6.5 3.207 6.52 3.469 ;
      RECT 6.44 3.202 6.5 3.466 ;
      RECT 6.405 3.177 6.44 3.462 ;
      RECT 6.395 3.154 6.405 3.46 ;
      RECT 6.365 3.131 6.395 3.46 ;
      RECT 6.355 3.11 6.365 3.46 ;
      RECT 6.33 3.092 6.355 3.458 ;
      RECT 6.315 3.07 6.33 3.455 ;
      RECT 6.3 3.052 6.315 3.453 ;
      RECT 6.28 3.042 6.3 3.451 ;
      RECT 6.265 3.037 6.28 3.45 ;
      RECT 6.25 3.035 6.265 3.449 ;
      RECT 6.22 3.036 6.25 3.447 ;
      RECT 6.2 3.039 6.22 3.445 ;
      RECT 6.143 3.043 6.2 3.445 ;
      RECT 6.057 3.052 6.143 3.445 ;
      RECT 5.971 3.063 6.057 3.445 ;
      RECT 5.885 3.074 5.971 3.445 ;
      RECT 5.865 3.081 5.885 3.453 ;
      RECT 5.855 3.084 5.865 3.46 ;
      RECT 5.79 3.089 5.855 3.478 ;
      RECT 5.76 3.096 5.79 3.503 ;
      RECT 5.75 3.099 5.76 3.51 ;
      RECT 5.705 3.103 5.75 3.515 ;
      RECT 5.675 3.108 5.705 3.52 ;
      RECT 5.674 3.11 5.675 3.52 ;
      RECT 5.588 3.116 5.674 3.52 ;
      RECT 5.502 3.127 5.588 3.52 ;
      RECT 5.416 3.139 5.502 3.52 ;
      RECT 5.33 3.15 5.416 3.52 ;
      RECT 5.315 3.157 5.33 3.515 ;
      RECT 5.31 3.159 5.315 3.509 ;
      RECT 5.29 3.17 5.31 3.504 ;
      RECT 5.28 3.188 5.29 3.498 ;
      RECT 5.275 3.2 5.28 3.298 ;
      RECT 7.57 1.953 7.59 2.04 ;
      RECT 7.565 1.888 7.57 2.072 ;
      RECT 7.555 1.855 7.565 2.077 ;
      RECT 7.55 1.835 7.555 2.083 ;
      RECT 7.52 1.835 7.55 2.1 ;
      RECT 7.471 1.835 7.52 2.136 ;
      RECT 7.385 1.835 7.471 2.194 ;
      RECT 7.356 1.845 7.385 2.243 ;
      RECT 7.27 1.887 7.356 2.296 ;
      RECT 7.25 1.925 7.27 2.343 ;
      RECT 7.225 1.942 7.25 2.363 ;
      RECT 7.215 1.956 7.225 2.383 ;
      RECT 7.21 1.962 7.215 2.393 ;
      RECT 7.205 1.966 7.21 2.4 ;
      RECT 7.155 1.986 7.205 2.405 ;
      RECT 7.09 2.03 7.155 2.405 ;
      RECT 7.065 2.08 7.09 2.405 ;
      RECT 7.055 2.11 7.065 2.405 ;
      RECT 7.05 2.137 7.055 2.405 ;
      RECT 7.045 2.155 7.05 2.405 ;
      RECT 7.035 2.197 7.045 2.405 ;
      RECT 7.385 2.755 7.555 2.93 ;
      RECT 7.325 2.583 7.385 2.918 ;
      RECT 7.315 2.576 7.325 2.901 ;
      RECT 7.27 2.755 7.555 2.881 ;
      RECT 7.251 2.755 7.555 2.859 ;
      RECT 7.165 2.755 7.555 2.824 ;
      RECT 7.145 2.575 7.315 2.78 ;
      RECT 7.145 2.722 7.55 2.78 ;
      RECT 7.145 2.67 7.525 2.78 ;
      RECT 7.145 2.625 7.49 2.78 ;
      RECT 7.145 2.607 7.455 2.78 ;
      RECT 7.145 2.597 7.45 2.78 ;
      RECT 6.865 3.555 7.055 3.78 ;
      RECT 6.855 3.556 7.06 3.775 ;
      RECT 6.855 3.558 7.07 3.755 ;
      RECT 6.855 3.562 7.075 3.74 ;
      RECT 6.855 3.549 7.025 3.775 ;
      RECT 6.855 3.552 7.05 3.775 ;
      RECT 6.865 3.548 7.025 3.78 ;
      RECT 6.951 3.546 7.025 3.78 ;
      RECT 6.575 2.797 6.745 3.035 ;
      RECT 6.575 2.797 6.831 2.949 ;
      RECT 6.575 2.797 6.835 2.859 ;
      RECT 6.625 2.57 6.845 2.838 ;
      RECT 6.62 2.587 6.85 2.811 ;
      RECT 6.585 2.745 6.85 2.811 ;
      RECT 6.605 2.595 6.745 3.035 ;
      RECT 6.595 2.677 6.855 2.794 ;
      RECT 6.59 2.725 6.855 2.794 ;
      RECT 6.595 2.635 6.85 2.811 ;
      RECT 6.62 2.572 6.845 2.838 ;
      RECT 6.185 2.547 6.355 2.745 ;
      RECT 6.185 2.547 6.4 2.72 ;
      RECT 6.255 2.49 6.425 2.678 ;
      RECT 6.23 2.505 6.425 2.678 ;
      RECT 5.845 2.551 5.875 2.745 ;
      RECT 5.84 2.523 5.845 2.745 ;
      RECT 5.81 2.497 5.84 2.747 ;
      RECT 5.785 2.455 5.81 2.75 ;
      RECT 5.775 2.427 5.785 2.752 ;
      RECT 5.74 2.407 5.775 2.754 ;
      RECT 5.675 2.392 5.74 2.76 ;
      RECT 5.625 2.39 5.675 2.766 ;
      RECT 5.602 2.392 5.625 2.771 ;
      RECT 5.516 2.403 5.602 2.777 ;
      RECT 5.43 2.421 5.516 2.787 ;
      RECT 5.415 2.432 5.43 2.793 ;
      RECT 5.345 2.455 5.415 2.799 ;
      RECT 5.29 2.487 5.345 2.807 ;
      RECT 5.25 2.51 5.29 2.813 ;
      RECT 5.236 2.523 5.25 2.816 ;
      RECT 5.15 2.545 5.236 2.822 ;
      RECT 5.135 2.57 5.15 2.828 ;
      RECT 5.095 2.585 5.135 2.832 ;
      RECT 5.045 2.6 5.095 2.837 ;
      RECT 5.02 2.607 5.045 2.841 ;
      RECT 4.96 2.602 5.02 2.845 ;
      RECT 4.945 2.593 4.96 2.849 ;
      RECT 4.875 2.583 4.945 2.845 ;
      RECT 4.85 2.575 4.87 2.835 ;
      RECT 4.791 2.575 4.85 2.813 ;
      RECT 4.705 2.575 4.791 2.77 ;
      RECT 4.87 2.575 4.875 2.84 ;
      RECT 5.565 1.806 5.735 2.14 ;
      RECT 5.535 1.806 5.735 2.135 ;
      RECT 5.475 1.773 5.535 2.123 ;
      RECT 5.475 1.829 5.745 2.118 ;
      RECT 5.45 1.829 5.745 2.112 ;
      RECT 5.445 1.77 5.475 2.109 ;
      RECT 5.43 1.776 5.565 2.107 ;
      RECT 5.425 1.784 5.65 2.095 ;
      RECT 5.425 1.836 5.76 2.048 ;
      RECT 5.41 1.792 5.65 2.043 ;
      RECT 5.41 1.862 5.77 1.984 ;
      RECT 5.38 1.812 5.735 1.945 ;
      RECT 5.38 1.902 5.78 1.941 ;
      RECT 5.43 1.781 5.65 2.107 ;
      RECT 4.77 2.111 4.825 2.375 ;
      RECT 4.77 2.111 4.89 2.374 ;
      RECT 4.77 2.111 4.915 2.373 ;
      RECT 4.77 2.111 4.98 2.372 ;
      RECT 4.915 2.077 4.995 2.371 ;
      RECT 4.73 2.121 5.14 2.37 ;
      RECT 4.77 2.118 5.14 2.37 ;
      RECT 4.73 2.126 5.145 2.363 ;
      RECT 4.715 2.128 5.145 2.362 ;
      RECT 4.715 2.135 5.15 2.358 ;
      RECT 4.695 2.134 5.145 2.354 ;
      RECT 4.695 2.142 5.155 2.353 ;
      RECT 4.69 2.139 5.15 2.349 ;
      RECT 4.69 2.152 5.165 2.348 ;
      RECT 4.675 2.142 5.155 2.347 ;
      RECT 4.64 2.155 5.165 2.34 ;
      RECT 4.825 2.11 5.135 2.37 ;
      RECT 4.825 2.095 5.085 2.37 ;
      RECT 4.89 2.082 5.02 2.37 ;
      RECT 4.435 3.171 4.45 3.564 ;
      RECT 4.4 3.176 4.45 3.563 ;
      RECT 4.435 3.175 4.495 3.562 ;
      RECT 4.38 3.186 4.495 3.561 ;
      RECT 4.395 3.182 4.495 3.561 ;
      RECT 4.36 3.192 4.57 3.558 ;
      RECT 4.36 3.211 4.615 3.556 ;
      RECT 4.36 3.218 4.62 3.553 ;
      RECT 4.345 3.195 4.57 3.55 ;
      RECT 4.325 3.2 4.57 3.543 ;
      RECT 4.32 3.204 4.57 3.539 ;
      RECT 4.32 3.221 4.63 3.538 ;
      RECT 4.3 3.215 4.615 3.534 ;
      RECT 4.3 3.224 4.635 3.528 ;
      RECT 4.295 3.23 4.635 3.3 ;
      RECT 4.36 3.19 4.495 3.558 ;
      RECT 4.235 2.553 4.435 2.865 ;
      RECT 4.31 2.531 4.435 2.865 ;
      RECT 4.25 2.55 4.44 2.85 ;
      RECT 4.22 2.561 4.44 2.848 ;
      RECT 4.235 2.556 4.445 2.814 ;
      RECT 4.22 2.66 4.45 2.781 ;
      RECT 4.25 2.532 4.435 2.865 ;
      RECT 4.31 2.51 4.41 2.865 ;
      RECT 4.335 2.507 4.41 2.865 ;
      RECT 4.335 2.502 4.355 2.865 ;
      RECT 3.74 2.57 3.915 2.745 ;
      RECT 3.735 2.57 3.915 2.743 ;
      RECT 3.71 2.57 3.915 2.738 ;
      RECT 3.655 2.55 3.825 2.728 ;
      RECT 3.655 2.557 3.89 2.728 ;
      RECT 3.74 3.237 3.755 3.42 ;
      RECT 3.73 3.215 3.74 3.42 ;
      RECT 3.715 3.195 3.73 3.42 ;
      RECT 3.705 3.17 3.715 3.42 ;
      RECT 3.675 3.135 3.705 3.42 ;
      RECT 3.64 3.075 3.675 3.42 ;
      RECT 3.635 3.037 3.64 3.42 ;
      RECT 3.585 2.988 3.635 3.42 ;
      RECT 3.575 2.938 3.585 3.408 ;
      RECT 3.56 2.917 3.575 3.368 ;
      RECT 3.54 2.885 3.56 3.318 ;
      RECT 3.515 2.841 3.54 3.258 ;
      RECT 3.51 2.813 3.515 3.213 ;
      RECT 3.505 2.804 3.51 3.199 ;
      RECT 3.5 2.797 3.505 3.186 ;
      RECT 3.495 2.792 3.5 3.175 ;
      RECT 3.49 2.777 3.495 3.165 ;
      RECT 3.485 2.755 3.49 3.152 ;
      RECT 3.475 2.715 3.485 3.127 ;
      RECT 3.45 2.645 3.475 3.083 ;
      RECT 3.445 2.585 3.45 3.048 ;
      RECT 3.43 2.565 3.445 3.015 ;
      RECT 3.425 2.565 3.43 2.99 ;
      RECT 3.395 2.565 3.425 2.945 ;
      RECT 3.35 2.565 3.395 2.885 ;
      RECT 3.275 2.565 3.35 2.833 ;
      RECT 3.27 2.565 3.275 2.798 ;
      RECT 3.265 2.565 3.27 2.788 ;
      RECT 3.26 2.565 3.265 2.768 ;
      RECT 3.525 1.785 3.695 2.255 ;
      RECT 3.47 1.778 3.665 2.239 ;
      RECT 3.47 1.792 3.7 2.238 ;
      RECT 3.455 1.793 3.7 2.219 ;
      RECT 3.45 1.811 3.7 2.205 ;
      RECT 3.455 1.794 3.705 2.203 ;
      RECT 3.44 1.825 3.705 2.188 ;
      RECT 3.455 1.8 3.71 2.173 ;
      RECT 3.435 1.84 3.71 2.17 ;
      RECT 3.45 1.812 3.715 2.155 ;
      RECT 3.45 1.824 3.72 2.135 ;
      RECT 3.435 1.84 3.725 2.118 ;
      RECT 3.435 1.85 3.73 1.973 ;
      RECT 3.43 1.85 3.73 1.93 ;
      RECT 3.43 1.865 3.735 1.908 ;
      RECT 3.525 1.775 3.665 2.255 ;
      RECT 3.525 1.773 3.635 2.255 ;
      RECT 3.611 1.77 3.635 2.255 ;
      RECT 3.27 3.437 3.275 3.483 ;
      RECT 3.26 3.285 3.27 3.507 ;
      RECT 3.255 3.13 3.26 3.532 ;
      RECT 3.24 3.092 3.255 3.543 ;
      RECT 3.235 3.075 3.24 3.55 ;
      RECT 3.225 3.063 3.235 3.557 ;
      RECT 3.22 3.054 3.225 3.559 ;
      RECT 3.215 3.052 3.22 3.563 ;
      RECT 3.17 3.043 3.215 3.578 ;
      RECT 3.165 3.035 3.17 3.592 ;
      RECT 3.16 3.032 3.165 3.596 ;
      RECT 3.145 3.027 3.16 3.604 ;
      RECT 3.09 3.017 3.145 3.615 ;
      RECT 3.055 3.005 3.09 3.616 ;
      RECT 3.046 3 3.055 3.61 ;
      RECT 2.96 3 3.046 3.6 ;
      RECT 2.93 3 2.96 3.578 ;
      RECT 2.92 3 2.925 3.558 ;
      RECT 2.915 3 2.92 3.52 ;
      RECT 2.91 3 2.915 3.478 ;
      RECT 2.905 3 2.91 3.438 ;
      RECT 2.9 3 2.905 3.368 ;
      RECT 2.89 3 2.9 3.29 ;
      RECT 2.885 3 2.89 3.19 ;
      RECT 2.925 3 2.93 3.56 ;
      RECT 2.42 3.082 2.51 3.56 ;
      RECT 2.405 3.085 2.525 3.558 ;
      RECT 2.42 3.084 2.525 3.558 ;
      RECT 2.385 3.091 2.55 3.548 ;
      RECT 2.405 3.085 2.55 3.548 ;
      RECT 2.37 3.097 2.55 3.536 ;
      RECT 2.405 3.088 2.6 3.529 ;
      RECT 2.356 3.105 2.6 3.527 ;
      RECT 2.385 3.095 2.61 3.515 ;
      RECT 2.356 3.116 2.64 3.506 ;
      RECT 2.27 3.14 2.64 3.5 ;
      RECT 2.27 3.153 2.68 3.483 ;
      RECT 2.265 3.175 2.68 3.476 ;
      RECT 2.235 3.19 2.68 3.466 ;
      RECT 2.23 3.201 2.68 3.456 ;
      RECT 2.2 3.214 2.68 3.447 ;
      RECT 2.185 3.232 2.68 3.436 ;
      RECT 2.16 3.245 2.68 3.426 ;
      RECT 2.42 3.081 2.43 3.56 ;
      RECT 2.466 2.505 2.505 2.75 ;
      RECT 2.38 2.505 2.515 2.748 ;
      RECT 2.265 2.53 2.515 2.745 ;
      RECT 2.265 2.53 2.52 2.743 ;
      RECT 2.265 2.53 2.535 2.738 ;
      RECT 2.371 2.505 2.55 2.718 ;
      RECT 2.285 2.513 2.55 2.718 ;
      RECT 1.955 1.865 2.125 2.3 ;
      RECT 1.945 1.899 2.125 2.283 ;
      RECT 2.025 1.835 2.195 2.27 ;
      RECT 1.93 1.91 2.195 2.248 ;
      RECT 2.025 1.845 2.2 2.238 ;
      RECT 1.955 1.897 2.23 2.223 ;
      RECT 1.915 1.923 2.23 2.208 ;
      RECT 1.915 1.965 2.24 2.188 ;
      RECT 1.91 1.99 2.245 2.17 ;
      RECT 1.91 2 2.25 2.155 ;
      RECT 1.905 1.937 2.23 2.153 ;
      RECT 1.905 2.01 2.255 2.138 ;
      RECT 1.9 1.947 2.23 2.135 ;
      RECT 1.895 2.031 2.26 2.118 ;
      RECT 1.895 2.063 2.265 2.098 ;
      RECT 1.89 1.977 2.24 2.09 ;
      RECT 1.895 1.962 2.23 2.118 ;
      RECT 1.91 1.932 2.23 2.17 ;
      RECT 1.755 2.519 1.98 2.775 ;
      RECT 1.755 2.552 2 2.765 ;
      RECT 1.72 2.552 2 2.763 ;
      RECT 1.72 2.565 2.005 2.753 ;
      RECT 1.72 2.585 2.015 2.745 ;
      RECT 1.72 2.682 2.02 2.738 ;
      RECT 1.7 2.43 1.83 2.728 ;
      RECT 1.655 2.585 2.015 2.67 ;
      RECT 1.645 2.43 1.83 2.615 ;
      RECT 1.645 2.462 1.916 2.615 ;
      RECT 1.61 2.992 1.63 3.17 ;
      RECT 1.575 2.945 1.61 3.17 ;
      RECT 1.56 2.885 1.575 3.17 ;
      RECT 1.535 2.832 1.56 3.17 ;
      RECT 1.52 2.785 1.535 3.17 ;
      RECT 1.5 2.762 1.52 3.17 ;
      RECT 1.475 2.727 1.5 3.17 ;
      RECT 1.465 2.573 1.475 3.17 ;
      RECT 1.435 2.568 1.465 3.161 ;
      RECT 1.43 2.565 1.435 3.151 ;
      RECT 1.415 2.565 1.43 3.125 ;
      RECT 1.41 2.565 1.415 3.088 ;
      RECT 1.385 2.565 1.41 3.04 ;
      RECT 1.365 2.565 1.385 2.965 ;
      RECT 1.355 2.565 1.365 2.925 ;
      RECT 1.35 2.565 1.355 2.9 ;
      RECT 1.345 2.565 1.35 2.883 ;
      RECT 1.34 2.565 1.345 2.865 ;
      RECT 1.335 2.566 1.34 2.855 ;
      RECT 1.325 2.568 1.335 2.823 ;
      RECT 1.315 2.57 1.325 2.79 ;
      RECT 1.305 2.573 1.315 2.763 ;
      RECT 1.63 3 1.855 3.17 ;
      RECT 0.96 1.812 1.13 2.265 ;
      RECT 0.96 1.812 1.22 2.231 ;
      RECT 0.96 1.812 1.25 2.215 ;
      RECT 0.96 1.812 1.28 2.188 ;
      RECT 1.216 1.79 1.295 2.17 ;
      RECT 0.995 1.797 1.3 2.155 ;
      RECT 0.995 1.805 1.31 2.118 ;
      RECT 0.955 1.832 1.31 2.09 ;
      RECT 0.94 1.845 1.31 2.055 ;
      RECT 0.96 1.82 1.33 2.045 ;
      RECT 0.935 1.885 1.33 2.015 ;
      RECT 0.935 1.915 1.335 1.998 ;
      RECT 0.93 1.945 1.335 1.985 ;
      RECT 0.995 1.794 1.295 2.17 ;
      RECT 1.13 1.791 1.216 2.249 ;
      RECT 1.081 1.792 1.295 2.17 ;
      RECT 1.225 3.452 1.27 3.645 ;
      RECT 1.215 3.422 1.225 3.645 ;
      RECT 1.21 3.407 1.215 3.645 ;
      RECT 1.17 3.317 1.21 3.645 ;
      RECT 1.165 3.23 1.17 3.645 ;
      RECT 1.155 3.2 1.165 3.645 ;
      RECT 1.15 3.16 1.155 3.645 ;
      RECT 1.14 3.122 1.15 3.645 ;
      RECT 1.135 3.087 1.14 3.645 ;
      RECT 1.115 3.04 1.135 3.645 ;
      RECT 1.1 2.965 1.115 3.645 ;
      RECT 1.095 2.92 1.1 3.64 ;
      RECT 1.09 2.9 1.095 3.613 ;
      RECT 1.085 2.88 1.09 3.598 ;
      RECT 1.08 2.855 1.085 3.578 ;
      RECT 1.075 2.833 1.08 3.563 ;
      RECT 1.07 2.811 1.075 3.545 ;
      RECT 1.065 2.79 1.07 3.535 ;
      RECT 1.055 2.762 1.065 3.505 ;
      RECT 1.045 2.725 1.055 3.473 ;
      RECT 1.035 2.685 1.045 3.44 ;
      RECT 1.025 2.663 1.035 3.41 ;
      RECT 0.995 2.615 1.025 3.342 ;
      RECT 0.98 2.575 0.995 3.269 ;
      RECT 0.97 2.575 0.98 3.235 ;
      RECT 0.965 2.575 0.97 3.21 ;
      RECT 0.96 2.575 0.965 3.195 ;
      RECT 0.955 2.575 0.96 3.173 ;
      RECT 0.95 2.575 0.955 3.16 ;
      RECT 0.935 2.575 0.95 3.125 ;
      RECT 0.915 2.575 0.935 3.065 ;
      RECT 0.905 2.575 0.915 3.015 ;
      RECT 0.885 2.575 0.905 2.963 ;
      RECT 0.865 2.575 0.885 2.92 ;
      RECT 0.855 2.575 0.865 2.908 ;
      RECT 0.825 2.575 0.855 2.895 ;
      RECT 0.795 2.596 0.825 2.875 ;
      RECT 0.785 2.624 0.795 2.855 ;
      RECT 0.77 2.641 0.785 2.823 ;
      RECT 0.765 2.655 0.77 2.79 ;
      RECT 0.76 2.663 0.765 2.763 ;
      RECT 0.755 2.671 0.76 2.725 ;
      RECT 0.76 3.195 0.765 3.53 ;
      RECT 0.725 3.182 0.76 3.529 ;
      RECT 0.655 3.122 0.725 3.528 ;
      RECT 0.575 3.065 0.655 3.527 ;
      RECT 0.44 3.025 0.575 3.526 ;
      RECT 0.44 3.212 0.775 3.515 ;
      RECT 0.4 3.212 0.775 3.505 ;
      RECT 0.4 3.23 0.78 3.5 ;
      RECT 0.4 3.32 0.785 3.49 ;
      RECT 0.395 3.015 0.56 3.47 ;
      RECT 0.39 3.015 0.56 3.213 ;
      RECT 0.39 3.172 0.755 3.213 ;
      RECT 0.39 3.16 0.75 3.213 ;
      RECT 78.71 0.575 78.88 1.085 ;
      RECT 78.71 5.015 78.88 6.485 ;
      RECT 78.71 7.795 78.88 8.305 ;
      RECT 77.72 0.575 77.89 1.085 ;
      RECT 77.72 2.395 77.89 3.865 ;
      RECT 77.72 5.015 77.89 6.485 ;
      RECT 77.72 7.795 77.89 8.305 ;
      RECT 76.355 0.575 76.525 3.865 ;
      RECT 76.355 5.015 76.525 8.305 ;
      RECT 75.925 0.575 76.095 1.085 ;
      RECT 75.925 1.655 76.095 3.865 ;
      RECT 75.925 5.015 76.095 7.225 ;
      RECT 75.925 7.795 76.095 8.305 ;
      RECT 74.555 1.66 74.725 2.935 ;
      RECT 74.555 5.945 74.725 7.22 ;
      RECT 62.86 0.575 63.03 1.085 ;
      RECT 62.86 2.395 63.03 3.865 ;
      RECT 62.86 5.015 63.03 6.485 ;
      RECT 62.86 7.795 63.03 8.305 ;
      RECT 61.87 0.575 62.04 1.085 ;
      RECT 61.87 2.395 62.04 3.865 ;
      RECT 61.87 5.015 62.04 6.485 ;
      RECT 61.87 7.795 62.04 8.305 ;
      RECT 60.505 0.575 60.675 3.865 ;
      RECT 60.505 5.015 60.675 8.305 ;
      RECT 60.075 0.575 60.245 1.085 ;
      RECT 60.075 1.655 60.245 3.865 ;
      RECT 60.075 5.015 60.245 7.225 ;
      RECT 60.075 7.795 60.245 8.305 ;
      RECT 58.705 1.66 58.875 2.935 ;
      RECT 58.705 5.945 58.875 7.22 ;
      RECT 47.01 0.575 47.18 1.085 ;
      RECT 47.01 2.395 47.18 3.865 ;
      RECT 47.01 5.015 47.18 6.485 ;
      RECT 47.01 7.795 47.18 8.305 ;
      RECT 46.02 0.575 46.19 1.085 ;
      RECT 46.02 2.395 46.19 3.865 ;
      RECT 46.02 5.015 46.19 6.485 ;
      RECT 46.02 7.795 46.19 8.305 ;
      RECT 44.655 0.575 44.825 3.865 ;
      RECT 44.655 5.015 44.825 8.305 ;
      RECT 44.225 0.575 44.395 1.085 ;
      RECT 44.225 1.655 44.395 3.865 ;
      RECT 44.225 5.015 44.395 7.225 ;
      RECT 44.225 7.795 44.395 8.305 ;
      RECT 42.855 1.66 43.025 2.935 ;
      RECT 42.855 5.945 43.025 7.22 ;
      RECT 31.16 0.575 31.33 1.085 ;
      RECT 31.16 2.395 31.33 3.865 ;
      RECT 31.16 5.015 31.33 6.485 ;
      RECT 31.16 7.795 31.33 8.305 ;
      RECT 30.17 0.575 30.34 1.085 ;
      RECT 30.17 2.395 30.34 3.865 ;
      RECT 30.17 5.015 30.34 6.485 ;
      RECT 30.17 7.795 30.34 8.305 ;
      RECT 28.805 0.575 28.975 3.865 ;
      RECT 28.805 5.015 28.975 8.305 ;
      RECT 28.375 0.575 28.545 1.085 ;
      RECT 28.375 1.655 28.545 3.865 ;
      RECT 28.375 5.015 28.545 7.225 ;
      RECT 28.375 7.795 28.545 8.305 ;
      RECT 27.005 1.66 27.175 2.935 ;
      RECT 27.005 5.945 27.175 7.22 ;
      RECT 15.31 0.575 15.48 1.085 ;
      RECT 15.31 2.395 15.48 3.865 ;
      RECT 15.31 5.015 15.48 6.485 ;
      RECT 15.31 7.795 15.48 8.305 ;
      RECT 14.32 0.575 14.49 1.085 ;
      RECT 14.32 2.395 14.49 3.865 ;
      RECT 14.32 5.015 14.49 6.485 ;
      RECT 14.32 7.795 14.49 8.305 ;
      RECT 12.955 0.575 13.125 3.865 ;
      RECT 12.955 5.015 13.125 8.305 ;
      RECT 12.525 0.575 12.695 1.085 ;
      RECT 12.525 1.655 12.695 3.865 ;
      RECT 12.525 5.015 12.695 7.225 ;
      RECT 12.525 7.795 12.695 8.305 ;
      RECT 11.155 1.66 11.325 2.935 ;
      RECT 11.155 5.945 11.325 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2aa_8

MACRO sky130_osu_ring_oscillator_mpr2at_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2at_8 0 0 ;
  SIZE 89.605 BY 8.88 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT 81.36 3.685 81.915 4.015 ;
      RECT 81.36 2.02 81.66 4.015 ;
      RECT 77.425 3.125 77.98 3.455 ;
      RECT 77.68 2.02 77.98 3.455 ;
      RECT 78.475 1.885 78.625 2.535 ;
      RECT 77.68 2.02 81.66 2.32 ;
      RECT 63.44 3.685 63.995 4.015 ;
      RECT 63.44 2.02 63.74 4.015 ;
      RECT 59.505 3.125 60.06 3.455 ;
      RECT 59.76 2.02 60.06 3.455 ;
      RECT 60.555 1.885 60.705 2.535 ;
      RECT 59.76 2.02 63.74 2.32 ;
      RECT 45.52 3.685 46.075 4.015 ;
      RECT 45.52 2.02 45.82 4.015 ;
      RECT 41.585 3.125 42.14 3.455 ;
      RECT 41.84 2.02 42.14 3.455 ;
      RECT 42.635 1.885 42.785 2.535 ;
      RECT 41.84 2.02 45.82 2.32 ;
      RECT 27.605 3.685 28.16 4.015 ;
      RECT 27.605 2.02 27.905 4.015 ;
      RECT 23.67 3.125 24.225 3.455 ;
      RECT 23.925 2.02 24.225 3.455 ;
      RECT 24.72 1.885 24.87 2.535 ;
      RECT 23.925 2.02 27.905 2.32 ;
      RECT 9.685 3.685 10.24 4.015 ;
      RECT 9.685 2.02 9.985 4.015 ;
      RECT 5.75 3.125 6.305 3.455 ;
      RECT 6.005 2.02 6.305 3.455 ;
      RECT 6.8 1.885 6.95 2.535 ;
      RECT 6.005 2.02 9.985 2.32 ;
      RECT 82.545 2.005 83.275 2.335 ;
      RECT 80.325 3.685 81.055 4.015 ;
      RECT 78.625 3.685 79.355 4.015 ;
      RECT 76.185 2.565 76.915 2.895 ;
      RECT 74.745 3.125 75.475 3.455 ;
      RECT 73.67 2.565 74.4 2.895 ;
      RECT 72.635 2.565 73.365 2.895 ;
      RECT 72.305 3.685 73.035 4.015 ;
      RECT 64.625 2.005 65.355 2.335 ;
      RECT 62.405 3.685 63.135 4.015 ;
      RECT 60.705 3.685 61.435 4.015 ;
      RECT 58.265 2.565 58.995 2.895 ;
      RECT 56.825 3.125 57.555 3.455 ;
      RECT 55.75 2.565 56.48 2.895 ;
      RECT 54.715 2.565 55.445 2.895 ;
      RECT 54.385 3.685 55.115 4.015 ;
      RECT 46.705 2.005 47.435 2.335 ;
      RECT 44.485 3.685 45.215 4.015 ;
      RECT 42.785 3.685 43.515 4.015 ;
      RECT 40.345 2.565 41.075 2.895 ;
      RECT 38.905 3.125 39.635 3.455 ;
      RECT 37.83 2.565 38.56 2.895 ;
      RECT 36.795 2.565 37.525 2.895 ;
      RECT 36.465 3.685 37.195 4.015 ;
      RECT 28.79 2.005 29.52 2.335 ;
      RECT 26.57 3.685 27.3 4.015 ;
      RECT 24.87 3.685 25.6 4.015 ;
      RECT 22.43 2.565 23.16 2.895 ;
      RECT 20.99 3.125 21.72 3.455 ;
      RECT 19.915 2.565 20.645 2.895 ;
      RECT 18.88 2.565 19.61 2.895 ;
      RECT 18.55 3.685 19.28 4.015 ;
      RECT 10.87 2.005 11.6 2.335 ;
      RECT 8.65 3.685 9.38 4.015 ;
      RECT 6.95 3.685 7.68 4.015 ;
      RECT 4.51 2.565 5.24 2.895 ;
      RECT 3.07 3.125 3.8 3.455 ;
      RECT 1.995 2.565 2.725 2.895 ;
      RECT 0.96 2.565 1.69 2.895 ;
      RECT 0.63 3.685 1.36 4.015 ;
    LAYER via2 ;
      RECT 82.61 2.07 82.81 2.27 ;
      RECT 81.65 3.75 81.85 3.95 ;
      RECT 80.65 3.75 80.85 3.95 ;
      RECT 78.69 3.75 78.89 3.95 ;
      RECT 77.49 3.19 77.69 3.39 ;
      RECT 76.25 2.63 76.45 2.83 ;
      RECT 74.81 3.19 75.01 3.39 ;
      RECT 74.07 2.63 74.27 2.83 ;
      RECT 72.85 2.63 73.05 2.83 ;
      RECT 72.37 3.75 72.57 3.95 ;
      RECT 64.69 2.07 64.89 2.27 ;
      RECT 63.73 3.75 63.93 3.95 ;
      RECT 62.73 3.75 62.93 3.95 ;
      RECT 60.77 3.75 60.97 3.95 ;
      RECT 59.57 3.19 59.77 3.39 ;
      RECT 58.33 2.63 58.53 2.83 ;
      RECT 56.89 3.19 57.09 3.39 ;
      RECT 56.15 2.63 56.35 2.83 ;
      RECT 54.93 2.63 55.13 2.83 ;
      RECT 54.45 3.75 54.65 3.95 ;
      RECT 46.77 2.07 46.97 2.27 ;
      RECT 45.81 3.75 46.01 3.95 ;
      RECT 44.81 3.75 45.01 3.95 ;
      RECT 42.85 3.75 43.05 3.95 ;
      RECT 41.65 3.19 41.85 3.39 ;
      RECT 40.41 2.63 40.61 2.83 ;
      RECT 38.97 3.19 39.17 3.39 ;
      RECT 38.23 2.63 38.43 2.83 ;
      RECT 37.01 2.63 37.21 2.83 ;
      RECT 36.53 3.75 36.73 3.95 ;
      RECT 28.855 2.07 29.055 2.27 ;
      RECT 27.895 3.75 28.095 3.95 ;
      RECT 26.895 3.75 27.095 3.95 ;
      RECT 24.935 3.75 25.135 3.95 ;
      RECT 23.735 3.19 23.935 3.39 ;
      RECT 22.495 2.63 22.695 2.83 ;
      RECT 21.055 3.19 21.255 3.39 ;
      RECT 20.315 2.63 20.515 2.83 ;
      RECT 19.095 2.63 19.295 2.83 ;
      RECT 18.615 3.75 18.815 3.95 ;
      RECT 10.935 2.07 11.135 2.27 ;
      RECT 9.975 3.75 10.175 3.95 ;
      RECT 8.975 3.75 9.175 3.95 ;
      RECT 7.015 3.75 7.215 3.95 ;
      RECT 5.815 3.19 6.015 3.39 ;
      RECT 4.575 2.63 4.775 2.83 ;
      RECT 3.135 3.19 3.335 3.39 ;
      RECT 2.395 2.63 2.595 2.83 ;
      RECT 1.175 2.63 1.375 2.83 ;
      RECT 0.695 3.75 0.895 3.95 ;
    LAYER met2 ;
      RECT 14.2 6.28 14.52 6.605 ;
      RECT 14.23 5.695 14.4 6.605 ;
      RECT 14.23 5.695 14.405 6.045 ;
      RECT 14.23 5.695 15.205 5.87 ;
      RECT 15.03 1.965 15.205 5.87 ;
      RECT 2.365 2.59 2.56 3.375 ;
      RECT 2.39 1.47 2.56 3.375 ;
      RECT 2.3 3.115 2.36 3.375 ;
      RECT 3.67 2.635 3.93 2.895 ;
      RECT 2.355 2.59 2.56 2.87 ;
      RECT 3.665 2.645 3.93 2.83 ;
      RECT 3.38 2.62 3.39 2.77 ;
      RECT 14.975 1.965 15.325 2.315 ;
      RECT 12.69 2.025 15.325 2.195 ;
      RECT 12.69 1.47 12.86 2.195 ;
      RECT 12.65 0.105 12.84 1.65 ;
      RECT 2.39 1.47 12.86 1.64 ;
      RECT 89.03 1.1 89.38 1.45 ;
      RECT 89.065 0.105 89.255 1.45 ;
      RECT 12.65 0.105 89.255 0.295 ;
      RECT 3.655 2.645 3.665 2.829 ;
      RECT 3.645 2.644 3.655 2.826 ;
      RECT 3.636 2.643 3.645 2.824 ;
      RECT 3.55 2.639 3.636 2.814 ;
      RECT 3.476 2.631 3.55 2.796 ;
      RECT 3.39 2.624 3.476 2.779 ;
      RECT 3.33 2.62 3.38 2.769 ;
      RECT 3.295 2.619 3.33 2.766 ;
      RECT 3.24 2.619 3.295 2.768 ;
      RECT 3.205 2.619 3.24 2.772 ;
      RECT 3.119 2.618 3.205 2.779 ;
      RECT 3.033 2.617 3.119 2.789 ;
      RECT 2.947 2.616 3.033 2.8 ;
      RECT 2.861 2.616 2.947 2.81 ;
      RECT 2.775 2.615 2.861 2.82 ;
      RECT 2.74 2.615 2.775 2.86 ;
      RECT 2.735 2.615 2.74 2.903 ;
      RECT 2.71 2.615 2.735 2.92 ;
      RECT 2.635 2.615 2.71 2.935 ;
      RECT 2.61 2.59 2.635 2.95 ;
      RECT 2.585 2.59 2.61 3 ;
      RECT 2.56 2.59 2.585 3.078 ;
      RECT 2.36 2.997 2.365 3.375 ;
      RECT 85.875 6.28 86.195 6.605 ;
      RECT 85.905 5.695 86.075 6.605 ;
      RECT 85.905 5.695 86.08 6.045 ;
      RECT 85.905 5.695 86.88 5.87 ;
      RECT 86.705 1.965 86.88 5.87 ;
      RECT 74.04 2.59 74.235 3.375 ;
      RECT 73.975 3.115 74.035 3.375 ;
      RECT 75.345 2.635 75.605 2.895 ;
      RECT 74.03 2.59 74.235 2.87 ;
      RECT 75.34 2.645 75.605 2.83 ;
      RECT 75.055 2.62 75.065 2.77 ;
      RECT 74.065 1.47 74.235 3.375 ;
      RECT 86.65 1.965 87 2.315 ;
      RECT 84.365 2.025 87 2.195 ;
      RECT 84.365 1.47 84.535 2.195 ;
      RECT 74.065 1.47 84.535 1.64 ;
      RECT 74.12 1.165 74.305 1.64 ;
      RECT 71.12 1.095 71.47 1.445 ;
      RECT 71.12 1.165 74.305 1.335 ;
      RECT 75.33 2.645 75.34 2.829 ;
      RECT 75.32 2.644 75.33 2.826 ;
      RECT 75.311 2.643 75.32 2.824 ;
      RECT 75.225 2.639 75.311 2.814 ;
      RECT 75.151 2.631 75.225 2.796 ;
      RECT 75.065 2.624 75.151 2.779 ;
      RECT 75.005 2.62 75.055 2.769 ;
      RECT 74.97 2.619 75.005 2.766 ;
      RECT 74.915 2.619 74.97 2.768 ;
      RECT 74.88 2.619 74.915 2.772 ;
      RECT 74.794 2.618 74.88 2.779 ;
      RECT 74.708 2.617 74.794 2.789 ;
      RECT 74.622 2.616 74.708 2.8 ;
      RECT 74.536 2.616 74.622 2.81 ;
      RECT 74.45 2.615 74.536 2.82 ;
      RECT 74.415 2.615 74.45 2.86 ;
      RECT 74.41 2.615 74.415 2.903 ;
      RECT 74.385 2.615 74.41 2.92 ;
      RECT 74.31 2.615 74.385 2.935 ;
      RECT 74.285 2.59 74.31 2.95 ;
      RECT 74.26 2.59 74.285 3 ;
      RECT 74.235 2.59 74.26 3.078 ;
      RECT 74.035 2.997 74.04 3.375 ;
      RECT 86.675 6.655 87 6.98 ;
      RECT 85.56 6.745 87 6.915 ;
      RECT 85.56 2.395 85.72 6.915 ;
      RECT 85.875 2.365 86.195 2.685 ;
      RECT 85.56 2.395 86.195 2.565 ;
      RECT 84.82 5.84 85.17 6.19 ;
      RECT 84.895 2.705 85.07 6.19 ;
      RECT 84.83 2.705 85.18 3.055 ;
      RECT 78.845 4.36 84.515 4.53 ;
      RECT 84.345 3.425 84.515 4.53 ;
      RECT 78.9 3.71 78.93 3.99 ;
      RECT 78.65 3.6 78.67 3.99 ;
      RECT 78.605 3.6 78.67 3.86 ;
      RECT 84.255 3.43 84.605 3.78 ;
      RECT 78.435 2.225 78.47 2.485 ;
      RECT 78.21 2.225 78.27 2.485 ;
      RECT 78.89 3.69 78.9 3.99 ;
      RECT 78.885 3.65 78.89 3.99 ;
      RECT 78.87 3.605 78.885 3.99 ;
      RECT 78.865 3.57 78.87 3.99 ;
      RECT 78.86 3.55 78.865 3.99 ;
      RECT 78.845 3.508 78.86 3.99 ;
      RECT 78.83 3.446 78.845 4.53 ;
      RECT 78.81 3.375 78.83 4.53 ;
      RECT 78.8 3.305 78.81 4.53 ;
      RECT 78.755 3.245 78.8 4.53 ;
      RECT 78.675 3.207 78.755 4.53 ;
      RECT 78.67 3.198 78.675 3.99 ;
      RECT 78.665 3.197 78.67 3.57 ;
      RECT 78.655 3.196 78.665 3.553 ;
      RECT 78.63 3.177 78.655 3.523 ;
      RECT 78.625 3.152 78.63 3.502 ;
      RECT 78.615 3.13 78.625 3.493 ;
      RECT 78.61 3.101 78.615 3.483 ;
      RECT 78.57 3.027 78.61 3.455 ;
      RECT 78.55 2.928 78.57 3.42 ;
      RECT 78.535 2.864 78.55 3.403 ;
      RECT 78.505 2.788 78.535 3.375 ;
      RECT 78.485 2.703 78.505 3.348 ;
      RECT 78.445 2.599 78.485 3.255 ;
      RECT 78.44 2.52 78.445 3.163 ;
      RECT 78.435 2.503 78.44 3.14 ;
      RECT 78.43 2.225 78.435 3.12 ;
      RECT 78.4 2.225 78.43 3.058 ;
      RECT 78.395 2.225 78.4 2.99 ;
      RECT 78.385 2.225 78.395 2.955 ;
      RECT 78.375 2.225 78.385 2.92 ;
      RECT 78.31 2.225 78.375 2.775 ;
      RECT 78.305 2.225 78.31 2.645 ;
      RECT 78.275 2.225 78.305 2.578 ;
      RECT 78.27 2.225 78.275 2.503 ;
      RECT 82.605 2.16 82.865 2.42 ;
      RECT 82.6 2.16 82.865 2.368 ;
      RECT 82.595 2.16 82.865 2.338 ;
      RECT 82.57 2.03 82.85 2.31 ;
      RECT 81.61 3.71 81.89 3.99 ;
      RECT 81.65 3.665 81.915 3.925 ;
      RECT 81.64 3.7 81.915 3.925 ;
      RECT 81.645 3.685 81.89 3.99 ;
      RECT 81.65 3.662 81.86 3.99 ;
      RECT 81.65 3.66 81.845 3.99 ;
      RECT 81.69 3.65 81.845 3.99 ;
      RECT 81.66 3.655 81.845 3.99 ;
      RECT 81.69 3.647 81.79 3.99 ;
      RECT 81.715 3.64 81.79 3.99 ;
      RECT 81.695 3.642 81.79 3.99 ;
      RECT 81.025 3.155 81.285 3.415 ;
      RECT 81.075 3.147 81.265 3.415 ;
      RECT 81.08 3.067 81.265 3.415 ;
      RECT 81.2 2.455 81.265 3.415 ;
      RECT 81.105 2.852 81.265 3.415 ;
      RECT 81.18 2.54 81.265 3.415 ;
      RECT 81.215 2.165 81.351 2.893 ;
      RECT 81.16 2.662 81.351 2.893 ;
      RECT 81.175 2.602 81.265 3.415 ;
      RECT 81.215 2.165 81.375 2.558 ;
      RECT 81.215 2.165 81.385 2.455 ;
      RECT 81.205 2.165 81.465 2.425 ;
      RECT 80.61 3.71 80.89 3.99 ;
      RECT 80.63 3.67 80.89 3.99 ;
      RECT 80.27 3.625 80.375 3.885 ;
      RECT 80.125 2.115 80.215 2.375 ;
      RECT 80.665 3.18 80.67 3.22 ;
      RECT 80.66 3.17 80.665 3.305 ;
      RECT 80.655 3.16 80.66 3.398 ;
      RECT 80.645 3.14 80.655 3.454 ;
      RECT 80.565 3.068 80.645 3.534 ;
      RECT 80.6 3.712 80.61 3.937 ;
      RECT 80.595 3.709 80.6 3.932 ;
      RECT 80.58 3.706 80.595 3.925 ;
      RECT 80.545 3.7 80.58 3.907 ;
      RECT 80.56 3.003 80.565 3.608 ;
      RECT 80.54 2.954 80.56 3.623 ;
      RECT 80.53 3.687 80.545 3.89 ;
      RECT 80.535 2.896 80.54 3.638 ;
      RECT 80.53 2.874 80.535 3.648 ;
      RECT 80.495 2.784 80.53 3.885 ;
      RECT 80.48 2.662 80.495 3.885 ;
      RECT 80.475 2.615 80.48 3.885 ;
      RECT 80.45 2.54 80.475 3.885 ;
      RECT 80.435 2.455 80.45 3.885 ;
      RECT 80.43 2.402 80.435 3.885 ;
      RECT 80.425 2.382 80.43 3.885 ;
      RECT 80.42 2.357 80.425 3.119 ;
      RECT 80.405 3.317 80.425 3.885 ;
      RECT 80.415 2.335 80.42 3.096 ;
      RECT 80.405 2.287 80.415 3.061 ;
      RECT 80.4 2.25 80.405 3.027 ;
      RECT 80.4 3.397 80.405 3.885 ;
      RECT 80.385 2.227 80.4 2.982 ;
      RECT 80.38 3.495 80.4 3.885 ;
      RECT 80.33 2.115 80.385 2.824 ;
      RECT 80.375 3.617 80.38 3.885 ;
      RECT 80.315 2.115 80.33 2.663 ;
      RECT 80.31 2.115 80.315 2.615 ;
      RECT 80.305 2.115 80.31 2.603 ;
      RECT 80.26 2.115 80.305 2.54 ;
      RECT 80.235 2.115 80.26 2.458 ;
      RECT 80.22 2.115 80.235 2.41 ;
      RECT 80.215 2.115 80.22 2.38 ;
      RECT 79.54 3.565 79.585 3.825 ;
      RECT 79.445 2.1 79.59 2.36 ;
      RECT 79.95 2.722 79.96 2.813 ;
      RECT 79.935 2.66 79.95 2.869 ;
      RECT 79.93 2.607 79.935 2.915 ;
      RECT 79.88 2.554 79.93 3.041 ;
      RECT 79.875 2.509 79.88 3.188 ;
      RECT 79.865 2.497 79.875 3.23 ;
      RECT 79.83 2.461 79.865 3.335 ;
      RECT 79.825 2.429 79.83 3.441 ;
      RECT 79.81 2.411 79.825 3.486 ;
      RECT 79.805 2.394 79.81 2.72 ;
      RECT 79.8 2.775 79.81 3.543 ;
      RECT 79.795 2.38 79.805 2.693 ;
      RECT 79.79 2.83 79.8 3.825 ;
      RECT 79.785 2.366 79.795 2.678 ;
      RECT 79.785 2.88 79.79 3.825 ;
      RECT 79.77 2.343 79.785 2.658 ;
      RECT 79.75 3.002 79.785 3.825 ;
      RECT 79.765 2.325 79.77 2.64 ;
      RECT 79.76 2.317 79.765 2.63 ;
      RECT 79.73 2.285 79.76 2.594 ;
      RECT 79.74 3.13 79.75 3.825 ;
      RECT 79.735 3.157 79.74 3.825 ;
      RECT 79.73 3.207 79.735 3.825 ;
      RECT 79.72 2.251 79.73 2.559 ;
      RECT 79.68 3.275 79.73 3.825 ;
      RECT 79.705 2.228 79.72 2.535 ;
      RECT 79.68 2.1 79.705 2.498 ;
      RECT 79.675 2.1 79.68 2.47 ;
      RECT 79.645 3.375 79.68 3.825 ;
      RECT 79.67 2.1 79.675 2.463 ;
      RECT 79.665 2.1 79.67 2.453 ;
      RECT 79.65 2.1 79.665 2.438 ;
      RECT 79.635 2.1 79.65 2.41 ;
      RECT 79.6 3.48 79.645 3.825 ;
      RECT 79.62 2.1 79.635 2.383 ;
      RECT 79.59 2.1 79.62 2.368 ;
      RECT 79.585 3.552 79.6 3.825 ;
      RECT 79.51 2.635 79.55 2.895 ;
      RECT 79.285 2.582 79.29 2.84 ;
      RECT 75.24 2.06 75.5 2.32 ;
      RECT 75.24 2.085 75.515 2.3 ;
      RECT 77.63 1.91 77.635 2.055 ;
      RECT 79.5 2.63 79.51 2.895 ;
      RECT 79.48 2.622 79.5 2.895 ;
      RECT 79.462 2.618 79.48 2.895 ;
      RECT 79.376 2.607 79.462 2.895 ;
      RECT 79.29 2.59 79.376 2.895 ;
      RECT 79.235 2.577 79.285 2.825 ;
      RECT 79.201 2.569 79.235 2.8 ;
      RECT 79.115 2.558 79.201 2.765 ;
      RECT 79.08 2.535 79.115 2.73 ;
      RECT 79.07 2.497 79.08 2.716 ;
      RECT 79.065 2.47 79.07 2.712 ;
      RECT 79.06 2.457 79.065 2.709 ;
      RECT 79.05 2.437 79.06 2.705 ;
      RECT 79.045 2.412 79.05 2.701 ;
      RECT 79.02 2.367 79.045 2.695 ;
      RECT 79.01 2.308 79.02 2.687 ;
      RECT 79 2.276 79.01 2.678 ;
      RECT 78.98 2.228 79 2.658 ;
      RECT 78.975 2.188 78.98 2.628 ;
      RECT 78.96 2.162 78.975 2.602 ;
      RECT 78.955 2.14 78.96 2.578 ;
      RECT 78.94 2.112 78.955 2.554 ;
      RECT 78.925 2.085 78.94 2.518 ;
      RECT 78.91 2.062 78.925 2.48 ;
      RECT 78.905 2.052 78.91 2.455 ;
      RECT 78.895 2.045 78.905 2.438 ;
      RECT 78.88 2.032 78.895 2.408 ;
      RECT 78.875 2.022 78.88 2.383 ;
      RECT 78.87 2.017 78.875 2.37 ;
      RECT 78.86 2.01 78.87 2.35 ;
      RECT 78.855 2.003 78.86 2.335 ;
      RECT 78.83 1.996 78.855 2.293 ;
      RECT 78.815 1.986 78.83 2.243 ;
      RECT 78.805 1.981 78.815 2.213 ;
      RECT 78.795 1.977 78.805 2.188 ;
      RECT 78.78 1.974 78.795 2.178 ;
      RECT 78.73 1.971 78.78 2.163 ;
      RECT 78.71 1.969 78.73 2.148 ;
      RECT 78.661 1.967 78.71 2.143 ;
      RECT 78.575 1.963 78.661 2.138 ;
      RECT 78.536 1.96 78.575 2.134 ;
      RECT 78.45 1.956 78.536 2.129 ;
      RECT 78.4 1.953 78.45 2.123 ;
      RECT 78.351 1.95 78.4 2.118 ;
      RECT 78.265 1.947 78.351 2.113 ;
      RECT 78.261 1.945 78.265 2.11 ;
      RECT 78.175 1.942 78.261 2.105 ;
      RECT 78.126 1.938 78.175 2.098 ;
      RECT 78.04 1.935 78.126 2.093 ;
      RECT 78.016 1.932 78.04 2.089 ;
      RECT 77.93 1.93 78.016 2.084 ;
      RECT 77.865 1.926 77.93 2.077 ;
      RECT 77.862 1.925 77.865 2.074 ;
      RECT 77.776 1.922 77.862 2.071 ;
      RECT 77.69 1.916 77.776 2.064 ;
      RECT 77.66 1.912 77.69 2.06 ;
      RECT 77.635 1.91 77.66 2.058 ;
      RECT 77.58 1.907 77.63 2.055 ;
      RECT 77.5 1.906 77.58 2.055 ;
      RECT 77.445 1.908 77.5 2.058 ;
      RECT 77.43 1.909 77.445 2.062 ;
      RECT 77.375 1.917 77.43 2.072 ;
      RECT 77.345 1.925 77.375 2.085 ;
      RECT 77.326 1.926 77.345 2.091 ;
      RECT 77.24 1.929 77.326 2.096 ;
      RECT 77.17 1.934 77.24 2.105 ;
      RECT 77.151 1.937 77.17 2.111 ;
      RECT 77.065 1.941 77.151 2.116 ;
      RECT 77.025 1.945 77.065 2.123 ;
      RECT 77.016 1.947 77.025 2.126 ;
      RECT 76.93 1.951 77.016 2.131 ;
      RECT 76.927 1.954 76.93 2.135 ;
      RECT 76.841 1.957 76.927 2.139 ;
      RECT 76.755 1.963 76.841 2.147 ;
      RECT 76.731 1.967 76.755 2.151 ;
      RECT 76.645 1.971 76.731 2.156 ;
      RECT 76.6 1.976 76.645 2.163 ;
      RECT 76.52 1.981 76.6 2.17 ;
      RECT 76.44 1.987 76.52 2.185 ;
      RECT 76.415 1.991 76.44 2.198 ;
      RECT 76.35 1.994 76.415 2.21 ;
      RECT 76.295 1.999 76.35 2.225 ;
      RECT 76.265 2.002 76.295 2.243 ;
      RECT 76.255 2.004 76.265 2.256 ;
      RECT 76.195 2.019 76.255 2.266 ;
      RECT 76.18 2.036 76.195 2.275 ;
      RECT 76.175 2.045 76.18 2.275 ;
      RECT 76.165 2.055 76.175 2.275 ;
      RECT 76.155 2.072 76.165 2.275 ;
      RECT 76.135 2.082 76.155 2.276 ;
      RECT 76.09 2.092 76.135 2.277 ;
      RECT 76.055 2.101 76.09 2.279 ;
      RECT 75.99 2.106 76.055 2.281 ;
      RECT 75.91 2.107 75.99 2.284 ;
      RECT 75.906 2.105 75.91 2.285 ;
      RECT 75.82 2.102 75.906 2.287 ;
      RECT 75.773 2.099 75.82 2.289 ;
      RECT 75.687 2.095 75.773 2.292 ;
      RECT 75.601 2.091 75.687 2.295 ;
      RECT 75.515 2.087 75.601 2.299 ;
      RECT 77.45 3.15 77.73 3.43 ;
      RECT 77.49 3.13 77.75 3.39 ;
      RECT 77.48 3.14 77.75 3.39 ;
      RECT 77.49 3.067 77.705 3.43 ;
      RECT 77.545 2.99 77.7 3.43 ;
      RECT 77.55 2.775 77.7 3.43 ;
      RECT 77.54 2.577 77.69 2.828 ;
      RECT 77.53 2.577 77.69 2.695 ;
      RECT 77.525 2.455 77.685 2.598 ;
      RECT 77.51 2.455 77.685 2.503 ;
      RECT 77.505 2.165 77.68 2.48 ;
      RECT 77.49 2.165 77.68 2.45 ;
      RECT 77.45 2.165 77.71 2.425 ;
      RECT 77.36 3.635 77.44 3.895 ;
      RECT 76.765 2.355 76.77 2.62 ;
      RECT 76.645 2.355 76.77 2.615 ;
      RECT 77.32 3.6 77.36 3.895 ;
      RECT 77.275 3.522 77.32 3.895 ;
      RECT 77.255 3.45 77.275 3.895 ;
      RECT 77.245 3.402 77.255 3.895 ;
      RECT 77.21 3.335 77.245 3.895 ;
      RECT 77.18 3.235 77.21 3.895 ;
      RECT 77.16 3.16 77.18 3.695 ;
      RECT 77.15 3.11 77.16 3.65 ;
      RECT 77.145 3.087 77.15 3.623 ;
      RECT 77.14 3.072 77.145 3.61 ;
      RECT 77.135 3.057 77.14 3.588 ;
      RECT 77.13 3.042 77.135 3.57 ;
      RECT 77.105 2.997 77.13 3.525 ;
      RECT 77.095 2.945 77.105 3.468 ;
      RECT 77.085 2.915 77.095 3.435 ;
      RECT 77.075 2.88 77.085 3.403 ;
      RECT 77.04 2.812 77.075 3.335 ;
      RECT 77.035 2.751 77.04 3.27 ;
      RECT 77.025 2.739 77.035 3.25 ;
      RECT 77.02 2.727 77.025 3.23 ;
      RECT 77.015 2.719 77.02 3.218 ;
      RECT 77.01 2.711 77.015 3.198 ;
      RECT 77 2.699 77.01 3.17 ;
      RECT 76.99 2.683 77 3.14 ;
      RECT 76.965 2.655 76.99 3.078 ;
      RECT 76.955 2.626 76.965 3.023 ;
      RECT 76.94 2.605 76.955 2.983 ;
      RECT 76.935 2.589 76.94 2.955 ;
      RECT 76.93 2.577 76.935 2.945 ;
      RECT 76.925 2.572 76.93 2.918 ;
      RECT 76.92 2.565 76.925 2.905 ;
      RECT 76.905 2.548 76.92 2.878 ;
      RECT 76.895 2.355 76.905 2.838 ;
      RECT 76.885 2.355 76.895 2.805 ;
      RECT 76.875 2.355 76.885 2.78 ;
      RECT 76.805 2.355 76.875 2.715 ;
      RECT 76.795 2.355 76.805 2.663 ;
      RECT 76.78 2.355 76.795 2.645 ;
      RECT 76.77 2.355 76.78 2.63 ;
      RECT 76.6 3.225 76.86 3.485 ;
      RECT 75.135 3.26 75.14 3.467 ;
      RECT 74.77 3.15 74.845 3.465 ;
      RECT 74.585 3.205 74.74 3.465 ;
      RECT 74.77 3.15 74.875 3.43 ;
      RECT 76.585 3.322 76.6 3.483 ;
      RECT 76.56 3.33 76.585 3.488 ;
      RECT 76.535 3.337 76.56 3.493 ;
      RECT 76.472 3.348 76.535 3.502 ;
      RECT 76.386 3.367 76.472 3.519 ;
      RECT 76.3 3.389 76.386 3.538 ;
      RECT 76.285 3.402 76.3 3.549 ;
      RECT 76.245 3.41 76.285 3.556 ;
      RECT 76.225 3.415 76.245 3.563 ;
      RECT 76.187 3.416 76.225 3.566 ;
      RECT 76.101 3.419 76.187 3.567 ;
      RECT 76.015 3.423 76.101 3.568 ;
      RECT 75.966 3.425 76.015 3.57 ;
      RECT 75.88 3.425 75.966 3.572 ;
      RECT 75.84 3.42 75.88 3.574 ;
      RECT 75.83 3.414 75.84 3.575 ;
      RECT 75.79 3.409 75.83 3.572 ;
      RECT 75.78 3.402 75.79 3.568 ;
      RECT 75.765 3.398 75.78 3.566 ;
      RECT 75.748 3.394 75.765 3.564 ;
      RECT 75.662 3.384 75.748 3.556 ;
      RECT 75.576 3.366 75.662 3.542 ;
      RECT 75.49 3.349 75.576 3.528 ;
      RECT 75.465 3.337 75.49 3.519 ;
      RECT 75.395 3.327 75.465 3.512 ;
      RECT 75.35 3.315 75.395 3.503 ;
      RECT 75.29 3.302 75.35 3.495 ;
      RECT 75.285 3.294 75.29 3.49 ;
      RECT 75.25 3.289 75.285 3.488 ;
      RECT 75.195 3.28 75.25 3.481 ;
      RECT 75.155 3.269 75.195 3.473 ;
      RECT 75.14 3.262 75.155 3.469 ;
      RECT 75.12 3.255 75.135 3.466 ;
      RECT 75.105 3.245 75.12 3.464 ;
      RECT 75.09 3.232 75.105 3.461 ;
      RECT 75.065 3.215 75.09 3.457 ;
      RECT 75.05 3.197 75.065 3.454 ;
      RECT 75.025 3.15 75.05 3.452 ;
      RECT 75.001 3.15 75.025 3.449 ;
      RECT 74.915 3.15 75.001 3.441 ;
      RECT 74.875 3.15 74.915 3.433 ;
      RECT 74.74 3.197 74.77 3.465 ;
      RECT 76.42 2.78 76.68 3.04 ;
      RECT 76.38 2.78 76.68 2.918 ;
      RECT 76.345 2.78 76.68 2.903 ;
      RECT 76.29 2.78 76.68 2.883 ;
      RECT 76.21 2.59 76.49 2.87 ;
      RECT 76.21 2.772 76.56 2.87 ;
      RECT 76.21 2.715 76.545 2.87 ;
      RECT 76.21 2.662 76.495 2.87 ;
      RECT 73.37 2.949 73.385 3.405 ;
      RECT 73.365 3.021 73.471 3.403 ;
      RECT 73.385 2.115 73.52 3.401 ;
      RECT 73.37 2.965 73.525 3.4 ;
      RECT 73.37 3.015 73.53 3.398 ;
      RECT 73.355 3.08 73.53 3.397 ;
      RECT 73.365 3.072 73.535 3.394 ;
      RECT 73.345 3.12 73.535 3.389 ;
      RECT 73.345 3.12 73.55 3.386 ;
      RECT 73.34 3.12 73.55 3.383 ;
      RECT 73.315 3.12 73.575 3.38 ;
      RECT 73.385 2.115 73.545 2.768 ;
      RECT 73.38 2.115 73.545 2.74 ;
      RECT 73.375 2.115 73.545 2.568 ;
      RECT 73.375 2.115 73.565 2.508 ;
      RECT 73.33 2.115 73.59 2.375 ;
      RECT 72.81 2.59 73.09 2.87 ;
      RECT 72.8 2.605 73.09 2.865 ;
      RECT 72.755 2.667 73.09 2.863 ;
      RECT 72.83 2.582 72.995 2.87 ;
      RECT 72.83 2.567 72.951 2.87 ;
      RECT 72.865 2.56 72.951 2.87 ;
      RECT 72.33 3.71 72.61 3.99 ;
      RECT 72.29 3.672 72.585 3.783 ;
      RECT 72.275 3.622 72.565 3.678 ;
      RECT 72.22 3.385 72.48 3.645 ;
      RECT 72.22 3.587 72.56 3.645 ;
      RECT 72.22 3.527 72.555 3.645 ;
      RECT 72.22 3.477 72.535 3.645 ;
      RECT 72.22 3.457 72.53 3.645 ;
      RECT 72.22 3.435 72.525 3.645 ;
      RECT 72.22 3.42 72.495 3.645 ;
      RECT 67.955 6.28 68.275 6.605 ;
      RECT 67.985 5.695 68.155 6.605 ;
      RECT 67.985 5.695 68.16 6.045 ;
      RECT 67.985 5.695 68.96 5.87 ;
      RECT 68.785 1.965 68.96 5.87 ;
      RECT 56.12 2.59 56.315 3.375 ;
      RECT 56.055 3.115 56.115 3.375 ;
      RECT 57.425 2.635 57.685 2.895 ;
      RECT 56.11 2.59 56.315 2.87 ;
      RECT 57.42 2.645 57.685 2.83 ;
      RECT 57.135 2.62 57.145 2.77 ;
      RECT 56.145 1.47 56.315 3.375 ;
      RECT 68.73 1.965 69.08 2.315 ;
      RECT 66.445 2.025 69.08 2.195 ;
      RECT 66.445 1.47 66.615 2.195 ;
      RECT 56.145 1.47 66.615 1.64 ;
      RECT 56.19 1.17 56.36 1.64 ;
      RECT 53.195 1.1 53.545 1.45 ;
      RECT 53.195 1.17 56.36 1.34 ;
      RECT 57.41 2.645 57.42 2.829 ;
      RECT 57.4 2.644 57.41 2.826 ;
      RECT 57.391 2.643 57.4 2.824 ;
      RECT 57.305 2.639 57.391 2.814 ;
      RECT 57.231 2.631 57.305 2.796 ;
      RECT 57.145 2.624 57.231 2.779 ;
      RECT 57.085 2.62 57.135 2.769 ;
      RECT 57.05 2.619 57.085 2.766 ;
      RECT 56.995 2.619 57.05 2.768 ;
      RECT 56.96 2.619 56.995 2.772 ;
      RECT 56.874 2.618 56.96 2.779 ;
      RECT 56.788 2.617 56.874 2.789 ;
      RECT 56.702 2.616 56.788 2.8 ;
      RECT 56.616 2.616 56.702 2.81 ;
      RECT 56.53 2.615 56.616 2.82 ;
      RECT 56.495 2.615 56.53 2.86 ;
      RECT 56.49 2.615 56.495 2.903 ;
      RECT 56.465 2.615 56.49 2.92 ;
      RECT 56.39 2.615 56.465 2.935 ;
      RECT 56.365 2.59 56.39 2.95 ;
      RECT 56.34 2.59 56.365 3 ;
      RECT 56.315 2.59 56.34 3.078 ;
      RECT 56.115 2.997 56.12 3.375 ;
      RECT 68.755 6.655 69.08 6.98 ;
      RECT 67.64 6.745 69.08 6.915 ;
      RECT 67.64 2.395 67.8 6.915 ;
      RECT 67.955 2.365 68.275 2.685 ;
      RECT 67.64 2.395 68.275 2.565 ;
      RECT 66.9 5.84 67.25 6.19 ;
      RECT 66.975 2.705 67.15 6.19 ;
      RECT 66.91 2.705 67.26 3.055 ;
      RECT 60.925 4.36 66.595 4.53 ;
      RECT 66.425 3.425 66.595 4.53 ;
      RECT 60.98 3.71 61.01 3.99 ;
      RECT 60.73 3.6 60.75 3.99 ;
      RECT 60.685 3.6 60.75 3.86 ;
      RECT 66.335 3.43 66.685 3.78 ;
      RECT 60.515 2.225 60.55 2.485 ;
      RECT 60.29 2.225 60.35 2.485 ;
      RECT 60.97 3.69 60.98 3.99 ;
      RECT 60.965 3.65 60.97 3.99 ;
      RECT 60.95 3.605 60.965 3.99 ;
      RECT 60.945 3.57 60.95 3.99 ;
      RECT 60.94 3.55 60.945 3.99 ;
      RECT 60.925 3.508 60.94 3.99 ;
      RECT 60.91 3.446 60.925 4.53 ;
      RECT 60.89 3.375 60.91 4.53 ;
      RECT 60.88 3.305 60.89 4.53 ;
      RECT 60.835 3.245 60.88 4.53 ;
      RECT 60.755 3.207 60.835 4.53 ;
      RECT 60.75 3.198 60.755 3.99 ;
      RECT 60.745 3.197 60.75 3.57 ;
      RECT 60.735 3.196 60.745 3.553 ;
      RECT 60.71 3.177 60.735 3.523 ;
      RECT 60.705 3.152 60.71 3.502 ;
      RECT 60.695 3.13 60.705 3.493 ;
      RECT 60.69 3.101 60.695 3.483 ;
      RECT 60.65 3.027 60.69 3.455 ;
      RECT 60.63 2.928 60.65 3.42 ;
      RECT 60.615 2.864 60.63 3.403 ;
      RECT 60.585 2.788 60.615 3.375 ;
      RECT 60.565 2.703 60.585 3.348 ;
      RECT 60.525 2.599 60.565 3.255 ;
      RECT 60.52 2.52 60.525 3.163 ;
      RECT 60.515 2.503 60.52 3.14 ;
      RECT 60.51 2.225 60.515 3.12 ;
      RECT 60.48 2.225 60.51 3.058 ;
      RECT 60.475 2.225 60.48 2.99 ;
      RECT 60.465 2.225 60.475 2.955 ;
      RECT 60.455 2.225 60.465 2.92 ;
      RECT 60.39 2.225 60.455 2.775 ;
      RECT 60.385 2.225 60.39 2.645 ;
      RECT 60.355 2.225 60.385 2.578 ;
      RECT 60.35 2.225 60.355 2.503 ;
      RECT 64.685 2.16 64.945 2.42 ;
      RECT 64.68 2.16 64.945 2.368 ;
      RECT 64.675 2.16 64.945 2.338 ;
      RECT 64.65 2.03 64.93 2.31 ;
      RECT 63.69 3.71 63.97 3.99 ;
      RECT 63.73 3.665 63.995 3.925 ;
      RECT 63.72 3.7 63.995 3.925 ;
      RECT 63.725 3.685 63.97 3.99 ;
      RECT 63.73 3.662 63.94 3.99 ;
      RECT 63.73 3.66 63.925 3.99 ;
      RECT 63.77 3.65 63.925 3.99 ;
      RECT 63.74 3.655 63.925 3.99 ;
      RECT 63.77 3.647 63.87 3.99 ;
      RECT 63.795 3.64 63.87 3.99 ;
      RECT 63.775 3.642 63.87 3.99 ;
      RECT 63.105 3.155 63.365 3.415 ;
      RECT 63.155 3.147 63.345 3.415 ;
      RECT 63.16 3.067 63.345 3.415 ;
      RECT 63.28 2.455 63.345 3.415 ;
      RECT 63.185 2.852 63.345 3.415 ;
      RECT 63.26 2.54 63.345 3.415 ;
      RECT 63.295 2.165 63.431 2.893 ;
      RECT 63.24 2.662 63.431 2.893 ;
      RECT 63.255 2.602 63.345 3.415 ;
      RECT 63.295 2.165 63.455 2.558 ;
      RECT 63.295 2.165 63.465 2.455 ;
      RECT 63.285 2.165 63.545 2.425 ;
      RECT 62.69 3.71 62.97 3.99 ;
      RECT 62.71 3.67 62.97 3.99 ;
      RECT 62.35 3.625 62.455 3.885 ;
      RECT 62.205 2.115 62.295 2.375 ;
      RECT 62.745 3.18 62.75 3.22 ;
      RECT 62.74 3.17 62.745 3.305 ;
      RECT 62.735 3.16 62.74 3.398 ;
      RECT 62.725 3.14 62.735 3.454 ;
      RECT 62.645 3.068 62.725 3.534 ;
      RECT 62.68 3.712 62.69 3.937 ;
      RECT 62.675 3.709 62.68 3.932 ;
      RECT 62.66 3.706 62.675 3.925 ;
      RECT 62.625 3.7 62.66 3.907 ;
      RECT 62.64 3.003 62.645 3.608 ;
      RECT 62.62 2.954 62.64 3.623 ;
      RECT 62.61 3.687 62.625 3.89 ;
      RECT 62.615 2.896 62.62 3.638 ;
      RECT 62.61 2.874 62.615 3.648 ;
      RECT 62.575 2.784 62.61 3.885 ;
      RECT 62.56 2.662 62.575 3.885 ;
      RECT 62.555 2.615 62.56 3.885 ;
      RECT 62.53 2.54 62.555 3.885 ;
      RECT 62.515 2.455 62.53 3.885 ;
      RECT 62.51 2.402 62.515 3.885 ;
      RECT 62.505 2.382 62.51 3.885 ;
      RECT 62.5 2.357 62.505 3.119 ;
      RECT 62.485 3.317 62.505 3.885 ;
      RECT 62.495 2.335 62.5 3.096 ;
      RECT 62.485 2.287 62.495 3.061 ;
      RECT 62.48 2.25 62.485 3.027 ;
      RECT 62.48 3.397 62.485 3.885 ;
      RECT 62.465 2.227 62.48 2.982 ;
      RECT 62.46 3.495 62.48 3.885 ;
      RECT 62.41 2.115 62.465 2.824 ;
      RECT 62.455 3.617 62.46 3.885 ;
      RECT 62.395 2.115 62.41 2.663 ;
      RECT 62.39 2.115 62.395 2.615 ;
      RECT 62.385 2.115 62.39 2.603 ;
      RECT 62.34 2.115 62.385 2.54 ;
      RECT 62.315 2.115 62.34 2.458 ;
      RECT 62.3 2.115 62.315 2.41 ;
      RECT 62.295 2.115 62.3 2.38 ;
      RECT 61.62 3.565 61.665 3.825 ;
      RECT 61.525 2.1 61.67 2.36 ;
      RECT 62.03 2.722 62.04 2.813 ;
      RECT 62.015 2.66 62.03 2.869 ;
      RECT 62.01 2.607 62.015 2.915 ;
      RECT 61.96 2.554 62.01 3.041 ;
      RECT 61.955 2.509 61.96 3.188 ;
      RECT 61.945 2.497 61.955 3.23 ;
      RECT 61.91 2.461 61.945 3.335 ;
      RECT 61.905 2.429 61.91 3.441 ;
      RECT 61.89 2.411 61.905 3.486 ;
      RECT 61.885 2.394 61.89 2.72 ;
      RECT 61.88 2.775 61.89 3.543 ;
      RECT 61.875 2.38 61.885 2.693 ;
      RECT 61.87 2.83 61.88 3.825 ;
      RECT 61.865 2.366 61.875 2.678 ;
      RECT 61.865 2.88 61.87 3.825 ;
      RECT 61.85 2.343 61.865 2.658 ;
      RECT 61.83 3.002 61.865 3.825 ;
      RECT 61.845 2.325 61.85 2.64 ;
      RECT 61.84 2.317 61.845 2.63 ;
      RECT 61.81 2.285 61.84 2.594 ;
      RECT 61.82 3.13 61.83 3.825 ;
      RECT 61.815 3.157 61.82 3.825 ;
      RECT 61.81 3.207 61.815 3.825 ;
      RECT 61.8 2.251 61.81 2.559 ;
      RECT 61.76 3.275 61.81 3.825 ;
      RECT 61.785 2.228 61.8 2.535 ;
      RECT 61.76 2.1 61.785 2.498 ;
      RECT 61.755 2.1 61.76 2.47 ;
      RECT 61.725 3.375 61.76 3.825 ;
      RECT 61.75 2.1 61.755 2.463 ;
      RECT 61.745 2.1 61.75 2.453 ;
      RECT 61.73 2.1 61.745 2.438 ;
      RECT 61.715 2.1 61.73 2.41 ;
      RECT 61.68 3.48 61.725 3.825 ;
      RECT 61.7 2.1 61.715 2.383 ;
      RECT 61.67 2.1 61.7 2.368 ;
      RECT 61.665 3.552 61.68 3.825 ;
      RECT 61.59 2.635 61.63 2.895 ;
      RECT 61.365 2.582 61.37 2.84 ;
      RECT 57.32 2.06 57.58 2.32 ;
      RECT 57.32 2.085 57.595 2.3 ;
      RECT 59.71 1.91 59.715 2.055 ;
      RECT 61.58 2.63 61.59 2.895 ;
      RECT 61.56 2.622 61.58 2.895 ;
      RECT 61.542 2.618 61.56 2.895 ;
      RECT 61.456 2.607 61.542 2.895 ;
      RECT 61.37 2.59 61.456 2.895 ;
      RECT 61.315 2.577 61.365 2.825 ;
      RECT 61.281 2.569 61.315 2.8 ;
      RECT 61.195 2.558 61.281 2.765 ;
      RECT 61.16 2.535 61.195 2.73 ;
      RECT 61.15 2.497 61.16 2.716 ;
      RECT 61.145 2.47 61.15 2.712 ;
      RECT 61.14 2.457 61.145 2.709 ;
      RECT 61.13 2.437 61.14 2.705 ;
      RECT 61.125 2.412 61.13 2.701 ;
      RECT 61.1 2.367 61.125 2.695 ;
      RECT 61.09 2.308 61.1 2.687 ;
      RECT 61.08 2.276 61.09 2.678 ;
      RECT 61.06 2.228 61.08 2.658 ;
      RECT 61.055 2.188 61.06 2.628 ;
      RECT 61.04 2.162 61.055 2.602 ;
      RECT 61.035 2.14 61.04 2.578 ;
      RECT 61.02 2.112 61.035 2.554 ;
      RECT 61.005 2.085 61.02 2.518 ;
      RECT 60.99 2.062 61.005 2.48 ;
      RECT 60.985 2.052 60.99 2.455 ;
      RECT 60.975 2.045 60.985 2.438 ;
      RECT 60.96 2.032 60.975 2.408 ;
      RECT 60.955 2.022 60.96 2.383 ;
      RECT 60.95 2.017 60.955 2.37 ;
      RECT 60.94 2.01 60.95 2.35 ;
      RECT 60.935 2.003 60.94 2.335 ;
      RECT 60.91 1.996 60.935 2.293 ;
      RECT 60.895 1.986 60.91 2.243 ;
      RECT 60.885 1.981 60.895 2.213 ;
      RECT 60.875 1.977 60.885 2.188 ;
      RECT 60.86 1.974 60.875 2.178 ;
      RECT 60.81 1.971 60.86 2.163 ;
      RECT 60.79 1.969 60.81 2.148 ;
      RECT 60.741 1.967 60.79 2.143 ;
      RECT 60.655 1.963 60.741 2.138 ;
      RECT 60.616 1.96 60.655 2.134 ;
      RECT 60.53 1.956 60.616 2.129 ;
      RECT 60.48 1.953 60.53 2.123 ;
      RECT 60.431 1.95 60.48 2.118 ;
      RECT 60.345 1.947 60.431 2.113 ;
      RECT 60.341 1.945 60.345 2.11 ;
      RECT 60.255 1.942 60.341 2.105 ;
      RECT 60.206 1.938 60.255 2.098 ;
      RECT 60.12 1.935 60.206 2.093 ;
      RECT 60.096 1.932 60.12 2.089 ;
      RECT 60.01 1.93 60.096 2.084 ;
      RECT 59.945 1.926 60.01 2.077 ;
      RECT 59.942 1.925 59.945 2.074 ;
      RECT 59.856 1.922 59.942 2.071 ;
      RECT 59.77 1.916 59.856 2.064 ;
      RECT 59.74 1.912 59.77 2.06 ;
      RECT 59.715 1.91 59.74 2.058 ;
      RECT 59.66 1.907 59.71 2.055 ;
      RECT 59.58 1.906 59.66 2.055 ;
      RECT 59.525 1.908 59.58 2.058 ;
      RECT 59.51 1.909 59.525 2.062 ;
      RECT 59.455 1.917 59.51 2.072 ;
      RECT 59.425 1.925 59.455 2.085 ;
      RECT 59.406 1.926 59.425 2.091 ;
      RECT 59.32 1.929 59.406 2.096 ;
      RECT 59.25 1.934 59.32 2.105 ;
      RECT 59.231 1.937 59.25 2.111 ;
      RECT 59.145 1.941 59.231 2.116 ;
      RECT 59.105 1.945 59.145 2.123 ;
      RECT 59.096 1.947 59.105 2.126 ;
      RECT 59.01 1.951 59.096 2.131 ;
      RECT 59.007 1.954 59.01 2.135 ;
      RECT 58.921 1.957 59.007 2.139 ;
      RECT 58.835 1.963 58.921 2.147 ;
      RECT 58.811 1.967 58.835 2.151 ;
      RECT 58.725 1.971 58.811 2.156 ;
      RECT 58.68 1.976 58.725 2.163 ;
      RECT 58.6 1.981 58.68 2.17 ;
      RECT 58.52 1.987 58.6 2.185 ;
      RECT 58.495 1.991 58.52 2.198 ;
      RECT 58.43 1.994 58.495 2.21 ;
      RECT 58.375 1.999 58.43 2.225 ;
      RECT 58.345 2.002 58.375 2.243 ;
      RECT 58.335 2.004 58.345 2.256 ;
      RECT 58.275 2.019 58.335 2.266 ;
      RECT 58.26 2.036 58.275 2.275 ;
      RECT 58.255 2.045 58.26 2.275 ;
      RECT 58.245 2.055 58.255 2.275 ;
      RECT 58.235 2.072 58.245 2.275 ;
      RECT 58.215 2.082 58.235 2.276 ;
      RECT 58.17 2.092 58.215 2.277 ;
      RECT 58.135 2.101 58.17 2.279 ;
      RECT 58.07 2.106 58.135 2.281 ;
      RECT 57.99 2.107 58.07 2.284 ;
      RECT 57.986 2.105 57.99 2.285 ;
      RECT 57.9 2.102 57.986 2.287 ;
      RECT 57.853 2.099 57.9 2.289 ;
      RECT 57.767 2.095 57.853 2.292 ;
      RECT 57.681 2.091 57.767 2.295 ;
      RECT 57.595 2.087 57.681 2.299 ;
      RECT 59.53 3.15 59.81 3.43 ;
      RECT 59.57 3.13 59.83 3.39 ;
      RECT 59.56 3.14 59.83 3.39 ;
      RECT 59.57 3.067 59.785 3.43 ;
      RECT 59.625 2.99 59.78 3.43 ;
      RECT 59.63 2.775 59.78 3.43 ;
      RECT 59.62 2.577 59.77 2.828 ;
      RECT 59.61 2.577 59.77 2.695 ;
      RECT 59.605 2.455 59.765 2.598 ;
      RECT 59.59 2.455 59.765 2.503 ;
      RECT 59.585 2.165 59.76 2.48 ;
      RECT 59.57 2.165 59.76 2.45 ;
      RECT 59.53 2.165 59.79 2.425 ;
      RECT 59.44 3.635 59.52 3.895 ;
      RECT 58.845 2.355 58.85 2.62 ;
      RECT 58.725 2.355 58.85 2.615 ;
      RECT 59.4 3.6 59.44 3.895 ;
      RECT 59.355 3.522 59.4 3.895 ;
      RECT 59.335 3.45 59.355 3.895 ;
      RECT 59.325 3.402 59.335 3.895 ;
      RECT 59.29 3.335 59.325 3.895 ;
      RECT 59.26 3.235 59.29 3.895 ;
      RECT 59.24 3.16 59.26 3.695 ;
      RECT 59.23 3.11 59.24 3.65 ;
      RECT 59.225 3.087 59.23 3.623 ;
      RECT 59.22 3.072 59.225 3.61 ;
      RECT 59.215 3.057 59.22 3.588 ;
      RECT 59.21 3.042 59.215 3.57 ;
      RECT 59.185 2.997 59.21 3.525 ;
      RECT 59.175 2.945 59.185 3.468 ;
      RECT 59.165 2.915 59.175 3.435 ;
      RECT 59.155 2.88 59.165 3.403 ;
      RECT 59.12 2.812 59.155 3.335 ;
      RECT 59.115 2.751 59.12 3.27 ;
      RECT 59.105 2.739 59.115 3.25 ;
      RECT 59.1 2.727 59.105 3.23 ;
      RECT 59.095 2.719 59.1 3.218 ;
      RECT 59.09 2.711 59.095 3.198 ;
      RECT 59.08 2.699 59.09 3.17 ;
      RECT 59.07 2.683 59.08 3.14 ;
      RECT 59.045 2.655 59.07 3.078 ;
      RECT 59.035 2.626 59.045 3.023 ;
      RECT 59.02 2.605 59.035 2.983 ;
      RECT 59.015 2.589 59.02 2.955 ;
      RECT 59.01 2.577 59.015 2.945 ;
      RECT 59.005 2.572 59.01 2.918 ;
      RECT 59 2.565 59.005 2.905 ;
      RECT 58.985 2.548 59 2.878 ;
      RECT 58.975 2.355 58.985 2.838 ;
      RECT 58.965 2.355 58.975 2.805 ;
      RECT 58.955 2.355 58.965 2.78 ;
      RECT 58.885 2.355 58.955 2.715 ;
      RECT 58.875 2.355 58.885 2.663 ;
      RECT 58.86 2.355 58.875 2.645 ;
      RECT 58.85 2.355 58.86 2.63 ;
      RECT 58.68 3.225 58.94 3.485 ;
      RECT 57.215 3.26 57.22 3.467 ;
      RECT 56.85 3.15 56.925 3.465 ;
      RECT 56.665 3.205 56.82 3.465 ;
      RECT 56.85 3.15 56.955 3.43 ;
      RECT 58.665 3.322 58.68 3.483 ;
      RECT 58.64 3.33 58.665 3.488 ;
      RECT 58.615 3.337 58.64 3.493 ;
      RECT 58.552 3.348 58.615 3.502 ;
      RECT 58.466 3.367 58.552 3.519 ;
      RECT 58.38 3.389 58.466 3.538 ;
      RECT 58.365 3.402 58.38 3.549 ;
      RECT 58.325 3.41 58.365 3.556 ;
      RECT 58.305 3.415 58.325 3.563 ;
      RECT 58.267 3.416 58.305 3.566 ;
      RECT 58.181 3.419 58.267 3.567 ;
      RECT 58.095 3.423 58.181 3.568 ;
      RECT 58.046 3.425 58.095 3.57 ;
      RECT 57.96 3.425 58.046 3.572 ;
      RECT 57.92 3.42 57.96 3.574 ;
      RECT 57.91 3.414 57.92 3.575 ;
      RECT 57.87 3.409 57.91 3.572 ;
      RECT 57.86 3.402 57.87 3.568 ;
      RECT 57.845 3.398 57.86 3.566 ;
      RECT 57.828 3.394 57.845 3.564 ;
      RECT 57.742 3.384 57.828 3.556 ;
      RECT 57.656 3.366 57.742 3.542 ;
      RECT 57.57 3.349 57.656 3.528 ;
      RECT 57.545 3.337 57.57 3.519 ;
      RECT 57.475 3.327 57.545 3.512 ;
      RECT 57.43 3.315 57.475 3.503 ;
      RECT 57.37 3.302 57.43 3.495 ;
      RECT 57.365 3.294 57.37 3.49 ;
      RECT 57.33 3.289 57.365 3.488 ;
      RECT 57.275 3.28 57.33 3.481 ;
      RECT 57.235 3.269 57.275 3.473 ;
      RECT 57.22 3.262 57.235 3.469 ;
      RECT 57.2 3.255 57.215 3.466 ;
      RECT 57.185 3.245 57.2 3.464 ;
      RECT 57.17 3.232 57.185 3.461 ;
      RECT 57.145 3.215 57.17 3.457 ;
      RECT 57.13 3.197 57.145 3.454 ;
      RECT 57.105 3.15 57.13 3.452 ;
      RECT 57.081 3.15 57.105 3.449 ;
      RECT 56.995 3.15 57.081 3.441 ;
      RECT 56.955 3.15 56.995 3.433 ;
      RECT 56.82 3.197 56.85 3.465 ;
      RECT 58.5 2.78 58.76 3.04 ;
      RECT 58.46 2.78 58.76 2.918 ;
      RECT 58.425 2.78 58.76 2.903 ;
      RECT 58.37 2.78 58.76 2.883 ;
      RECT 58.29 2.59 58.57 2.87 ;
      RECT 58.29 2.772 58.64 2.87 ;
      RECT 58.29 2.715 58.625 2.87 ;
      RECT 58.29 2.662 58.575 2.87 ;
      RECT 55.45 2.949 55.465 3.405 ;
      RECT 55.445 3.021 55.551 3.403 ;
      RECT 55.465 2.115 55.6 3.401 ;
      RECT 55.45 2.965 55.605 3.4 ;
      RECT 55.45 3.015 55.61 3.398 ;
      RECT 55.435 3.08 55.61 3.397 ;
      RECT 55.445 3.072 55.615 3.394 ;
      RECT 55.425 3.12 55.615 3.389 ;
      RECT 55.425 3.12 55.63 3.386 ;
      RECT 55.42 3.12 55.63 3.383 ;
      RECT 55.395 3.12 55.655 3.38 ;
      RECT 55.465 2.115 55.625 2.768 ;
      RECT 55.46 2.115 55.625 2.74 ;
      RECT 55.455 2.115 55.625 2.568 ;
      RECT 55.455 2.115 55.645 2.508 ;
      RECT 55.41 2.115 55.67 2.375 ;
      RECT 54.89 2.59 55.17 2.87 ;
      RECT 54.88 2.605 55.17 2.865 ;
      RECT 54.835 2.667 55.17 2.863 ;
      RECT 54.91 2.582 55.075 2.87 ;
      RECT 54.91 2.567 55.031 2.87 ;
      RECT 54.945 2.56 55.031 2.87 ;
      RECT 54.41 3.71 54.69 3.99 ;
      RECT 54.37 3.672 54.665 3.783 ;
      RECT 54.355 3.622 54.645 3.678 ;
      RECT 54.3 3.385 54.56 3.645 ;
      RECT 54.3 3.587 54.64 3.645 ;
      RECT 54.3 3.527 54.635 3.645 ;
      RECT 54.3 3.477 54.615 3.645 ;
      RECT 54.3 3.457 54.61 3.645 ;
      RECT 54.3 3.435 54.605 3.645 ;
      RECT 54.3 3.42 54.575 3.645 ;
      RECT 50.035 6.28 50.355 6.605 ;
      RECT 50.065 5.695 50.235 6.605 ;
      RECT 50.065 5.695 50.24 6.045 ;
      RECT 50.065 5.695 51.04 5.87 ;
      RECT 50.865 1.965 51.04 5.87 ;
      RECT 38.2 2.59 38.395 3.375 ;
      RECT 38.135 3.115 38.195 3.375 ;
      RECT 39.505 2.635 39.765 2.895 ;
      RECT 38.19 2.59 38.395 2.87 ;
      RECT 39.5 2.645 39.765 2.83 ;
      RECT 39.215 2.62 39.225 2.77 ;
      RECT 38.225 1.47 38.395 3.375 ;
      RECT 50.81 1.965 51.16 2.315 ;
      RECT 48.525 2.025 51.16 2.195 ;
      RECT 48.525 1.47 48.695 2.195 ;
      RECT 38.225 1.47 48.695 1.64 ;
      RECT 38.28 1.165 38.475 1.64 ;
      RECT 35.275 1.095 35.625 1.445 ;
      RECT 35.275 1.165 38.475 1.335 ;
      RECT 39.49 2.645 39.5 2.829 ;
      RECT 39.48 2.644 39.49 2.826 ;
      RECT 39.471 2.643 39.48 2.824 ;
      RECT 39.385 2.639 39.471 2.814 ;
      RECT 39.311 2.631 39.385 2.796 ;
      RECT 39.225 2.624 39.311 2.779 ;
      RECT 39.165 2.62 39.215 2.769 ;
      RECT 39.13 2.619 39.165 2.766 ;
      RECT 39.075 2.619 39.13 2.768 ;
      RECT 39.04 2.619 39.075 2.772 ;
      RECT 38.954 2.618 39.04 2.779 ;
      RECT 38.868 2.617 38.954 2.789 ;
      RECT 38.782 2.616 38.868 2.8 ;
      RECT 38.696 2.616 38.782 2.81 ;
      RECT 38.61 2.615 38.696 2.82 ;
      RECT 38.575 2.615 38.61 2.86 ;
      RECT 38.57 2.615 38.575 2.903 ;
      RECT 38.545 2.615 38.57 2.92 ;
      RECT 38.47 2.615 38.545 2.935 ;
      RECT 38.445 2.59 38.47 2.95 ;
      RECT 38.42 2.59 38.445 3 ;
      RECT 38.395 2.59 38.42 3.078 ;
      RECT 38.195 2.997 38.2 3.375 ;
      RECT 50.835 6.655 51.16 6.98 ;
      RECT 49.72 6.745 51.16 6.915 ;
      RECT 49.72 2.395 49.88 6.915 ;
      RECT 50.035 2.365 50.355 2.685 ;
      RECT 49.72 2.395 50.355 2.565 ;
      RECT 48.98 5.84 49.33 6.19 ;
      RECT 49.055 2.705 49.23 6.19 ;
      RECT 48.99 2.705 49.34 3.055 ;
      RECT 43.005 4.36 48.675 4.53 ;
      RECT 48.505 3.425 48.675 4.53 ;
      RECT 43.06 3.71 43.09 3.99 ;
      RECT 42.81 3.6 42.83 3.99 ;
      RECT 42.765 3.6 42.83 3.86 ;
      RECT 48.415 3.43 48.765 3.78 ;
      RECT 42.595 2.225 42.63 2.485 ;
      RECT 42.37 2.225 42.43 2.485 ;
      RECT 43.05 3.69 43.06 3.99 ;
      RECT 43.045 3.65 43.05 3.99 ;
      RECT 43.03 3.605 43.045 3.99 ;
      RECT 43.025 3.57 43.03 3.99 ;
      RECT 43.02 3.55 43.025 3.99 ;
      RECT 43.005 3.508 43.02 3.99 ;
      RECT 42.99 3.446 43.005 4.53 ;
      RECT 42.97 3.375 42.99 4.53 ;
      RECT 42.96 3.305 42.97 4.53 ;
      RECT 42.915 3.245 42.96 4.53 ;
      RECT 42.835 3.207 42.915 4.53 ;
      RECT 42.83 3.198 42.835 3.99 ;
      RECT 42.825 3.197 42.83 3.57 ;
      RECT 42.815 3.196 42.825 3.553 ;
      RECT 42.79 3.177 42.815 3.523 ;
      RECT 42.785 3.152 42.79 3.502 ;
      RECT 42.775 3.13 42.785 3.493 ;
      RECT 42.77 3.101 42.775 3.483 ;
      RECT 42.73 3.027 42.77 3.455 ;
      RECT 42.71 2.928 42.73 3.42 ;
      RECT 42.695 2.864 42.71 3.403 ;
      RECT 42.665 2.788 42.695 3.375 ;
      RECT 42.645 2.703 42.665 3.348 ;
      RECT 42.605 2.599 42.645 3.255 ;
      RECT 42.6 2.52 42.605 3.163 ;
      RECT 42.595 2.503 42.6 3.14 ;
      RECT 42.59 2.225 42.595 3.12 ;
      RECT 42.56 2.225 42.59 3.058 ;
      RECT 42.555 2.225 42.56 2.99 ;
      RECT 42.545 2.225 42.555 2.955 ;
      RECT 42.535 2.225 42.545 2.92 ;
      RECT 42.47 2.225 42.535 2.775 ;
      RECT 42.465 2.225 42.47 2.645 ;
      RECT 42.435 2.225 42.465 2.578 ;
      RECT 42.43 2.225 42.435 2.503 ;
      RECT 46.765 2.16 47.025 2.42 ;
      RECT 46.76 2.16 47.025 2.368 ;
      RECT 46.755 2.16 47.025 2.338 ;
      RECT 46.73 2.03 47.01 2.31 ;
      RECT 45.77 3.71 46.05 3.99 ;
      RECT 45.81 3.665 46.075 3.925 ;
      RECT 45.8 3.7 46.075 3.925 ;
      RECT 45.805 3.685 46.05 3.99 ;
      RECT 45.81 3.662 46.02 3.99 ;
      RECT 45.81 3.66 46.005 3.99 ;
      RECT 45.85 3.65 46.005 3.99 ;
      RECT 45.82 3.655 46.005 3.99 ;
      RECT 45.85 3.647 45.95 3.99 ;
      RECT 45.875 3.64 45.95 3.99 ;
      RECT 45.855 3.642 45.95 3.99 ;
      RECT 45.185 3.155 45.445 3.415 ;
      RECT 45.235 3.147 45.425 3.415 ;
      RECT 45.24 3.067 45.425 3.415 ;
      RECT 45.36 2.455 45.425 3.415 ;
      RECT 45.265 2.852 45.425 3.415 ;
      RECT 45.34 2.54 45.425 3.415 ;
      RECT 45.375 2.165 45.511 2.893 ;
      RECT 45.32 2.662 45.511 2.893 ;
      RECT 45.335 2.602 45.425 3.415 ;
      RECT 45.375 2.165 45.535 2.558 ;
      RECT 45.375 2.165 45.545 2.455 ;
      RECT 45.365 2.165 45.625 2.425 ;
      RECT 44.77 3.71 45.05 3.99 ;
      RECT 44.79 3.67 45.05 3.99 ;
      RECT 44.43 3.625 44.535 3.885 ;
      RECT 44.285 2.115 44.375 2.375 ;
      RECT 44.825 3.18 44.83 3.22 ;
      RECT 44.82 3.17 44.825 3.305 ;
      RECT 44.815 3.16 44.82 3.398 ;
      RECT 44.805 3.14 44.815 3.454 ;
      RECT 44.725 3.068 44.805 3.534 ;
      RECT 44.76 3.712 44.77 3.937 ;
      RECT 44.755 3.709 44.76 3.932 ;
      RECT 44.74 3.706 44.755 3.925 ;
      RECT 44.705 3.7 44.74 3.907 ;
      RECT 44.72 3.003 44.725 3.608 ;
      RECT 44.7 2.954 44.72 3.623 ;
      RECT 44.69 3.687 44.705 3.89 ;
      RECT 44.695 2.896 44.7 3.638 ;
      RECT 44.69 2.874 44.695 3.648 ;
      RECT 44.655 2.784 44.69 3.885 ;
      RECT 44.64 2.662 44.655 3.885 ;
      RECT 44.635 2.615 44.64 3.885 ;
      RECT 44.61 2.54 44.635 3.885 ;
      RECT 44.595 2.455 44.61 3.885 ;
      RECT 44.59 2.402 44.595 3.885 ;
      RECT 44.585 2.382 44.59 3.885 ;
      RECT 44.58 2.357 44.585 3.119 ;
      RECT 44.565 3.317 44.585 3.885 ;
      RECT 44.575 2.335 44.58 3.096 ;
      RECT 44.565 2.287 44.575 3.061 ;
      RECT 44.56 2.25 44.565 3.027 ;
      RECT 44.56 3.397 44.565 3.885 ;
      RECT 44.545 2.227 44.56 2.982 ;
      RECT 44.54 3.495 44.56 3.885 ;
      RECT 44.49 2.115 44.545 2.824 ;
      RECT 44.535 3.617 44.54 3.885 ;
      RECT 44.475 2.115 44.49 2.663 ;
      RECT 44.47 2.115 44.475 2.615 ;
      RECT 44.465 2.115 44.47 2.603 ;
      RECT 44.42 2.115 44.465 2.54 ;
      RECT 44.395 2.115 44.42 2.458 ;
      RECT 44.38 2.115 44.395 2.41 ;
      RECT 44.375 2.115 44.38 2.38 ;
      RECT 43.7 3.565 43.745 3.825 ;
      RECT 43.605 2.1 43.75 2.36 ;
      RECT 44.11 2.722 44.12 2.813 ;
      RECT 44.095 2.66 44.11 2.869 ;
      RECT 44.09 2.607 44.095 2.915 ;
      RECT 44.04 2.554 44.09 3.041 ;
      RECT 44.035 2.509 44.04 3.188 ;
      RECT 44.025 2.497 44.035 3.23 ;
      RECT 43.99 2.461 44.025 3.335 ;
      RECT 43.985 2.429 43.99 3.441 ;
      RECT 43.97 2.411 43.985 3.486 ;
      RECT 43.965 2.394 43.97 2.72 ;
      RECT 43.96 2.775 43.97 3.543 ;
      RECT 43.955 2.38 43.965 2.693 ;
      RECT 43.95 2.83 43.96 3.825 ;
      RECT 43.945 2.366 43.955 2.678 ;
      RECT 43.945 2.88 43.95 3.825 ;
      RECT 43.93 2.343 43.945 2.658 ;
      RECT 43.91 3.002 43.945 3.825 ;
      RECT 43.925 2.325 43.93 2.64 ;
      RECT 43.92 2.317 43.925 2.63 ;
      RECT 43.89 2.285 43.92 2.594 ;
      RECT 43.9 3.13 43.91 3.825 ;
      RECT 43.895 3.157 43.9 3.825 ;
      RECT 43.89 3.207 43.895 3.825 ;
      RECT 43.88 2.251 43.89 2.559 ;
      RECT 43.84 3.275 43.89 3.825 ;
      RECT 43.865 2.228 43.88 2.535 ;
      RECT 43.84 2.1 43.865 2.498 ;
      RECT 43.835 2.1 43.84 2.47 ;
      RECT 43.805 3.375 43.84 3.825 ;
      RECT 43.83 2.1 43.835 2.463 ;
      RECT 43.825 2.1 43.83 2.453 ;
      RECT 43.81 2.1 43.825 2.438 ;
      RECT 43.795 2.1 43.81 2.41 ;
      RECT 43.76 3.48 43.805 3.825 ;
      RECT 43.78 2.1 43.795 2.383 ;
      RECT 43.75 2.1 43.78 2.368 ;
      RECT 43.745 3.552 43.76 3.825 ;
      RECT 43.67 2.635 43.71 2.895 ;
      RECT 43.445 2.582 43.45 2.84 ;
      RECT 39.4 2.06 39.66 2.32 ;
      RECT 39.4 2.085 39.675 2.3 ;
      RECT 41.79 1.91 41.795 2.055 ;
      RECT 43.66 2.63 43.67 2.895 ;
      RECT 43.64 2.622 43.66 2.895 ;
      RECT 43.622 2.618 43.64 2.895 ;
      RECT 43.536 2.607 43.622 2.895 ;
      RECT 43.45 2.59 43.536 2.895 ;
      RECT 43.395 2.577 43.445 2.825 ;
      RECT 43.361 2.569 43.395 2.8 ;
      RECT 43.275 2.558 43.361 2.765 ;
      RECT 43.24 2.535 43.275 2.73 ;
      RECT 43.23 2.497 43.24 2.716 ;
      RECT 43.225 2.47 43.23 2.712 ;
      RECT 43.22 2.457 43.225 2.709 ;
      RECT 43.21 2.437 43.22 2.705 ;
      RECT 43.205 2.412 43.21 2.701 ;
      RECT 43.18 2.367 43.205 2.695 ;
      RECT 43.17 2.308 43.18 2.687 ;
      RECT 43.16 2.276 43.17 2.678 ;
      RECT 43.14 2.228 43.16 2.658 ;
      RECT 43.135 2.188 43.14 2.628 ;
      RECT 43.12 2.162 43.135 2.602 ;
      RECT 43.115 2.14 43.12 2.578 ;
      RECT 43.1 2.112 43.115 2.554 ;
      RECT 43.085 2.085 43.1 2.518 ;
      RECT 43.07 2.062 43.085 2.48 ;
      RECT 43.065 2.052 43.07 2.455 ;
      RECT 43.055 2.045 43.065 2.438 ;
      RECT 43.04 2.032 43.055 2.408 ;
      RECT 43.035 2.022 43.04 2.383 ;
      RECT 43.03 2.017 43.035 2.37 ;
      RECT 43.02 2.01 43.03 2.35 ;
      RECT 43.015 2.003 43.02 2.335 ;
      RECT 42.99 1.996 43.015 2.293 ;
      RECT 42.975 1.986 42.99 2.243 ;
      RECT 42.965 1.981 42.975 2.213 ;
      RECT 42.955 1.977 42.965 2.188 ;
      RECT 42.94 1.974 42.955 2.178 ;
      RECT 42.89 1.971 42.94 2.163 ;
      RECT 42.87 1.969 42.89 2.148 ;
      RECT 42.821 1.967 42.87 2.143 ;
      RECT 42.735 1.963 42.821 2.138 ;
      RECT 42.696 1.96 42.735 2.134 ;
      RECT 42.61 1.956 42.696 2.129 ;
      RECT 42.56 1.953 42.61 2.123 ;
      RECT 42.511 1.95 42.56 2.118 ;
      RECT 42.425 1.947 42.511 2.113 ;
      RECT 42.421 1.945 42.425 2.11 ;
      RECT 42.335 1.942 42.421 2.105 ;
      RECT 42.286 1.938 42.335 2.098 ;
      RECT 42.2 1.935 42.286 2.093 ;
      RECT 42.176 1.932 42.2 2.089 ;
      RECT 42.09 1.93 42.176 2.084 ;
      RECT 42.025 1.926 42.09 2.077 ;
      RECT 42.022 1.925 42.025 2.074 ;
      RECT 41.936 1.922 42.022 2.071 ;
      RECT 41.85 1.916 41.936 2.064 ;
      RECT 41.82 1.912 41.85 2.06 ;
      RECT 41.795 1.91 41.82 2.058 ;
      RECT 41.74 1.907 41.79 2.055 ;
      RECT 41.66 1.906 41.74 2.055 ;
      RECT 41.605 1.908 41.66 2.058 ;
      RECT 41.59 1.909 41.605 2.062 ;
      RECT 41.535 1.917 41.59 2.072 ;
      RECT 41.505 1.925 41.535 2.085 ;
      RECT 41.486 1.926 41.505 2.091 ;
      RECT 41.4 1.929 41.486 2.096 ;
      RECT 41.33 1.934 41.4 2.105 ;
      RECT 41.311 1.937 41.33 2.111 ;
      RECT 41.225 1.941 41.311 2.116 ;
      RECT 41.185 1.945 41.225 2.123 ;
      RECT 41.176 1.947 41.185 2.126 ;
      RECT 41.09 1.951 41.176 2.131 ;
      RECT 41.087 1.954 41.09 2.135 ;
      RECT 41.001 1.957 41.087 2.139 ;
      RECT 40.915 1.963 41.001 2.147 ;
      RECT 40.891 1.967 40.915 2.151 ;
      RECT 40.805 1.971 40.891 2.156 ;
      RECT 40.76 1.976 40.805 2.163 ;
      RECT 40.68 1.981 40.76 2.17 ;
      RECT 40.6 1.987 40.68 2.185 ;
      RECT 40.575 1.991 40.6 2.198 ;
      RECT 40.51 1.994 40.575 2.21 ;
      RECT 40.455 1.999 40.51 2.225 ;
      RECT 40.425 2.002 40.455 2.243 ;
      RECT 40.415 2.004 40.425 2.256 ;
      RECT 40.355 2.019 40.415 2.266 ;
      RECT 40.34 2.036 40.355 2.275 ;
      RECT 40.335 2.045 40.34 2.275 ;
      RECT 40.325 2.055 40.335 2.275 ;
      RECT 40.315 2.072 40.325 2.275 ;
      RECT 40.295 2.082 40.315 2.276 ;
      RECT 40.25 2.092 40.295 2.277 ;
      RECT 40.215 2.101 40.25 2.279 ;
      RECT 40.15 2.106 40.215 2.281 ;
      RECT 40.07 2.107 40.15 2.284 ;
      RECT 40.066 2.105 40.07 2.285 ;
      RECT 39.98 2.102 40.066 2.287 ;
      RECT 39.933 2.099 39.98 2.289 ;
      RECT 39.847 2.095 39.933 2.292 ;
      RECT 39.761 2.091 39.847 2.295 ;
      RECT 39.675 2.087 39.761 2.299 ;
      RECT 41.61 3.15 41.89 3.43 ;
      RECT 41.65 3.13 41.91 3.39 ;
      RECT 41.64 3.14 41.91 3.39 ;
      RECT 41.65 3.067 41.865 3.43 ;
      RECT 41.705 2.99 41.86 3.43 ;
      RECT 41.71 2.775 41.86 3.43 ;
      RECT 41.7 2.577 41.85 2.828 ;
      RECT 41.69 2.577 41.85 2.695 ;
      RECT 41.685 2.455 41.845 2.598 ;
      RECT 41.67 2.455 41.845 2.503 ;
      RECT 41.665 2.165 41.84 2.48 ;
      RECT 41.65 2.165 41.84 2.45 ;
      RECT 41.61 2.165 41.87 2.425 ;
      RECT 41.52 3.635 41.6 3.895 ;
      RECT 40.925 2.355 40.93 2.62 ;
      RECT 40.805 2.355 40.93 2.615 ;
      RECT 41.48 3.6 41.52 3.895 ;
      RECT 41.435 3.522 41.48 3.895 ;
      RECT 41.415 3.45 41.435 3.895 ;
      RECT 41.405 3.402 41.415 3.895 ;
      RECT 41.37 3.335 41.405 3.895 ;
      RECT 41.34 3.235 41.37 3.895 ;
      RECT 41.32 3.16 41.34 3.695 ;
      RECT 41.31 3.11 41.32 3.65 ;
      RECT 41.305 3.087 41.31 3.623 ;
      RECT 41.3 3.072 41.305 3.61 ;
      RECT 41.295 3.057 41.3 3.588 ;
      RECT 41.29 3.042 41.295 3.57 ;
      RECT 41.265 2.997 41.29 3.525 ;
      RECT 41.255 2.945 41.265 3.468 ;
      RECT 41.245 2.915 41.255 3.435 ;
      RECT 41.235 2.88 41.245 3.403 ;
      RECT 41.2 2.812 41.235 3.335 ;
      RECT 41.195 2.751 41.2 3.27 ;
      RECT 41.185 2.739 41.195 3.25 ;
      RECT 41.18 2.727 41.185 3.23 ;
      RECT 41.175 2.719 41.18 3.218 ;
      RECT 41.17 2.711 41.175 3.198 ;
      RECT 41.16 2.699 41.17 3.17 ;
      RECT 41.15 2.683 41.16 3.14 ;
      RECT 41.125 2.655 41.15 3.078 ;
      RECT 41.115 2.626 41.125 3.023 ;
      RECT 41.1 2.605 41.115 2.983 ;
      RECT 41.095 2.589 41.1 2.955 ;
      RECT 41.09 2.577 41.095 2.945 ;
      RECT 41.085 2.572 41.09 2.918 ;
      RECT 41.08 2.565 41.085 2.905 ;
      RECT 41.065 2.548 41.08 2.878 ;
      RECT 41.055 2.355 41.065 2.838 ;
      RECT 41.045 2.355 41.055 2.805 ;
      RECT 41.035 2.355 41.045 2.78 ;
      RECT 40.965 2.355 41.035 2.715 ;
      RECT 40.955 2.355 40.965 2.663 ;
      RECT 40.94 2.355 40.955 2.645 ;
      RECT 40.93 2.355 40.94 2.63 ;
      RECT 40.76 3.225 41.02 3.485 ;
      RECT 39.295 3.26 39.3 3.467 ;
      RECT 38.93 3.15 39.005 3.465 ;
      RECT 38.745 3.205 38.9 3.465 ;
      RECT 38.93 3.15 39.035 3.43 ;
      RECT 40.745 3.322 40.76 3.483 ;
      RECT 40.72 3.33 40.745 3.488 ;
      RECT 40.695 3.337 40.72 3.493 ;
      RECT 40.632 3.348 40.695 3.502 ;
      RECT 40.546 3.367 40.632 3.519 ;
      RECT 40.46 3.389 40.546 3.538 ;
      RECT 40.445 3.402 40.46 3.549 ;
      RECT 40.405 3.41 40.445 3.556 ;
      RECT 40.385 3.415 40.405 3.563 ;
      RECT 40.347 3.416 40.385 3.566 ;
      RECT 40.261 3.419 40.347 3.567 ;
      RECT 40.175 3.423 40.261 3.568 ;
      RECT 40.126 3.425 40.175 3.57 ;
      RECT 40.04 3.425 40.126 3.572 ;
      RECT 40 3.42 40.04 3.574 ;
      RECT 39.99 3.414 40 3.575 ;
      RECT 39.95 3.409 39.99 3.572 ;
      RECT 39.94 3.402 39.95 3.568 ;
      RECT 39.925 3.398 39.94 3.566 ;
      RECT 39.908 3.394 39.925 3.564 ;
      RECT 39.822 3.384 39.908 3.556 ;
      RECT 39.736 3.366 39.822 3.542 ;
      RECT 39.65 3.349 39.736 3.528 ;
      RECT 39.625 3.337 39.65 3.519 ;
      RECT 39.555 3.327 39.625 3.512 ;
      RECT 39.51 3.315 39.555 3.503 ;
      RECT 39.45 3.302 39.51 3.495 ;
      RECT 39.445 3.294 39.45 3.49 ;
      RECT 39.41 3.289 39.445 3.488 ;
      RECT 39.355 3.28 39.41 3.481 ;
      RECT 39.315 3.269 39.355 3.473 ;
      RECT 39.3 3.262 39.315 3.469 ;
      RECT 39.28 3.255 39.295 3.466 ;
      RECT 39.265 3.245 39.28 3.464 ;
      RECT 39.25 3.232 39.265 3.461 ;
      RECT 39.225 3.215 39.25 3.457 ;
      RECT 39.21 3.197 39.225 3.454 ;
      RECT 39.185 3.15 39.21 3.452 ;
      RECT 39.161 3.15 39.185 3.449 ;
      RECT 39.075 3.15 39.161 3.441 ;
      RECT 39.035 3.15 39.075 3.433 ;
      RECT 38.9 3.197 38.93 3.465 ;
      RECT 40.58 2.78 40.84 3.04 ;
      RECT 40.54 2.78 40.84 2.918 ;
      RECT 40.505 2.78 40.84 2.903 ;
      RECT 40.45 2.78 40.84 2.883 ;
      RECT 40.37 2.59 40.65 2.87 ;
      RECT 40.37 2.772 40.72 2.87 ;
      RECT 40.37 2.715 40.705 2.87 ;
      RECT 40.37 2.662 40.655 2.87 ;
      RECT 37.53 2.949 37.545 3.405 ;
      RECT 37.525 3.021 37.631 3.403 ;
      RECT 37.545 2.115 37.68 3.401 ;
      RECT 37.53 2.965 37.685 3.4 ;
      RECT 37.53 3.015 37.69 3.398 ;
      RECT 37.515 3.08 37.69 3.397 ;
      RECT 37.525 3.072 37.695 3.394 ;
      RECT 37.505 3.12 37.695 3.389 ;
      RECT 37.505 3.12 37.71 3.386 ;
      RECT 37.5 3.12 37.71 3.383 ;
      RECT 37.475 3.12 37.735 3.38 ;
      RECT 37.545 2.115 37.705 2.768 ;
      RECT 37.54 2.115 37.705 2.74 ;
      RECT 37.535 2.115 37.705 2.568 ;
      RECT 37.535 2.115 37.725 2.508 ;
      RECT 37.49 2.115 37.75 2.375 ;
      RECT 36.97 2.59 37.25 2.87 ;
      RECT 36.96 2.605 37.25 2.865 ;
      RECT 36.915 2.667 37.25 2.863 ;
      RECT 36.99 2.582 37.155 2.87 ;
      RECT 36.99 2.567 37.111 2.87 ;
      RECT 37.025 2.56 37.111 2.87 ;
      RECT 36.49 3.71 36.77 3.99 ;
      RECT 36.45 3.672 36.745 3.783 ;
      RECT 36.435 3.622 36.725 3.678 ;
      RECT 36.38 3.385 36.64 3.645 ;
      RECT 36.38 3.587 36.72 3.645 ;
      RECT 36.38 3.527 36.715 3.645 ;
      RECT 36.38 3.477 36.695 3.645 ;
      RECT 36.38 3.457 36.69 3.645 ;
      RECT 36.38 3.435 36.685 3.645 ;
      RECT 36.38 3.42 36.655 3.645 ;
      RECT 32.12 6.28 32.44 6.605 ;
      RECT 32.15 5.695 32.32 6.605 ;
      RECT 32.15 5.695 32.325 6.045 ;
      RECT 32.15 5.695 33.125 5.87 ;
      RECT 32.95 1.965 33.125 5.87 ;
      RECT 20.285 2.59 20.48 3.375 ;
      RECT 20.22 3.115 20.28 3.375 ;
      RECT 21.59 2.635 21.85 2.895 ;
      RECT 20.275 2.59 20.48 2.87 ;
      RECT 21.585 2.645 21.85 2.83 ;
      RECT 21.3 2.62 21.31 2.77 ;
      RECT 20.31 1.47 20.48 3.375 ;
      RECT 32.895 1.965 33.245 2.315 ;
      RECT 30.61 2.025 33.245 2.195 ;
      RECT 30.61 1.47 30.78 2.195 ;
      RECT 20.31 1.47 30.78 1.64 ;
      RECT 20.365 1.165 20.56 1.64 ;
      RECT 17.305 1.095 17.655 1.445 ;
      RECT 17.305 1.165 20.56 1.335 ;
      RECT 21.575 2.645 21.585 2.829 ;
      RECT 21.565 2.644 21.575 2.826 ;
      RECT 21.556 2.643 21.565 2.824 ;
      RECT 21.47 2.639 21.556 2.814 ;
      RECT 21.396 2.631 21.47 2.796 ;
      RECT 21.31 2.624 21.396 2.779 ;
      RECT 21.25 2.62 21.3 2.769 ;
      RECT 21.215 2.619 21.25 2.766 ;
      RECT 21.16 2.619 21.215 2.768 ;
      RECT 21.125 2.619 21.16 2.772 ;
      RECT 21.039 2.618 21.125 2.779 ;
      RECT 20.953 2.617 21.039 2.789 ;
      RECT 20.867 2.616 20.953 2.8 ;
      RECT 20.781 2.616 20.867 2.81 ;
      RECT 20.695 2.615 20.781 2.82 ;
      RECT 20.66 2.615 20.695 2.86 ;
      RECT 20.655 2.615 20.66 2.903 ;
      RECT 20.63 2.615 20.655 2.92 ;
      RECT 20.555 2.615 20.63 2.935 ;
      RECT 20.53 2.59 20.555 2.95 ;
      RECT 20.505 2.59 20.53 3 ;
      RECT 20.48 2.59 20.505 3.078 ;
      RECT 20.28 2.997 20.285 3.375 ;
      RECT 32.92 6.655 33.245 6.98 ;
      RECT 31.805 6.745 33.245 6.915 ;
      RECT 31.805 2.395 31.965 6.915 ;
      RECT 32.12 2.365 32.44 2.685 ;
      RECT 31.805 2.395 32.44 2.565 ;
      RECT 31.065 5.84 31.415 6.19 ;
      RECT 31.14 2.705 31.315 6.19 ;
      RECT 31.075 2.705 31.425 3.055 ;
      RECT 25.09 4.36 30.76 4.53 ;
      RECT 30.59 3.425 30.76 4.53 ;
      RECT 25.145 3.71 25.175 3.99 ;
      RECT 24.895 3.6 24.915 3.99 ;
      RECT 24.85 3.6 24.915 3.86 ;
      RECT 30.5 3.43 30.85 3.78 ;
      RECT 24.68 2.225 24.715 2.485 ;
      RECT 24.455 2.225 24.515 2.485 ;
      RECT 25.135 3.69 25.145 3.99 ;
      RECT 25.13 3.65 25.135 3.99 ;
      RECT 25.115 3.605 25.13 3.99 ;
      RECT 25.11 3.57 25.115 3.99 ;
      RECT 25.105 3.55 25.11 3.99 ;
      RECT 25.09 3.508 25.105 3.99 ;
      RECT 25.075 3.446 25.09 4.53 ;
      RECT 25.055 3.375 25.075 4.53 ;
      RECT 25.045 3.305 25.055 4.53 ;
      RECT 25 3.245 25.045 4.53 ;
      RECT 24.92 3.207 25 4.53 ;
      RECT 24.915 3.198 24.92 3.99 ;
      RECT 24.91 3.197 24.915 3.57 ;
      RECT 24.9 3.196 24.91 3.553 ;
      RECT 24.875 3.177 24.9 3.523 ;
      RECT 24.87 3.152 24.875 3.502 ;
      RECT 24.86 3.13 24.87 3.493 ;
      RECT 24.855 3.101 24.86 3.483 ;
      RECT 24.815 3.027 24.855 3.455 ;
      RECT 24.795 2.928 24.815 3.42 ;
      RECT 24.78 2.864 24.795 3.403 ;
      RECT 24.75 2.788 24.78 3.375 ;
      RECT 24.73 2.703 24.75 3.348 ;
      RECT 24.69 2.599 24.73 3.255 ;
      RECT 24.685 2.52 24.69 3.163 ;
      RECT 24.68 2.503 24.685 3.14 ;
      RECT 24.675 2.225 24.68 3.12 ;
      RECT 24.645 2.225 24.675 3.058 ;
      RECT 24.64 2.225 24.645 2.99 ;
      RECT 24.63 2.225 24.64 2.955 ;
      RECT 24.62 2.225 24.63 2.92 ;
      RECT 24.555 2.225 24.62 2.775 ;
      RECT 24.55 2.225 24.555 2.645 ;
      RECT 24.52 2.225 24.55 2.578 ;
      RECT 24.515 2.225 24.52 2.503 ;
      RECT 28.85 2.16 29.11 2.42 ;
      RECT 28.845 2.16 29.11 2.368 ;
      RECT 28.84 2.16 29.11 2.338 ;
      RECT 28.815 2.03 29.095 2.31 ;
      RECT 27.855 3.71 28.135 3.99 ;
      RECT 27.895 3.665 28.16 3.925 ;
      RECT 27.885 3.7 28.16 3.925 ;
      RECT 27.89 3.685 28.135 3.99 ;
      RECT 27.895 3.662 28.105 3.99 ;
      RECT 27.895 3.66 28.09 3.99 ;
      RECT 27.935 3.65 28.09 3.99 ;
      RECT 27.905 3.655 28.09 3.99 ;
      RECT 27.935 3.647 28.035 3.99 ;
      RECT 27.96 3.64 28.035 3.99 ;
      RECT 27.94 3.642 28.035 3.99 ;
      RECT 27.27 3.155 27.53 3.415 ;
      RECT 27.32 3.147 27.51 3.415 ;
      RECT 27.325 3.067 27.51 3.415 ;
      RECT 27.445 2.455 27.51 3.415 ;
      RECT 27.35 2.852 27.51 3.415 ;
      RECT 27.425 2.54 27.51 3.415 ;
      RECT 27.46 2.165 27.596 2.893 ;
      RECT 27.405 2.662 27.596 2.893 ;
      RECT 27.42 2.602 27.51 3.415 ;
      RECT 27.46 2.165 27.62 2.558 ;
      RECT 27.46 2.165 27.63 2.455 ;
      RECT 27.45 2.165 27.71 2.425 ;
      RECT 26.855 3.71 27.135 3.99 ;
      RECT 26.875 3.67 27.135 3.99 ;
      RECT 26.515 3.625 26.62 3.885 ;
      RECT 26.37 2.115 26.46 2.375 ;
      RECT 26.91 3.18 26.915 3.22 ;
      RECT 26.905 3.17 26.91 3.305 ;
      RECT 26.9 3.16 26.905 3.398 ;
      RECT 26.89 3.14 26.9 3.454 ;
      RECT 26.81 3.068 26.89 3.534 ;
      RECT 26.845 3.712 26.855 3.937 ;
      RECT 26.84 3.709 26.845 3.932 ;
      RECT 26.825 3.706 26.84 3.925 ;
      RECT 26.79 3.7 26.825 3.907 ;
      RECT 26.805 3.003 26.81 3.608 ;
      RECT 26.785 2.954 26.805 3.623 ;
      RECT 26.775 3.687 26.79 3.89 ;
      RECT 26.78 2.896 26.785 3.638 ;
      RECT 26.775 2.874 26.78 3.648 ;
      RECT 26.74 2.784 26.775 3.885 ;
      RECT 26.725 2.662 26.74 3.885 ;
      RECT 26.72 2.615 26.725 3.885 ;
      RECT 26.695 2.54 26.72 3.885 ;
      RECT 26.68 2.455 26.695 3.885 ;
      RECT 26.675 2.402 26.68 3.885 ;
      RECT 26.67 2.382 26.675 3.885 ;
      RECT 26.665 2.357 26.67 3.119 ;
      RECT 26.65 3.317 26.67 3.885 ;
      RECT 26.66 2.335 26.665 3.096 ;
      RECT 26.65 2.287 26.66 3.061 ;
      RECT 26.645 2.25 26.65 3.027 ;
      RECT 26.645 3.397 26.65 3.885 ;
      RECT 26.63 2.227 26.645 2.982 ;
      RECT 26.625 3.495 26.645 3.885 ;
      RECT 26.575 2.115 26.63 2.824 ;
      RECT 26.62 3.617 26.625 3.885 ;
      RECT 26.56 2.115 26.575 2.663 ;
      RECT 26.555 2.115 26.56 2.615 ;
      RECT 26.55 2.115 26.555 2.603 ;
      RECT 26.505 2.115 26.55 2.54 ;
      RECT 26.48 2.115 26.505 2.458 ;
      RECT 26.465 2.115 26.48 2.41 ;
      RECT 26.46 2.115 26.465 2.38 ;
      RECT 25.785 3.565 25.83 3.825 ;
      RECT 25.69 2.1 25.835 2.36 ;
      RECT 26.195 2.722 26.205 2.813 ;
      RECT 26.18 2.66 26.195 2.869 ;
      RECT 26.175 2.607 26.18 2.915 ;
      RECT 26.125 2.554 26.175 3.041 ;
      RECT 26.12 2.509 26.125 3.188 ;
      RECT 26.11 2.497 26.12 3.23 ;
      RECT 26.075 2.461 26.11 3.335 ;
      RECT 26.07 2.429 26.075 3.441 ;
      RECT 26.055 2.411 26.07 3.486 ;
      RECT 26.05 2.394 26.055 2.72 ;
      RECT 26.045 2.775 26.055 3.543 ;
      RECT 26.04 2.38 26.05 2.693 ;
      RECT 26.035 2.83 26.045 3.825 ;
      RECT 26.03 2.366 26.04 2.678 ;
      RECT 26.03 2.88 26.035 3.825 ;
      RECT 26.015 2.343 26.03 2.658 ;
      RECT 25.995 3.002 26.03 3.825 ;
      RECT 26.01 2.325 26.015 2.64 ;
      RECT 26.005 2.317 26.01 2.63 ;
      RECT 25.975 2.285 26.005 2.594 ;
      RECT 25.985 3.13 25.995 3.825 ;
      RECT 25.98 3.157 25.985 3.825 ;
      RECT 25.975 3.207 25.98 3.825 ;
      RECT 25.965 2.251 25.975 2.559 ;
      RECT 25.925 3.275 25.975 3.825 ;
      RECT 25.95 2.228 25.965 2.535 ;
      RECT 25.925 2.1 25.95 2.498 ;
      RECT 25.92 2.1 25.925 2.47 ;
      RECT 25.89 3.375 25.925 3.825 ;
      RECT 25.915 2.1 25.92 2.463 ;
      RECT 25.91 2.1 25.915 2.453 ;
      RECT 25.895 2.1 25.91 2.438 ;
      RECT 25.88 2.1 25.895 2.41 ;
      RECT 25.845 3.48 25.89 3.825 ;
      RECT 25.865 2.1 25.88 2.383 ;
      RECT 25.835 2.1 25.865 2.368 ;
      RECT 25.83 3.552 25.845 3.825 ;
      RECT 25.755 2.635 25.795 2.895 ;
      RECT 25.53 2.582 25.535 2.84 ;
      RECT 21.485 2.06 21.745 2.32 ;
      RECT 21.485 2.085 21.76 2.3 ;
      RECT 23.875 1.91 23.88 2.055 ;
      RECT 25.745 2.63 25.755 2.895 ;
      RECT 25.725 2.622 25.745 2.895 ;
      RECT 25.707 2.618 25.725 2.895 ;
      RECT 25.621 2.607 25.707 2.895 ;
      RECT 25.535 2.59 25.621 2.895 ;
      RECT 25.48 2.577 25.53 2.825 ;
      RECT 25.446 2.569 25.48 2.8 ;
      RECT 25.36 2.558 25.446 2.765 ;
      RECT 25.325 2.535 25.36 2.73 ;
      RECT 25.315 2.497 25.325 2.716 ;
      RECT 25.31 2.47 25.315 2.712 ;
      RECT 25.305 2.457 25.31 2.709 ;
      RECT 25.295 2.437 25.305 2.705 ;
      RECT 25.29 2.412 25.295 2.701 ;
      RECT 25.265 2.367 25.29 2.695 ;
      RECT 25.255 2.308 25.265 2.687 ;
      RECT 25.245 2.276 25.255 2.678 ;
      RECT 25.225 2.228 25.245 2.658 ;
      RECT 25.22 2.188 25.225 2.628 ;
      RECT 25.205 2.162 25.22 2.602 ;
      RECT 25.2 2.14 25.205 2.578 ;
      RECT 25.185 2.112 25.2 2.554 ;
      RECT 25.17 2.085 25.185 2.518 ;
      RECT 25.155 2.062 25.17 2.48 ;
      RECT 25.15 2.052 25.155 2.455 ;
      RECT 25.14 2.045 25.15 2.438 ;
      RECT 25.125 2.032 25.14 2.408 ;
      RECT 25.12 2.022 25.125 2.383 ;
      RECT 25.115 2.017 25.12 2.37 ;
      RECT 25.105 2.01 25.115 2.35 ;
      RECT 25.1 2.003 25.105 2.335 ;
      RECT 25.075 1.996 25.1 2.293 ;
      RECT 25.06 1.986 25.075 2.243 ;
      RECT 25.05 1.981 25.06 2.213 ;
      RECT 25.04 1.977 25.05 2.188 ;
      RECT 25.025 1.974 25.04 2.178 ;
      RECT 24.975 1.971 25.025 2.163 ;
      RECT 24.955 1.969 24.975 2.148 ;
      RECT 24.906 1.967 24.955 2.143 ;
      RECT 24.82 1.963 24.906 2.138 ;
      RECT 24.781 1.96 24.82 2.134 ;
      RECT 24.695 1.956 24.781 2.129 ;
      RECT 24.645 1.953 24.695 2.123 ;
      RECT 24.596 1.95 24.645 2.118 ;
      RECT 24.51 1.947 24.596 2.113 ;
      RECT 24.506 1.945 24.51 2.11 ;
      RECT 24.42 1.942 24.506 2.105 ;
      RECT 24.371 1.938 24.42 2.098 ;
      RECT 24.285 1.935 24.371 2.093 ;
      RECT 24.261 1.932 24.285 2.089 ;
      RECT 24.175 1.93 24.261 2.084 ;
      RECT 24.11 1.926 24.175 2.077 ;
      RECT 24.107 1.925 24.11 2.074 ;
      RECT 24.021 1.922 24.107 2.071 ;
      RECT 23.935 1.916 24.021 2.064 ;
      RECT 23.905 1.912 23.935 2.06 ;
      RECT 23.88 1.91 23.905 2.058 ;
      RECT 23.825 1.907 23.875 2.055 ;
      RECT 23.745 1.906 23.825 2.055 ;
      RECT 23.69 1.908 23.745 2.058 ;
      RECT 23.675 1.909 23.69 2.062 ;
      RECT 23.62 1.917 23.675 2.072 ;
      RECT 23.59 1.925 23.62 2.085 ;
      RECT 23.571 1.926 23.59 2.091 ;
      RECT 23.485 1.929 23.571 2.096 ;
      RECT 23.415 1.934 23.485 2.105 ;
      RECT 23.396 1.937 23.415 2.111 ;
      RECT 23.31 1.941 23.396 2.116 ;
      RECT 23.27 1.945 23.31 2.123 ;
      RECT 23.261 1.947 23.27 2.126 ;
      RECT 23.175 1.951 23.261 2.131 ;
      RECT 23.172 1.954 23.175 2.135 ;
      RECT 23.086 1.957 23.172 2.139 ;
      RECT 23 1.963 23.086 2.147 ;
      RECT 22.976 1.967 23 2.151 ;
      RECT 22.89 1.971 22.976 2.156 ;
      RECT 22.845 1.976 22.89 2.163 ;
      RECT 22.765 1.981 22.845 2.17 ;
      RECT 22.685 1.987 22.765 2.185 ;
      RECT 22.66 1.991 22.685 2.198 ;
      RECT 22.595 1.994 22.66 2.21 ;
      RECT 22.54 1.999 22.595 2.225 ;
      RECT 22.51 2.002 22.54 2.243 ;
      RECT 22.5 2.004 22.51 2.256 ;
      RECT 22.44 2.019 22.5 2.266 ;
      RECT 22.425 2.036 22.44 2.275 ;
      RECT 22.42 2.045 22.425 2.275 ;
      RECT 22.41 2.055 22.42 2.275 ;
      RECT 22.4 2.072 22.41 2.275 ;
      RECT 22.38 2.082 22.4 2.276 ;
      RECT 22.335 2.092 22.38 2.277 ;
      RECT 22.3 2.101 22.335 2.279 ;
      RECT 22.235 2.106 22.3 2.281 ;
      RECT 22.155 2.107 22.235 2.284 ;
      RECT 22.151 2.105 22.155 2.285 ;
      RECT 22.065 2.102 22.151 2.287 ;
      RECT 22.018 2.099 22.065 2.289 ;
      RECT 21.932 2.095 22.018 2.292 ;
      RECT 21.846 2.091 21.932 2.295 ;
      RECT 21.76 2.087 21.846 2.299 ;
      RECT 23.695 3.15 23.975 3.43 ;
      RECT 23.735 3.13 23.995 3.39 ;
      RECT 23.725 3.14 23.995 3.39 ;
      RECT 23.735 3.067 23.95 3.43 ;
      RECT 23.79 2.99 23.945 3.43 ;
      RECT 23.795 2.775 23.945 3.43 ;
      RECT 23.785 2.577 23.935 2.828 ;
      RECT 23.775 2.577 23.935 2.695 ;
      RECT 23.77 2.455 23.93 2.598 ;
      RECT 23.755 2.455 23.93 2.503 ;
      RECT 23.75 2.165 23.925 2.48 ;
      RECT 23.735 2.165 23.925 2.45 ;
      RECT 23.695 2.165 23.955 2.425 ;
      RECT 23.605 3.635 23.685 3.895 ;
      RECT 23.01 2.355 23.015 2.62 ;
      RECT 22.89 2.355 23.015 2.615 ;
      RECT 23.565 3.6 23.605 3.895 ;
      RECT 23.52 3.522 23.565 3.895 ;
      RECT 23.5 3.45 23.52 3.895 ;
      RECT 23.49 3.402 23.5 3.895 ;
      RECT 23.455 3.335 23.49 3.895 ;
      RECT 23.425 3.235 23.455 3.895 ;
      RECT 23.405 3.16 23.425 3.695 ;
      RECT 23.395 3.11 23.405 3.65 ;
      RECT 23.39 3.087 23.395 3.623 ;
      RECT 23.385 3.072 23.39 3.61 ;
      RECT 23.38 3.057 23.385 3.588 ;
      RECT 23.375 3.042 23.38 3.57 ;
      RECT 23.35 2.997 23.375 3.525 ;
      RECT 23.34 2.945 23.35 3.468 ;
      RECT 23.33 2.915 23.34 3.435 ;
      RECT 23.32 2.88 23.33 3.403 ;
      RECT 23.285 2.812 23.32 3.335 ;
      RECT 23.28 2.751 23.285 3.27 ;
      RECT 23.27 2.739 23.28 3.25 ;
      RECT 23.265 2.727 23.27 3.23 ;
      RECT 23.26 2.719 23.265 3.218 ;
      RECT 23.255 2.711 23.26 3.198 ;
      RECT 23.245 2.699 23.255 3.17 ;
      RECT 23.235 2.683 23.245 3.14 ;
      RECT 23.21 2.655 23.235 3.078 ;
      RECT 23.2 2.626 23.21 3.023 ;
      RECT 23.185 2.605 23.2 2.983 ;
      RECT 23.18 2.589 23.185 2.955 ;
      RECT 23.175 2.577 23.18 2.945 ;
      RECT 23.17 2.572 23.175 2.918 ;
      RECT 23.165 2.565 23.17 2.905 ;
      RECT 23.15 2.548 23.165 2.878 ;
      RECT 23.14 2.355 23.15 2.838 ;
      RECT 23.13 2.355 23.14 2.805 ;
      RECT 23.12 2.355 23.13 2.78 ;
      RECT 23.05 2.355 23.12 2.715 ;
      RECT 23.04 2.355 23.05 2.663 ;
      RECT 23.025 2.355 23.04 2.645 ;
      RECT 23.015 2.355 23.025 2.63 ;
      RECT 22.845 3.225 23.105 3.485 ;
      RECT 21.38 3.26 21.385 3.467 ;
      RECT 21.015 3.15 21.09 3.465 ;
      RECT 20.83 3.205 20.985 3.465 ;
      RECT 21.015 3.15 21.12 3.43 ;
      RECT 22.83 3.322 22.845 3.483 ;
      RECT 22.805 3.33 22.83 3.488 ;
      RECT 22.78 3.337 22.805 3.493 ;
      RECT 22.717 3.348 22.78 3.502 ;
      RECT 22.631 3.367 22.717 3.519 ;
      RECT 22.545 3.389 22.631 3.538 ;
      RECT 22.53 3.402 22.545 3.549 ;
      RECT 22.49 3.41 22.53 3.556 ;
      RECT 22.47 3.415 22.49 3.563 ;
      RECT 22.432 3.416 22.47 3.566 ;
      RECT 22.346 3.419 22.432 3.567 ;
      RECT 22.26 3.423 22.346 3.568 ;
      RECT 22.211 3.425 22.26 3.57 ;
      RECT 22.125 3.425 22.211 3.572 ;
      RECT 22.085 3.42 22.125 3.574 ;
      RECT 22.075 3.414 22.085 3.575 ;
      RECT 22.035 3.409 22.075 3.572 ;
      RECT 22.025 3.402 22.035 3.568 ;
      RECT 22.01 3.398 22.025 3.566 ;
      RECT 21.993 3.394 22.01 3.564 ;
      RECT 21.907 3.384 21.993 3.556 ;
      RECT 21.821 3.366 21.907 3.542 ;
      RECT 21.735 3.349 21.821 3.528 ;
      RECT 21.71 3.337 21.735 3.519 ;
      RECT 21.64 3.327 21.71 3.512 ;
      RECT 21.595 3.315 21.64 3.503 ;
      RECT 21.535 3.302 21.595 3.495 ;
      RECT 21.53 3.294 21.535 3.49 ;
      RECT 21.495 3.289 21.53 3.488 ;
      RECT 21.44 3.28 21.495 3.481 ;
      RECT 21.4 3.269 21.44 3.473 ;
      RECT 21.385 3.262 21.4 3.469 ;
      RECT 21.365 3.255 21.38 3.466 ;
      RECT 21.35 3.245 21.365 3.464 ;
      RECT 21.335 3.232 21.35 3.461 ;
      RECT 21.31 3.215 21.335 3.457 ;
      RECT 21.295 3.197 21.31 3.454 ;
      RECT 21.27 3.15 21.295 3.452 ;
      RECT 21.246 3.15 21.27 3.449 ;
      RECT 21.16 3.15 21.246 3.441 ;
      RECT 21.12 3.15 21.16 3.433 ;
      RECT 20.985 3.197 21.015 3.465 ;
      RECT 22.665 2.78 22.925 3.04 ;
      RECT 22.625 2.78 22.925 2.918 ;
      RECT 22.59 2.78 22.925 2.903 ;
      RECT 22.535 2.78 22.925 2.883 ;
      RECT 22.455 2.59 22.735 2.87 ;
      RECT 22.455 2.772 22.805 2.87 ;
      RECT 22.455 2.715 22.79 2.87 ;
      RECT 22.455 2.662 22.74 2.87 ;
      RECT 19.615 2.949 19.63 3.405 ;
      RECT 19.61 3.021 19.716 3.403 ;
      RECT 19.63 2.115 19.765 3.401 ;
      RECT 19.615 2.965 19.77 3.4 ;
      RECT 19.615 3.015 19.775 3.398 ;
      RECT 19.6 3.08 19.775 3.397 ;
      RECT 19.61 3.072 19.78 3.394 ;
      RECT 19.59 3.12 19.78 3.389 ;
      RECT 19.59 3.12 19.795 3.386 ;
      RECT 19.585 3.12 19.795 3.383 ;
      RECT 19.56 3.12 19.82 3.38 ;
      RECT 19.63 2.115 19.79 2.768 ;
      RECT 19.625 2.115 19.79 2.74 ;
      RECT 19.62 2.115 19.79 2.568 ;
      RECT 19.62 2.115 19.81 2.508 ;
      RECT 19.575 2.115 19.835 2.375 ;
      RECT 19.055 2.59 19.335 2.87 ;
      RECT 19.045 2.605 19.335 2.865 ;
      RECT 19 2.667 19.335 2.863 ;
      RECT 19.075 2.582 19.24 2.87 ;
      RECT 19.075 2.567 19.196 2.87 ;
      RECT 19.11 2.56 19.196 2.87 ;
      RECT 18.575 3.71 18.855 3.99 ;
      RECT 18.535 3.672 18.83 3.783 ;
      RECT 18.52 3.622 18.81 3.678 ;
      RECT 18.465 3.385 18.725 3.645 ;
      RECT 18.465 3.587 18.805 3.645 ;
      RECT 18.465 3.527 18.8 3.645 ;
      RECT 18.465 3.477 18.78 3.645 ;
      RECT 18.465 3.457 18.775 3.645 ;
      RECT 18.465 3.435 18.77 3.645 ;
      RECT 18.465 3.42 18.74 3.645 ;
      RECT 15 6.655 15.325 6.98 ;
      RECT 13.885 6.745 15.325 6.915 ;
      RECT 13.885 2.395 14.045 6.915 ;
      RECT 14.2 2.365 14.52 2.685 ;
      RECT 13.885 2.395 14.52 2.565 ;
      RECT 13.145 5.84 13.495 6.19 ;
      RECT 13.22 2.705 13.395 6.19 ;
      RECT 13.155 2.705 13.505 3.055 ;
      RECT 7.17 4.36 12.84 4.53 ;
      RECT 12.67 3.425 12.84 4.53 ;
      RECT 7.225 3.71 7.255 3.99 ;
      RECT 6.975 3.6 6.995 3.99 ;
      RECT 6.93 3.6 6.995 3.86 ;
      RECT 12.58 3.43 12.93 3.78 ;
      RECT 6.76 2.225 6.795 2.485 ;
      RECT 6.535 2.225 6.595 2.485 ;
      RECT 7.215 3.69 7.225 3.99 ;
      RECT 7.21 3.65 7.215 3.99 ;
      RECT 7.195 3.605 7.21 3.99 ;
      RECT 7.19 3.57 7.195 3.99 ;
      RECT 7.185 3.55 7.19 3.99 ;
      RECT 7.17 3.508 7.185 3.99 ;
      RECT 7.155 3.446 7.17 4.53 ;
      RECT 7.135 3.375 7.155 4.53 ;
      RECT 7.125 3.305 7.135 4.53 ;
      RECT 7.08 3.245 7.125 4.53 ;
      RECT 7 3.207 7.08 4.53 ;
      RECT 6.995 3.198 7 3.99 ;
      RECT 6.99 3.197 6.995 3.57 ;
      RECT 6.98 3.196 6.99 3.553 ;
      RECT 6.955 3.177 6.98 3.523 ;
      RECT 6.95 3.152 6.955 3.502 ;
      RECT 6.94 3.13 6.95 3.493 ;
      RECT 6.935 3.101 6.94 3.483 ;
      RECT 6.895 3.027 6.935 3.455 ;
      RECT 6.875 2.928 6.895 3.42 ;
      RECT 6.86 2.864 6.875 3.403 ;
      RECT 6.83 2.788 6.86 3.375 ;
      RECT 6.81 2.703 6.83 3.348 ;
      RECT 6.77 2.599 6.81 3.255 ;
      RECT 6.765 2.52 6.77 3.163 ;
      RECT 6.76 2.503 6.765 3.14 ;
      RECT 6.755 2.225 6.76 3.12 ;
      RECT 6.725 2.225 6.755 3.058 ;
      RECT 6.72 2.225 6.725 2.99 ;
      RECT 6.71 2.225 6.72 2.955 ;
      RECT 6.7 2.225 6.71 2.92 ;
      RECT 6.635 2.225 6.7 2.775 ;
      RECT 6.63 2.225 6.635 2.645 ;
      RECT 6.6 2.225 6.63 2.578 ;
      RECT 6.595 2.225 6.6 2.503 ;
      RECT 10.93 2.16 11.19 2.42 ;
      RECT 10.925 2.16 11.19 2.368 ;
      RECT 10.92 2.16 11.19 2.338 ;
      RECT 10.895 2.03 11.175 2.31 ;
      RECT 9.935 3.71 10.215 3.99 ;
      RECT 9.975 3.665 10.24 3.925 ;
      RECT 9.965 3.7 10.24 3.925 ;
      RECT 9.97 3.685 10.215 3.99 ;
      RECT 9.975 3.662 10.185 3.99 ;
      RECT 9.975 3.66 10.17 3.99 ;
      RECT 10.015 3.65 10.17 3.99 ;
      RECT 9.985 3.655 10.17 3.99 ;
      RECT 10.015 3.647 10.115 3.99 ;
      RECT 10.04 3.64 10.115 3.99 ;
      RECT 10.02 3.642 10.115 3.99 ;
      RECT 9.35 3.155 9.61 3.415 ;
      RECT 9.4 3.147 9.59 3.415 ;
      RECT 9.405 3.067 9.59 3.415 ;
      RECT 9.525 2.455 9.59 3.415 ;
      RECT 9.43 2.852 9.59 3.415 ;
      RECT 9.505 2.54 9.59 3.415 ;
      RECT 9.54 2.165 9.676 2.893 ;
      RECT 9.485 2.662 9.676 2.893 ;
      RECT 9.5 2.602 9.59 3.415 ;
      RECT 9.54 2.165 9.7 2.558 ;
      RECT 9.54 2.165 9.71 2.455 ;
      RECT 9.53 2.165 9.79 2.425 ;
      RECT 8.935 3.71 9.215 3.99 ;
      RECT 8.955 3.67 9.215 3.99 ;
      RECT 8.595 3.625 8.7 3.885 ;
      RECT 8.45 2.115 8.54 2.375 ;
      RECT 8.99 3.18 8.995 3.22 ;
      RECT 8.985 3.17 8.99 3.305 ;
      RECT 8.98 3.16 8.985 3.398 ;
      RECT 8.97 3.14 8.98 3.454 ;
      RECT 8.89 3.068 8.97 3.534 ;
      RECT 8.925 3.712 8.935 3.937 ;
      RECT 8.92 3.709 8.925 3.932 ;
      RECT 8.905 3.706 8.92 3.925 ;
      RECT 8.87 3.7 8.905 3.907 ;
      RECT 8.885 3.003 8.89 3.608 ;
      RECT 8.865 2.954 8.885 3.623 ;
      RECT 8.855 3.687 8.87 3.89 ;
      RECT 8.86 2.896 8.865 3.638 ;
      RECT 8.855 2.874 8.86 3.648 ;
      RECT 8.82 2.784 8.855 3.885 ;
      RECT 8.805 2.662 8.82 3.885 ;
      RECT 8.8 2.615 8.805 3.885 ;
      RECT 8.775 2.54 8.8 3.885 ;
      RECT 8.76 2.455 8.775 3.885 ;
      RECT 8.755 2.402 8.76 3.885 ;
      RECT 8.75 2.382 8.755 3.885 ;
      RECT 8.745 2.357 8.75 3.119 ;
      RECT 8.73 3.317 8.75 3.885 ;
      RECT 8.74 2.335 8.745 3.096 ;
      RECT 8.73 2.287 8.74 3.061 ;
      RECT 8.725 2.25 8.73 3.027 ;
      RECT 8.725 3.397 8.73 3.885 ;
      RECT 8.71 2.227 8.725 2.982 ;
      RECT 8.705 3.495 8.725 3.885 ;
      RECT 8.655 2.115 8.71 2.824 ;
      RECT 8.7 3.617 8.705 3.885 ;
      RECT 8.64 2.115 8.655 2.663 ;
      RECT 8.635 2.115 8.64 2.615 ;
      RECT 8.63 2.115 8.635 2.603 ;
      RECT 8.585 2.115 8.63 2.54 ;
      RECT 8.56 2.115 8.585 2.458 ;
      RECT 8.545 2.115 8.56 2.41 ;
      RECT 8.54 2.115 8.545 2.38 ;
      RECT 7.865 3.565 7.91 3.825 ;
      RECT 7.77 2.1 7.915 2.36 ;
      RECT 8.275 2.722 8.285 2.813 ;
      RECT 8.26 2.66 8.275 2.869 ;
      RECT 8.255 2.607 8.26 2.915 ;
      RECT 8.205 2.554 8.255 3.041 ;
      RECT 8.2 2.509 8.205 3.188 ;
      RECT 8.19 2.497 8.2 3.23 ;
      RECT 8.155 2.461 8.19 3.335 ;
      RECT 8.15 2.429 8.155 3.441 ;
      RECT 8.135 2.411 8.15 3.486 ;
      RECT 8.13 2.394 8.135 2.72 ;
      RECT 8.125 2.775 8.135 3.543 ;
      RECT 8.12 2.38 8.13 2.693 ;
      RECT 8.115 2.83 8.125 3.825 ;
      RECT 8.11 2.366 8.12 2.678 ;
      RECT 8.11 2.88 8.115 3.825 ;
      RECT 8.095 2.343 8.11 2.658 ;
      RECT 8.075 3.002 8.11 3.825 ;
      RECT 8.09 2.325 8.095 2.64 ;
      RECT 8.085 2.317 8.09 2.63 ;
      RECT 8.055 2.285 8.085 2.594 ;
      RECT 8.065 3.13 8.075 3.825 ;
      RECT 8.06 3.157 8.065 3.825 ;
      RECT 8.055 3.207 8.06 3.825 ;
      RECT 8.045 2.251 8.055 2.559 ;
      RECT 8.005 3.275 8.055 3.825 ;
      RECT 8.03 2.228 8.045 2.535 ;
      RECT 8.005 2.1 8.03 2.498 ;
      RECT 8 2.1 8.005 2.47 ;
      RECT 7.97 3.375 8.005 3.825 ;
      RECT 7.995 2.1 8 2.463 ;
      RECT 7.99 2.1 7.995 2.453 ;
      RECT 7.975 2.1 7.99 2.438 ;
      RECT 7.96 2.1 7.975 2.41 ;
      RECT 7.925 3.48 7.97 3.825 ;
      RECT 7.945 2.1 7.96 2.383 ;
      RECT 7.915 2.1 7.945 2.368 ;
      RECT 7.91 3.552 7.925 3.825 ;
      RECT 7.835 2.635 7.875 2.895 ;
      RECT 7.61 2.582 7.615 2.84 ;
      RECT 3.565 2.06 3.825 2.32 ;
      RECT 3.565 2.085 3.84 2.3 ;
      RECT 5.955 1.91 5.96 2.055 ;
      RECT 7.825 2.63 7.835 2.895 ;
      RECT 7.805 2.622 7.825 2.895 ;
      RECT 7.787 2.618 7.805 2.895 ;
      RECT 7.701 2.607 7.787 2.895 ;
      RECT 7.615 2.59 7.701 2.895 ;
      RECT 7.56 2.577 7.61 2.825 ;
      RECT 7.526 2.569 7.56 2.8 ;
      RECT 7.44 2.558 7.526 2.765 ;
      RECT 7.405 2.535 7.44 2.73 ;
      RECT 7.395 2.497 7.405 2.716 ;
      RECT 7.39 2.47 7.395 2.712 ;
      RECT 7.385 2.457 7.39 2.709 ;
      RECT 7.375 2.437 7.385 2.705 ;
      RECT 7.37 2.412 7.375 2.701 ;
      RECT 7.345 2.367 7.37 2.695 ;
      RECT 7.335 2.308 7.345 2.687 ;
      RECT 7.325 2.276 7.335 2.678 ;
      RECT 7.305 2.228 7.325 2.658 ;
      RECT 7.3 2.188 7.305 2.628 ;
      RECT 7.285 2.162 7.3 2.602 ;
      RECT 7.28 2.14 7.285 2.578 ;
      RECT 7.265 2.112 7.28 2.554 ;
      RECT 7.25 2.085 7.265 2.518 ;
      RECT 7.235 2.062 7.25 2.48 ;
      RECT 7.23 2.052 7.235 2.455 ;
      RECT 7.22 2.045 7.23 2.438 ;
      RECT 7.205 2.032 7.22 2.408 ;
      RECT 7.2 2.022 7.205 2.383 ;
      RECT 7.195 2.017 7.2 2.37 ;
      RECT 7.185 2.01 7.195 2.35 ;
      RECT 7.18 2.003 7.185 2.335 ;
      RECT 7.155 1.996 7.18 2.293 ;
      RECT 7.14 1.986 7.155 2.243 ;
      RECT 7.13 1.981 7.14 2.213 ;
      RECT 7.12 1.977 7.13 2.188 ;
      RECT 7.105 1.974 7.12 2.178 ;
      RECT 7.055 1.971 7.105 2.163 ;
      RECT 7.035 1.969 7.055 2.148 ;
      RECT 6.986 1.967 7.035 2.143 ;
      RECT 6.9 1.963 6.986 2.138 ;
      RECT 6.861 1.96 6.9 2.134 ;
      RECT 6.775 1.956 6.861 2.129 ;
      RECT 6.725 1.953 6.775 2.123 ;
      RECT 6.676 1.95 6.725 2.118 ;
      RECT 6.59 1.947 6.676 2.113 ;
      RECT 6.586 1.945 6.59 2.11 ;
      RECT 6.5 1.942 6.586 2.105 ;
      RECT 6.451 1.938 6.5 2.098 ;
      RECT 6.365 1.935 6.451 2.093 ;
      RECT 6.341 1.932 6.365 2.089 ;
      RECT 6.255 1.93 6.341 2.084 ;
      RECT 6.19 1.926 6.255 2.077 ;
      RECT 6.187 1.925 6.19 2.074 ;
      RECT 6.101 1.922 6.187 2.071 ;
      RECT 6.015 1.916 6.101 2.064 ;
      RECT 5.985 1.912 6.015 2.06 ;
      RECT 5.96 1.91 5.985 2.058 ;
      RECT 5.905 1.907 5.955 2.055 ;
      RECT 5.825 1.906 5.905 2.055 ;
      RECT 5.77 1.908 5.825 2.058 ;
      RECT 5.755 1.909 5.77 2.062 ;
      RECT 5.7 1.917 5.755 2.072 ;
      RECT 5.67 1.925 5.7 2.085 ;
      RECT 5.651 1.926 5.67 2.091 ;
      RECT 5.565 1.929 5.651 2.096 ;
      RECT 5.495 1.934 5.565 2.105 ;
      RECT 5.476 1.937 5.495 2.111 ;
      RECT 5.39 1.941 5.476 2.116 ;
      RECT 5.35 1.945 5.39 2.123 ;
      RECT 5.341 1.947 5.35 2.126 ;
      RECT 5.255 1.951 5.341 2.131 ;
      RECT 5.252 1.954 5.255 2.135 ;
      RECT 5.166 1.957 5.252 2.139 ;
      RECT 5.08 1.963 5.166 2.147 ;
      RECT 5.056 1.967 5.08 2.151 ;
      RECT 4.97 1.971 5.056 2.156 ;
      RECT 4.925 1.976 4.97 2.163 ;
      RECT 4.845 1.981 4.925 2.17 ;
      RECT 4.765 1.987 4.845 2.185 ;
      RECT 4.74 1.991 4.765 2.198 ;
      RECT 4.675 1.994 4.74 2.21 ;
      RECT 4.62 1.999 4.675 2.225 ;
      RECT 4.59 2.002 4.62 2.243 ;
      RECT 4.58 2.004 4.59 2.256 ;
      RECT 4.52 2.019 4.58 2.266 ;
      RECT 4.505 2.036 4.52 2.275 ;
      RECT 4.5 2.045 4.505 2.275 ;
      RECT 4.49 2.055 4.5 2.275 ;
      RECT 4.48 2.072 4.49 2.275 ;
      RECT 4.46 2.082 4.48 2.276 ;
      RECT 4.415 2.092 4.46 2.277 ;
      RECT 4.38 2.101 4.415 2.279 ;
      RECT 4.315 2.106 4.38 2.281 ;
      RECT 4.235 2.107 4.315 2.284 ;
      RECT 4.231 2.105 4.235 2.285 ;
      RECT 4.145 2.102 4.231 2.287 ;
      RECT 4.098 2.099 4.145 2.289 ;
      RECT 4.012 2.095 4.098 2.292 ;
      RECT 3.926 2.091 4.012 2.295 ;
      RECT 3.84 2.087 3.926 2.299 ;
      RECT 5.775 3.15 6.055 3.43 ;
      RECT 5.815 3.13 6.075 3.39 ;
      RECT 5.805 3.14 6.075 3.39 ;
      RECT 5.815 3.067 6.03 3.43 ;
      RECT 5.87 2.99 6.025 3.43 ;
      RECT 5.875 2.775 6.025 3.43 ;
      RECT 5.865 2.577 6.015 2.828 ;
      RECT 5.855 2.577 6.015 2.695 ;
      RECT 5.85 2.455 6.01 2.598 ;
      RECT 5.835 2.455 6.01 2.503 ;
      RECT 5.83 2.165 6.005 2.48 ;
      RECT 5.815 2.165 6.005 2.45 ;
      RECT 5.775 2.165 6.035 2.425 ;
      RECT 5.685 3.635 5.765 3.895 ;
      RECT 5.09 2.355 5.095 2.62 ;
      RECT 4.97 2.355 5.095 2.615 ;
      RECT 5.645 3.6 5.685 3.895 ;
      RECT 5.6 3.522 5.645 3.895 ;
      RECT 5.58 3.45 5.6 3.895 ;
      RECT 5.57 3.402 5.58 3.895 ;
      RECT 5.535 3.335 5.57 3.895 ;
      RECT 5.505 3.235 5.535 3.895 ;
      RECT 5.485 3.16 5.505 3.695 ;
      RECT 5.475 3.11 5.485 3.65 ;
      RECT 5.47 3.087 5.475 3.623 ;
      RECT 5.465 3.072 5.47 3.61 ;
      RECT 5.46 3.057 5.465 3.588 ;
      RECT 5.455 3.042 5.46 3.57 ;
      RECT 5.43 2.997 5.455 3.525 ;
      RECT 5.42 2.945 5.43 3.468 ;
      RECT 5.41 2.915 5.42 3.435 ;
      RECT 5.4 2.88 5.41 3.403 ;
      RECT 5.365 2.812 5.4 3.335 ;
      RECT 5.36 2.751 5.365 3.27 ;
      RECT 5.35 2.739 5.36 3.25 ;
      RECT 5.345 2.727 5.35 3.23 ;
      RECT 5.34 2.719 5.345 3.218 ;
      RECT 5.335 2.711 5.34 3.198 ;
      RECT 5.325 2.699 5.335 3.17 ;
      RECT 5.315 2.683 5.325 3.14 ;
      RECT 5.29 2.655 5.315 3.078 ;
      RECT 5.28 2.626 5.29 3.023 ;
      RECT 5.265 2.605 5.28 2.983 ;
      RECT 5.26 2.589 5.265 2.955 ;
      RECT 5.255 2.577 5.26 2.945 ;
      RECT 5.25 2.572 5.255 2.918 ;
      RECT 5.245 2.565 5.25 2.905 ;
      RECT 5.23 2.548 5.245 2.878 ;
      RECT 5.22 2.355 5.23 2.838 ;
      RECT 5.21 2.355 5.22 2.805 ;
      RECT 5.2 2.355 5.21 2.78 ;
      RECT 5.13 2.355 5.2 2.715 ;
      RECT 5.12 2.355 5.13 2.663 ;
      RECT 5.105 2.355 5.12 2.645 ;
      RECT 5.095 2.355 5.105 2.63 ;
      RECT 4.925 3.225 5.185 3.485 ;
      RECT 3.46 3.26 3.465 3.467 ;
      RECT 3.095 3.15 3.17 3.465 ;
      RECT 2.91 3.205 3.065 3.465 ;
      RECT 3.095 3.15 3.2 3.43 ;
      RECT 4.91 3.322 4.925 3.483 ;
      RECT 4.885 3.33 4.91 3.488 ;
      RECT 4.86 3.337 4.885 3.493 ;
      RECT 4.797 3.348 4.86 3.502 ;
      RECT 4.711 3.367 4.797 3.519 ;
      RECT 4.625 3.389 4.711 3.538 ;
      RECT 4.61 3.402 4.625 3.549 ;
      RECT 4.57 3.41 4.61 3.556 ;
      RECT 4.55 3.415 4.57 3.563 ;
      RECT 4.512 3.416 4.55 3.566 ;
      RECT 4.426 3.419 4.512 3.567 ;
      RECT 4.34 3.423 4.426 3.568 ;
      RECT 4.291 3.425 4.34 3.57 ;
      RECT 4.205 3.425 4.291 3.572 ;
      RECT 4.165 3.42 4.205 3.574 ;
      RECT 4.155 3.414 4.165 3.575 ;
      RECT 4.115 3.409 4.155 3.572 ;
      RECT 4.105 3.402 4.115 3.568 ;
      RECT 4.09 3.398 4.105 3.566 ;
      RECT 4.073 3.394 4.09 3.564 ;
      RECT 3.987 3.384 4.073 3.556 ;
      RECT 3.901 3.366 3.987 3.542 ;
      RECT 3.815 3.349 3.901 3.528 ;
      RECT 3.79 3.337 3.815 3.519 ;
      RECT 3.72 3.327 3.79 3.512 ;
      RECT 3.675 3.315 3.72 3.503 ;
      RECT 3.615 3.302 3.675 3.495 ;
      RECT 3.61 3.294 3.615 3.49 ;
      RECT 3.575 3.289 3.61 3.488 ;
      RECT 3.52 3.28 3.575 3.481 ;
      RECT 3.48 3.269 3.52 3.473 ;
      RECT 3.465 3.262 3.48 3.469 ;
      RECT 3.445 3.255 3.46 3.466 ;
      RECT 3.43 3.245 3.445 3.464 ;
      RECT 3.415 3.232 3.43 3.461 ;
      RECT 3.39 3.215 3.415 3.457 ;
      RECT 3.375 3.197 3.39 3.454 ;
      RECT 3.35 3.15 3.375 3.452 ;
      RECT 3.326 3.15 3.35 3.449 ;
      RECT 3.24 3.15 3.326 3.441 ;
      RECT 3.2 3.15 3.24 3.433 ;
      RECT 3.065 3.197 3.095 3.465 ;
      RECT 4.745 2.78 5.005 3.04 ;
      RECT 4.705 2.78 5.005 2.918 ;
      RECT 4.67 2.78 5.005 2.903 ;
      RECT 4.615 2.78 5.005 2.883 ;
      RECT 4.535 2.59 4.815 2.87 ;
      RECT 4.535 2.772 4.885 2.87 ;
      RECT 4.535 2.715 4.87 2.87 ;
      RECT 4.535 2.662 4.82 2.87 ;
      RECT 1.695 2.949 1.71 3.405 ;
      RECT 1.69 3.021 1.796 3.403 ;
      RECT 1.71 2.115 1.845 3.401 ;
      RECT 1.695 2.965 1.85 3.4 ;
      RECT 1.695 3.015 1.855 3.398 ;
      RECT 1.68 3.08 1.855 3.397 ;
      RECT 1.69 3.072 1.86 3.394 ;
      RECT 1.67 3.12 1.86 3.389 ;
      RECT 1.67 3.12 1.875 3.386 ;
      RECT 1.665 3.12 1.875 3.383 ;
      RECT 1.64 3.12 1.9 3.38 ;
      RECT 1.71 2.115 1.87 2.768 ;
      RECT 1.705 2.115 1.87 2.74 ;
      RECT 1.7 2.115 1.87 2.568 ;
      RECT 1.7 2.115 1.89 2.508 ;
      RECT 1.655 2.115 1.915 2.375 ;
      RECT 1.135 2.59 1.415 2.87 ;
      RECT 1.125 2.605 1.415 2.865 ;
      RECT 1.08 2.667 1.415 2.863 ;
      RECT 1.155 2.582 1.32 2.87 ;
      RECT 1.155 2.567 1.276 2.87 ;
      RECT 1.19 2.56 1.276 2.87 ;
      RECT 0.655 3.71 0.935 3.99 ;
      RECT 0.615 3.672 0.91 3.783 ;
      RECT 0.6 3.622 0.89 3.678 ;
      RECT 0.545 3.385 0.805 3.645 ;
      RECT 0.545 3.587 0.885 3.645 ;
      RECT 0.545 3.527 0.88 3.645 ;
      RECT 0.545 3.477 0.86 3.645 ;
      RECT 0.545 3.457 0.855 3.645 ;
      RECT 0.545 3.435 0.85 3.645 ;
      RECT 0.545 3.42 0.82 3.645 ;
    LAYER via1 ;
      RECT 89.13 1.2 89.28 1.35 ;
      RECT 86.765 6.74 86.915 6.89 ;
      RECT 86.75 2.065 86.9 2.215 ;
      RECT 85.96 2.45 86.11 2.6 ;
      RECT 85.96 6.37 86.11 6.52 ;
      RECT 84.93 2.805 85.08 2.955 ;
      RECT 84.92 5.94 85.07 6.09 ;
      RECT 84.355 3.53 84.505 3.68 ;
      RECT 82.66 2.215 82.81 2.365 ;
      RECT 81.71 3.72 81.86 3.87 ;
      RECT 81.26 2.22 81.41 2.37 ;
      RECT 81.08 3.21 81.23 3.36 ;
      RECT 80.685 3.725 80.835 3.875 ;
      RECT 80.325 3.68 80.475 3.83 ;
      RECT 80.18 2.17 80.33 2.32 ;
      RECT 79.595 3.62 79.745 3.77 ;
      RECT 79.5 2.155 79.65 2.305 ;
      RECT 79.345 2.69 79.495 2.84 ;
      RECT 78.66 3.655 78.81 3.805 ;
      RECT 78.265 2.28 78.415 2.43 ;
      RECT 77.545 3.185 77.695 3.335 ;
      RECT 77.505 2.22 77.655 2.37 ;
      RECT 77.235 3.69 77.385 3.84 ;
      RECT 76.7 2.41 76.85 2.56 ;
      RECT 76.655 3.28 76.805 3.43 ;
      RECT 76.475 2.835 76.625 2.985 ;
      RECT 75.4 2.69 75.55 2.84 ;
      RECT 75.295 2.115 75.445 2.265 ;
      RECT 74.64 3.26 74.79 3.41 ;
      RECT 74.03 3.17 74.18 3.32 ;
      RECT 73.385 2.17 73.535 2.32 ;
      RECT 73.37 3.175 73.52 3.325 ;
      RECT 72.855 2.66 73.005 2.81 ;
      RECT 72.275 3.44 72.425 3.59 ;
      RECT 71.22 1.195 71.37 1.345 ;
      RECT 68.845 6.74 68.995 6.89 ;
      RECT 68.83 2.065 68.98 2.215 ;
      RECT 68.04 2.45 68.19 2.6 ;
      RECT 68.04 6.37 68.19 6.52 ;
      RECT 67.01 2.805 67.16 2.955 ;
      RECT 67 5.94 67.15 6.09 ;
      RECT 66.435 3.53 66.585 3.68 ;
      RECT 64.74 2.215 64.89 2.365 ;
      RECT 63.79 3.72 63.94 3.87 ;
      RECT 63.34 2.22 63.49 2.37 ;
      RECT 63.16 3.21 63.31 3.36 ;
      RECT 62.765 3.725 62.915 3.875 ;
      RECT 62.405 3.68 62.555 3.83 ;
      RECT 62.26 2.17 62.41 2.32 ;
      RECT 61.675 3.62 61.825 3.77 ;
      RECT 61.58 2.155 61.73 2.305 ;
      RECT 61.425 2.69 61.575 2.84 ;
      RECT 60.74 3.655 60.89 3.805 ;
      RECT 60.345 2.28 60.495 2.43 ;
      RECT 59.625 3.185 59.775 3.335 ;
      RECT 59.585 2.22 59.735 2.37 ;
      RECT 59.315 3.69 59.465 3.84 ;
      RECT 58.78 2.41 58.93 2.56 ;
      RECT 58.735 3.28 58.885 3.43 ;
      RECT 58.555 2.835 58.705 2.985 ;
      RECT 57.48 2.69 57.63 2.84 ;
      RECT 57.375 2.115 57.525 2.265 ;
      RECT 56.72 3.26 56.87 3.41 ;
      RECT 56.11 3.17 56.26 3.32 ;
      RECT 55.465 2.17 55.615 2.32 ;
      RECT 55.45 3.175 55.6 3.325 ;
      RECT 54.935 2.66 55.085 2.81 ;
      RECT 54.355 3.44 54.505 3.59 ;
      RECT 53.295 1.2 53.445 1.35 ;
      RECT 50.925 6.74 51.075 6.89 ;
      RECT 50.91 2.065 51.06 2.215 ;
      RECT 50.12 2.45 50.27 2.6 ;
      RECT 50.12 6.37 50.27 6.52 ;
      RECT 49.09 2.805 49.24 2.955 ;
      RECT 49.08 5.94 49.23 6.09 ;
      RECT 48.515 3.53 48.665 3.68 ;
      RECT 46.82 2.215 46.97 2.365 ;
      RECT 45.87 3.72 46.02 3.87 ;
      RECT 45.42 2.22 45.57 2.37 ;
      RECT 45.24 3.21 45.39 3.36 ;
      RECT 44.845 3.725 44.995 3.875 ;
      RECT 44.485 3.68 44.635 3.83 ;
      RECT 44.34 2.17 44.49 2.32 ;
      RECT 43.755 3.62 43.905 3.77 ;
      RECT 43.66 2.155 43.81 2.305 ;
      RECT 43.505 2.69 43.655 2.84 ;
      RECT 42.82 3.655 42.97 3.805 ;
      RECT 42.425 2.28 42.575 2.43 ;
      RECT 41.705 3.185 41.855 3.335 ;
      RECT 41.665 2.22 41.815 2.37 ;
      RECT 41.395 3.69 41.545 3.84 ;
      RECT 40.86 2.41 41.01 2.56 ;
      RECT 40.815 3.28 40.965 3.43 ;
      RECT 40.635 2.835 40.785 2.985 ;
      RECT 39.56 2.69 39.71 2.84 ;
      RECT 39.455 2.115 39.605 2.265 ;
      RECT 38.8 3.26 38.95 3.41 ;
      RECT 38.19 3.17 38.34 3.32 ;
      RECT 37.545 2.17 37.695 2.32 ;
      RECT 37.53 3.175 37.68 3.325 ;
      RECT 37.015 2.66 37.165 2.81 ;
      RECT 36.435 3.44 36.585 3.59 ;
      RECT 35.375 1.195 35.525 1.345 ;
      RECT 33.01 6.74 33.16 6.89 ;
      RECT 32.995 2.065 33.145 2.215 ;
      RECT 32.205 2.45 32.355 2.6 ;
      RECT 32.205 6.37 32.355 6.52 ;
      RECT 31.175 2.805 31.325 2.955 ;
      RECT 31.165 5.94 31.315 6.09 ;
      RECT 30.6 3.53 30.75 3.68 ;
      RECT 28.905 2.215 29.055 2.365 ;
      RECT 27.955 3.72 28.105 3.87 ;
      RECT 27.505 2.22 27.655 2.37 ;
      RECT 27.325 3.21 27.475 3.36 ;
      RECT 26.93 3.725 27.08 3.875 ;
      RECT 26.57 3.68 26.72 3.83 ;
      RECT 26.425 2.17 26.575 2.32 ;
      RECT 25.84 3.62 25.99 3.77 ;
      RECT 25.745 2.155 25.895 2.305 ;
      RECT 25.59 2.69 25.74 2.84 ;
      RECT 24.905 3.655 25.055 3.805 ;
      RECT 24.51 2.28 24.66 2.43 ;
      RECT 23.79 3.185 23.94 3.335 ;
      RECT 23.75 2.22 23.9 2.37 ;
      RECT 23.48 3.69 23.63 3.84 ;
      RECT 22.945 2.41 23.095 2.56 ;
      RECT 22.9 3.28 23.05 3.43 ;
      RECT 22.72 2.835 22.87 2.985 ;
      RECT 21.645 2.69 21.795 2.84 ;
      RECT 21.54 2.115 21.69 2.265 ;
      RECT 20.885 3.26 21.035 3.41 ;
      RECT 20.275 3.17 20.425 3.32 ;
      RECT 19.63 2.17 19.78 2.32 ;
      RECT 19.615 3.175 19.765 3.325 ;
      RECT 19.1 2.66 19.25 2.81 ;
      RECT 18.52 3.44 18.67 3.59 ;
      RECT 17.405 1.195 17.555 1.345 ;
      RECT 15.09 6.74 15.24 6.89 ;
      RECT 15.075 2.065 15.225 2.215 ;
      RECT 14.285 2.45 14.435 2.6 ;
      RECT 14.285 6.37 14.435 6.52 ;
      RECT 13.255 2.805 13.405 2.955 ;
      RECT 13.245 5.94 13.395 6.09 ;
      RECT 12.68 3.53 12.83 3.68 ;
      RECT 10.985 2.215 11.135 2.365 ;
      RECT 10.035 3.72 10.185 3.87 ;
      RECT 9.585 2.22 9.735 2.37 ;
      RECT 9.405 3.21 9.555 3.36 ;
      RECT 9.01 3.725 9.16 3.875 ;
      RECT 8.65 3.68 8.8 3.83 ;
      RECT 8.505 2.17 8.655 2.32 ;
      RECT 7.92 3.62 8.07 3.77 ;
      RECT 7.825 2.155 7.975 2.305 ;
      RECT 7.67 2.69 7.82 2.84 ;
      RECT 6.985 3.655 7.135 3.805 ;
      RECT 6.59 2.28 6.74 2.43 ;
      RECT 5.87 3.185 6.02 3.335 ;
      RECT 5.83 2.22 5.98 2.37 ;
      RECT 5.56 3.69 5.71 3.84 ;
      RECT 5.025 2.41 5.175 2.56 ;
      RECT 4.98 3.28 5.13 3.43 ;
      RECT 4.8 2.835 4.95 2.985 ;
      RECT 3.725 2.69 3.875 2.84 ;
      RECT 3.62 2.115 3.77 2.265 ;
      RECT 2.965 3.26 3.115 3.41 ;
      RECT 2.355 3.17 2.505 3.32 ;
      RECT 1.71 2.17 1.86 2.32 ;
      RECT 1.695 3.175 1.845 3.325 ;
      RECT 1.18 2.66 1.33 2.81 ;
      RECT 0.6 3.44 0.75 3.59 ;
    LAYER met1 ;
      RECT 72.055 0 84.015 1.89 ;
      RECT 54.135 0 66.095 1.89 ;
      RECT 36.215 0 48.175 1.89 ;
      RECT 18.3 0 30.26 1.89 ;
      RECT 0.38 0 12.34 1.89 ;
      RECT 72.05 0 84.015 1.68 ;
      RECT 54.13 0 66.095 1.68 ;
      RECT 36.21 0 48.175 1.68 ;
      RECT 18.295 0 30.26 1.68 ;
      RECT 0.375 0 12.34 1.68 ;
      RECT 0.005 0 89.605 0.305 ;
      RECT 0.005 4.285 89.605 4.745 ;
      RECT 72.055 4.135 89.605 4.745 ;
      RECT 54.135 4.135 71.685 4.745 ;
      RECT 36.215 4.135 53.765 4.745 ;
      RECT 18.3 4.135 35.85 4.745 ;
      RECT 0.38 4.135 17.93 4.745 ;
      RECT 72.055 4.13 84.015 4.745 ;
      RECT 54.135 4.13 66.095 4.745 ;
      RECT 36.215 4.13 48.175 4.745 ;
      RECT 18.3 4.13 30.26 4.745 ;
      RECT 0.38 4.13 12.34 4.745 ;
      RECT 89.005 2.365 89.295 2.595 ;
      RECT 89.065 0.885 89.235 2.595 ;
      RECT 89.03 1.1 89.38 1.45 ;
      RECT 89.005 0.885 89.295 1.115 ;
      RECT 89.005 7.765 89.295 7.995 ;
      RECT 89.065 6.285 89.235 7.995 ;
      RECT 89.005 6.285 89.295 6.515 ;
      RECT 88.595 2.735 88.925 2.965 ;
      RECT 88.595 2.765 89.095 2.935 ;
      RECT 88.595 2.395 88.785 2.965 ;
      RECT 88.015 2.365 88.305 2.595 ;
      RECT 88.015 2.395 88.785 2.565 ;
      RECT 88.075 0.885 88.245 2.595 ;
      RECT 88.015 0.885 88.305 1.115 ;
      RECT 88.015 7.765 88.305 7.995 ;
      RECT 88.075 6.285 88.245 7.995 ;
      RECT 88.015 6.285 88.305 6.515 ;
      RECT 88.015 6.325 88.865 6.485 ;
      RECT 88.695 5.915 88.865 6.485 ;
      RECT 88.015 6.32 88.405 6.485 ;
      RECT 88.635 5.915 88.925 6.145 ;
      RECT 88.635 5.945 89.095 6.115 ;
      RECT 87.645 2.735 87.935 2.965 ;
      RECT 87.645 2.765 88.105 2.935 ;
      RECT 87.705 1.655 87.87 2.965 ;
      RECT 86.22 1.625 86.51 1.855 ;
      RECT 86.22 1.655 87.87 1.825 ;
      RECT 86.28 0.885 86.45 1.855 ;
      RECT 86.22 0.885 86.51 1.115 ;
      RECT 86.22 7.765 86.51 7.995 ;
      RECT 86.28 7.025 86.45 7.995 ;
      RECT 86.28 7.12 87.87 7.29 ;
      RECT 87.7 5.915 87.87 7.29 ;
      RECT 86.22 7.025 86.51 7.255 ;
      RECT 87.645 5.915 87.935 6.145 ;
      RECT 87.645 5.945 88.105 6.115 ;
      RECT 86.65 1.965 87 2.315 ;
      RECT 86.48 2.025 87 2.195 ;
      RECT 86.675 6.655 87 6.98 ;
      RECT 86.65 6.655 87 6.885 ;
      RECT 86.48 6.685 87 6.855 ;
      RECT 84.255 3.43 84.605 3.78 ;
      RECT 84.345 2.395 84.515 3.78 ;
      RECT 85.875 2.365 86.195 2.685 ;
      RECT 85.845 2.365 86.195 2.595 ;
      RECT 84.345 2.395 86.195 2.565 ;
      RECT 85.875 6.28 86.195 6.605 ;
      RECT 85.845 6.285 86.195 6.515 ;
      RECT 85.675 6.315 86.195 6.485 ;
      RECT 84.83 2.705 85.18 3.055 ;
      RECT 84.83 2.765 85.31 2.935 ;
      RECT 84.82 5.84 85.17 6.19 ;
      RECT 84.82 5.945 85.31 6.115 ;
      RECT 81.655 3.665 81.695 3.925 ;
      RECT 81.695 3.645 81.7 3.655 ;
      RECT 83.035 2.735 83.19 3.055 ;
      RECT 82.955 2.735 83.035 3.22 ;
      RECT 82.945 2.735 82.955 3.363 ;
      RECT 82.92 2.735 82.945 3.41 ;
      RECT 82.895 2.735 82.92 3.488 ;
      RECT 82.875 2.735 82.895 3.558 ;
      RECT 82.87 2.735 82.875 3.588 ;
      RECT 82.85 2.885 82.87 3.6 ;
      RECT 82.84 2.885 82.85 3.618 ;
      RECT 82.83 2.887 82.84 3.626 ;
      RECT 82.825 2.892 82.83 3.083 ;
      RECT 82.825 3.092 82.83 3.627 ;
      RECT 82.82 3.137 82.825 3.628 ;
      RECT 82.81 3.202 82.82 3.629 ;
      RECT 82.8 3.297 82.81 3.631 ;
      RECT 82.795 3.35 82.8 3.633 ;
      RECT 82.79 3.37 82.795 3.634 ;
      RECT 82.735 3.395 82.79 3.64 ;
      RECT 82.695 3.43 82.735 3.649 ;
      RECT 82.685 3.447 82.695 3.654 ;
      RECT 82.676 3.453 82.685 3.656 ;
      RECT 82.59 3.491 82.676 3.667 ;
      RECT 82.585 3.53 82.59 3.677 ;
      RECT 82.51 3.537 82.585 3.687 ;
      RECT 82.49 3.547 82.51 3.698 ;
      RECT 82.46 3.554 82.49 3.706 ;
      RECT 82.435 3.561 82.46 3.713 ;
      RECT 82.411 3.567 82.435 3.718 ;
      RECT 82.325 3.58 82.411 3.73 ;
      RECT 82.247 3.587 82.325 3.748 ;
      RECT 82.161 3.582 82.247 3.766 ;
      RECT 82.075 3.577 82.161 3.786 ;
      RECT 81.995 3.571 82.075 3.803 ;
      RECT 81.93 3.567 81.995 3.832 ;
      RECT 81.925 3.281 81.93 3.305 ;
      RECT 81.915 3.557 81.93 3.86 ;
      RECT 81.92 3.275 81.925 3.345 ;
      RECT 81.915 3.269 81.92 3.415 ;
      RECT 81.91 3.263 81.915 3.493 ;
      RECT 81.91 3.54 81.915 3.925 ;
      RECT 81.902 3.26 81.91 3.925 ;
      RECT 81.816 3.258 81.902 3.925 ;
      RECT 81.73 3.256 81.816 3.925 ;
      RECT 81.72 3.257 81.73 3.925 ;
      RECT 81.715 3.262 81.72 3.925 ;
      RECT 81.705 3.275 81.715 3.925 ;
      RECT 81.7 3.297 81.705 3.925 ;
      RECT 81.695 3.657 81.7 3.925 ;
      RECT 82.325 3.125 82.33 3.345 ;
      RECT 82.83 2.16 82.865 2.42 ;
      RECT 82.815 2.16 82.83 2.428 ;
      RECT 82.786 2.16 82.815 2.45 ;
      RECT 82.7 2.16 82.786 2.51 ;
      RECT 82.68 2.16 82.7 2.575 ;
      RECT 82.62 2.16 82.68 2.74 ;
      RECT 82.615 2.16 82.62 2.888 ;
      RECT 82.61 2.16 82.615 2.9 ;
      RECT 82.605 2.16 82.61 2.926 ;
      RECT 82.575 2.346 82.605 3.006 ;
      RECT 82.57 2.394 82.575 3.095 ;
      RECT 82.565 2.408 82.57 3.11 ;
      RECT 82.56 2.427 82.565 3.14 ;
      RECT 82.555 2.442 82.56 3.156 ;
      RECT 82.55 2.457 82.555 3.178 ;
      RECT 82.545 2.477 82.55 3.2 ;
      RECT 82.535 2.497 82.545 3.233 ;
      RECT 82.52 2.539 82.535 3.295 ;
      RECT 82.515 2.57 82.52 3.335 ;
      RECT 82.51 2.582 82.515 3.34 ;
      RECT 82.505 2.594 82.51 3.345 ;
      RECT 82.5 2.607 82.505 3.345 ;
      RECT 82.495 2.625 82.5 3.345 ;
      RECT 82.49 2.645 82.495 3.345 ;
      RECT 82.485 2.657 82.49 3.345 ;
      RECT 82.48 2.67 82.485 3.345 ;
      RECT 82.46 2.705 82.48 3.345 ;
      RECT 82.41 2.807 82.46 3.345 ;
      RECT 82.405 2.892 82.41 3.345 ;
      RECT 82.4 2.9 82.405 3.345 ;
      RECT 82.395 2.917 82.4 3.345 ;
      RECT 82.39 2.932 82.395 3.345 ;
      RECT 82.355 2.997 82.39 3.345 ;
      RECT 82.34 3.062 82.355 3.345 ;
      RECT 82.335 3.092 82.34 3.345 ;
      RECT 82.33 3.117 82.335 3.345 ;
      RECT 82.315 3.127 82.325 3.345 ;
      RECT 82.3 3.14 82.315 3.338 ;
      RECT 82.045 2.73 82.115 2.94 ;
      RECT 81.835 2.707 81.84 2.9 ;
      RECT 79.29 2.635 79.55 2.895 ;
      RECT 82.125 2.917 82.13 2.92 ;
      RECT 82.115 2.735 82.125 2.935 ;
      RECT 82.016 2.728 82.045 2.94 ;
      RECT 81.93 2.72 82.016 2.94 ;
      RECT 81.915 2.714 81.93 2.938 ;
      RECT 81.895 2.713 81.915 2.925 ;
      RECT 81.89 2.712 81.895 2.908 ;
      RECT 81.84 2.709 81.89 2.903 ;
      RECT 81.81 2.706 81.835 2.898 ;
      RECT 81.79 2.704 81.81 2.893 ;
      RECT 81.775 2.702 81.79 2.89 ;
      RECT 81.745 2.7 81.775 2.888 ;
      RECT 81.68 2.696 81.745 2.88 ;
      RECT 81.65 2.691 81.68 2.875 ;
      RECT 81.63 2.689 81.65 2.873 ;
      RECT 81.6 2.686 81.63 2.868 ;
      RECT 81.54 2.682 81.6 2.86 ;
      RECT 81.535 2.679 81.54 2.855 ;
      RECT 81.465 2.677 81.535 2.85 ;
      RECT 81.436 2.673 81.465 2.843 ;
      RECT 81.35 2.668 81.436 2.835 ;
      RECT 81.316 2.663 81.35 2.827 ;
      RECT 81.23 2.655 81.316 2.819 ;
      RECT 81.191 2.648 81.23 2.811 ;
      RECT 81.105 2.643 81.191 2.803 ;
      RECT 81.04 2.637 81.105 2.793 ;
      RECT 81.02 2.632 81.04 2.788 ;
      RECT 81.011 2.629 81.02 2.787 ;
      RECT 80.925 2.625 81.011 2.781 ;
      RECT 80.885 2.621 80.925 2.773 ;
      RECT 80.865 2.617 80.885 2.771 ;
      RECT 80.805 2.617 80.865 2.768 ;
      RECT 80.785 2.62 80.805 2.766 ;
      RECT 80.764 2.62 80.785 2.766 ;
      RECT 80.678 2.622 80.764 2.77 ;
      RECT 80.592 2.624 80.678 2.776 ;
      RECT 80.506 2.626 80.592 2.783 ;
      RECT 80.42 2.629 80.506 2.789 ;
      RECT 80.386 2.63 80.42 2.794 ;
      RECT 80.3 2.633 80.386 2.799 ;
      RECT 80.271 2.64 80.3 2.804 ;
      RECT 80.185 2.64 80.271 2.809 ;
      RECT 80.152 2.64 80.185 2.814 ;
      RECT 80.066 2.642 80.152 2.819 ;
      RECT 79.98 2.644 80.066 2.826 ;
      RECT 79.916 2.646 79.98 2.832 ;
      RECT 79.83 2.648 79.916 2.838 ;
      RECT 79.827 2.65 79.83 2.841 ;
      RECT 79.741 2.651 79.827 2.845 ;
      RECT 79.655 2.654 79.741 2.852 ;
      RECT 79.636 2.656 79.655 2.856 ;
      RECT 79.55 2.658 79.636 2.861 ;
      RECT 79.28 2.67 79.29 2.865 ;
      RECT 81.515 2.25 81.7 2.46 ;
      RECT 81.51 2.251 81.705 2.458 ;
      RECT 81.505 2.256 81.715 2.453 ;
      RECT 81.5 2.232 81.505 2.45 ;
      RECT 81.47 2.229 81.5 2.443 ;
      RECT 81.465 2.225 81.47 2.434 ;
      RECT 81.43 2.256 81.715 2.429 ;
      RECT 81.205 2.165 81.465 2.425 ;
      RECT 81.505 2.234 81.51 2.453 ;
      RECT 81.51 2.235 81.515 2.458 ;
      RECT 81.205 2.247 81.585 2.425 ;
      RECT 81.205 2.245 81.57 2.425 ;
      RECT 81.205 2.24 81.56 2.425 ;
      RECT 81.16 3.155 81.21 3.44 ;
      RECT 81.105 3.125 81.11 3.44 ;
      RECT 81.075 3.105 81.08 3.44 ;
      RECT 81.225 3.155 81.285 3.415 ;
      RECT 81.22 3.155 81.225 3.423 ;
      RECT 81.21 3.155 81.22 3.435 ;
      RECT 81.125 3.145 81.16 3.44 ;
      RECT 81.12 3.132 81.125 3.44 ;
      RECT 81.11 3.127 81.12 3.44 ;
      RECT 81.09 3.117 81.105 3.44 ;
      RECT 81.08 3.11 81.09 3.44 ;
      RECT 81.07 3.102 81.075 3.44 ;
      RECT 81.04 3.092 81.07 3.44 ;
      RECT 81.025 3.08 81.04 3.44 ;
      RECT 81.01 3.07 81.025 3.435 ;
      RECT 80.99 3.06 81.01 3.41 ;
      RECT 80.98 3.052 80.99 3.387 ;
      RECT 80.95 3.035 80.98 3.377 ;
      RECT 80.945 3.012 80.95 3.368 ;
      RECT 80.94 2.999 80.945 3.366 ;
      RECT 80.925 2.975 80.94 3.36 ;
      RECT 80.92 2.951 80.925 3.354 ;
      RECT 80.91 2.94 80.92 3.349 ;
      RECT 80.905 2.93 80.91 3.345 ;
      RECT 80.9 2.922 80.905 3.342 ;
      RECT 80.89 2.917 80.9 3.338 ;
      RECT 80.885 2.912 80.89 3.334 ;
      RECT 80.8 2.91 80.885 3.309 ;
      RECT 80.77 2.91 80.8 3.275 ;
      RECT 80.755 2.91 80.77 3.258 ;
      RECT 80.7 2.91 80.755 3.203 ;
      RECT 80.695 2.915 80.7 3.152 ;
      RECT 80.685 2.92 80.695 3.142 ;
      RECT 80.68 2.93 80.685 3.128 ;
      RECT 80.63 3.67 80.89 3.93 ;
      RECT 80.55 3.685 80.89 3.906 ;
      RECT 80.53 3.685 80.89 3.901 ;
      RECT 80.506 3.685 80.89 3.899 ;
      RECT 80.42 3.685 80.89 3.894 ;
      RECT 80.27 3.625 80.53 3.89 ;
      RECT 80.225 3.685 80.89 3.885 ;
      RECT 80.22 3.692 80.89 3.88 ;
      RECT 80.235 3.68 80.55 3.89 ;
      RECT 80.125 2.115 80.385 2.375 ;
      RECT 80.125 2.172 80.39 2.368 ;
      RECT 80.125 2.202 80.395 2.3 ;
      RECT 80.185 2.633 80.3 2.635 ;
      RECT 80.271 2.63 80.3 2.635 ;
      RECT 79.295 3.634 79.32 3.874 ;
      RECT 79.28 3.637 79.37 3.868 ;
      RECT 79.275 3.642 79.456 3.863 ;
      RECT 79.27 3.65 79.52 3.861 ;
      RECT 79.27 3.65 79.53 3.86 ;
      RECT 79.265 3.657 79.54 3.853 ;
      RECT 79.265 3.657 79.626 3.842 ;
      RECT 79.26 3.692 79.626 3.838 ;
      RECT 79.26 3.692 79.635 3.827 ;
      RECT 79.54 3.565 79.8 3.825 ;
      RECT 79.25 3.742 79.8 3.823 ;
      RECT 79.52 3.61 79.54 3.858 ;
      RECT 79.456 3.613 79.52 3.862 ;
      RECT 79.37 3.618 79.456 3.867 ;
      RECT 79.3 3.629 79.8 3.825 ;
      RECT 79.32 3.623 79.37 3.872 ;
      RECT 79.445 2.1 79.455 2.362 ;
      RECT 79.435 2.157 79.445 2.365 ;
      RECT 79.41 2.162 79.435 2.371 ;
      RECT 79.385 2.166 79.41 2.383 ;
      RECT 79.375 2.169 79.385 2.393 ;
      RECT 79.37 2.17 79.375 2.398 ;
      RECT 79.365 2.171 79.37 2.403 ;
      RECT 79.36 2.172 79.365 2.405 ;
      RECT 79.335 2.175 79.36 2.408 ;
      RECT 79.305 2.181 79.335 2.411 ;
      RECT 79.24 2.192 79.305 2.414 ;
      RECT 79.195 2.2 79.24 2.418 ;
      RECT 79.18 2.2 79.195 2.426 ;
      RECT 79.175 2.201 79.18 2.433 ;
      RECT 79.17 2.203 79.175 2.436 ;
      RECT 79.165 2.207 79.17 2.439 ;
      RECT 79.155 2.215 79.165 2.443 ;
      RECT 79.15 2.228 79.155 2.448 ;
      RECT 79.145 2.236 79.15 2.45 ;
      RECT 79.14 2.242 79.145 2.45 ;
      RECT 79.135 2.246 79.14 2.453 ;
      RECT 79.13 2.248 79.135 2.456 ;
      RECT 79.125 2.251 79.13 2.459 ;
      RECT 79.115 2.256 79.125 2.463 ;
      RECT 79.11 2.262 79.115 2.468 ;
      RECT 79.1 2.268 79.11 2.472 ;
      RECT 79.085 2.275 79.1 2.478 ;
      RECT 79.056 2.289 79.085 2.488 ;
      RECT 78.97 2.324 79.056 2.52 ;
      RECT 78.95 2.357 78.97 2.549 ;
      RECT 78.93 2.37 78.95 2.56 ;
      RECT 78.91 2.382 78.93 2.571 ;
      RECT 78.86 2.404 78.91 2.591 ;
      RECT 78.845 2.422 78.86 2.608 ;
      RECT 78.84 2.428 78.845 2.611 ;
      RECT 78.835 2.432 78.84 2.614 ;
      RECT 78.83 2.436 78.835 2.618 ;
      RECT 78.825 2.438 78.83 2.621 ;
      RECT 78.815 2.445 78.825 2.624 ;
      RECT 78.81 2.45 78.815 2.628 ;
      RECT 78.805 2.452 78.81 2.631 ;
      RECT 78.8 2.456 78.805 2.634 ;
      RECT 78.795 2.458 78.8 2.638 ;
      RECT 78.78 2.463 78.795 2.643 ;
      RECT 78.775 2.468 78.78 2.646 ;
      RECT 78.77 2.476 78.775 2.649 ;
      RECT 78.765 2.478 78.77 2.652 ;
      RECT 78.76 2.48 78.765 2.655 ;
      RECT 78.75 2.482 78.76 2.661 ;
      RECT 78.715 2.496 78.75 2.673 ;
      RECT 78.705 2.511 78.715 2.683 ;
      RECT 78.63 2.54 78.705 2.707 ;
      RECT 78.625 2.565 78.63 2.73 ;
      RECT 78.61 2.569 78.625 2.736 ;
      RECT 78.6 2.577 78.61 2.741 ;
      RECT 78.57 2.59 78.6 2.745 ;
      RECT 78.56 2.605 78.57 2.75 ;
      RECT 78.55 2.61 78.56 2.753 ;
      RECT 78.545 2.612 78.55 2.755 ;
      RECT 78.53 2.615 78.545 2.758 ;
      RECT 78.525 2.617 78.53 2.761 ;
      RECT 78.505 2.622 78.525 2.765 ;
      RECT 78.475 2.627 78.505 2.773 ;
      RECT 78.45 2.634 78.475 2.781 ;
      RECT 78.445 2.639 78.45 2.786 ;
      RECT 78.415 2.642 78.445 2.79 ;
      RECT 78.375 2.645 78.415 2.8 ;
      RECT 78.34 2.642 78.375 2.812 ;
      RECT 78.33 2.638 78.34 2.819 ;
      RECT 78.305 2.634 78.33 2.825 ;
      RECT 78.3 2.63 78.305 2.83 ;
      RECT 78.26 2.627 78.3 2.83 ;
      RECT 78.245 2.612 78.26 2.831 ;
      RECT 78.222 2.6 78.245 2.831 ;
      RECT 78.136 2.6 78.222 2.832 ;
      RECT 78.05 2.6 78.136 2.834 ;
      RECT 78.03 2.6 78.05 2.831 ;
      RECT 78.025 2.605 78.03 2.826 ;
      RECT 78.02 2.61 78.025 2.824 ;
      RECT 78.01 2.62 78.02 2.822 ;
      RECT 78.005 2.626 78.01 2.815 ;
      RECT 78 2.628 78.005 2.8 ;
      RECT 77.995 2.632 78 2.79 ;
      RECT 79.455 2.1 79.705 2.36 ;
      RECT 77.18 3.635 77.44 3.895 ;
      RECT 79.475 3.125 79.48 3.335 ;
      RECT 79.48 3.13 79.49 3.33 ;
      RECT 79.43 3.125 79.475 3.35 ;
      RECT 79.42 3.125 79.43 3.37 ;
      RECT 79.401 3.125 79.42 3.375 ;
      RECT 79.315 3.125 79.401 3.372 ;
      RECT 79.285 3.127 79.315 3.37 ;
      RECT 79.23 3.137 79.285 3.368 ;
      RECT 79.165 3.151 79.23 3.366 ;
      RECT 79.16 3.159 79.165 3.365 ;
      RECT 79.145 3.162 79.16 3.363 ;
      RECT 79.08 3.172 79.145 3.359 ;
      RECT 79.032 3.186 79.08 3.36 ;
      RECT 78.946 3.203 79.032 3.374 ;
      RECT 78.86 3.224 78.946 3.391 ;
      RECT 78.84 3.237 78.86 3.401 ;
      RECT 78.795 3.245 78.84 3.408 ;
      RECT 78.76 3.253 78.795 3.416 ;
      RECT 78.726 3.261 78.76 3.424 ;
      RECT 78.64 3.275 78.726 3.436 ;
      RECT 78.605 3.292 78.64 3.448 ;
      RECT 78.596 3.301 78.605 3.452 ;
      RECT 78.51 3.319 78.596 3.469 ;
      RECT 78.451 3.346 78.51 3.496 ;
      RECT 78.365 3.373 78.451 3.524 ;
      RECT 78.345 3.395 78.365 3.544 ;
      RECT 78.285 3.41 78.345 3.56 ;
      RECT 78.275 3.422 78.285 3.573 ;
      RECT 78.27 3.427 78.275 3.576 ;
      RECT 78.26 3.43 78.27 3.579 ;
      RECT 78.255 3.432 78.26 3.582 ;
      RECT 78.225 3.44 78.255 3.589 ;
      RECT 78.21 3.447 78.225 3.597 ;
      RECT 78.2 3.452 78.21 3.601 ;
      RECT 78.195 3.455 78.2 3.604 ;
      RECT 78.185 3.457 78.195 3.607 ;
      RECT 78.15 3.467 78.185 3.616 ;
      RECT 78.075 3.49 78.15 3.638 ;
      RECT 78.055 3.508 78.075 3.656 ;
      RECT 78.025 3.515 78.055 3.666 ;
      RECT 78.005 3.523 78.025 3.676 ;
      RECT 77.995 3.529 78.005 3.683 ;
      RECT 77.976 3.534 77.995 3.689 ;
      RECT 77.89 3.554 77.976 3.709 ;
      RECT 77.875 3.574 77.89 3.728 ;
      RECT 77.83 3.586 77.875 3.739 ;
      RECT 77.765 3.607 77.83 3.762 ;
      RECT 77.725 3.627 77.765 3.783 ;
      RECT 77.715 3.637 77.725 3.793 ;
      RECT 77.665 3.649 77.715 3.804 ;
      RECT 77.645 3.665 77.665 3.816 ;
      RECT 77.615 3.675 77.645 3.822 ;
      RECT 77.605 3.68 77.615 3.824 ;
      RECT 77.536 3.681 77.605 3.83 ;
      RECT 77.45 3.683 77.536 3.84 ;
      RECT 77.44 3.684 77.45 3.845 ;
      RECT 78.71 3.71 78.9 3.92 ;
      RECT 78.7 3.715 78.91 3.913 ;
      RECT 78.685 3.715 78.91 3.878 ;
      RECT 78.605 3.6 78.865 3.86 ;
      RECT 77.52 3.13 77.705 3.425 ;
      RECT 77.51 3.13 77.705 3.423 ;
      RECT 77.495 3.13 77.71 3.418 ;
      RECT 77.495 3.13 77.715 3.415 ;
      RECT 77.49 3.13 77.715 3.413 ;
      RECT 77.485 3.385 77.715 3.403 ;
      RECT 77.49 3.13 77.75 3.39 ;
      RECT 77.45 2.165 77.71 2.425 ;
      RECT 77.26 2.09 77.346 2.423 ;
      RECT 77.235 2.094 77.39 2.419 ;
      RECT 77.346 2.086 77.39 2.419 ;
      RECT 77.346 2.087 77.395 2.418 ;
      RECT 77.26 2.092 77.41 2.417 ;
      RECT 77.235 2.1 77.45 2.416 ;
      RECT 77.23 2.095 77.41 2.411 ;
      RECT 77.22 2.11 77.45 2.318 ;
      RECT 77.22 2.162 77.65 2.318 ;
      RECT 77.22 2.155 77.63 2.318 ;
      RECT 77.22 2.142 77.6 2.318 ;
      RECT 77.22 2.13 77.54 2.318 ;
      RECT 77.22 2.115 77.515 2.318 ;
      RECT 76.42 2.745 76.555 3.04 ;
      RECT 76.68 2.768 76.685 2.955 ;
      RECT 77.4 2.665 77.545 2.9 ;
      RECT 77.56 2.665 77.565 2.89 ;
      RECT 77.595 2.676 77.6 2.87 ;
      RECT 77.59 2.668 77.595 2.875 ;
      RECT 77.57 2.665 77.59 2.88 ;
      RECT 77.565 2.665 77.57 2.888 ;
      RECT 77.555 2.665 77.56 2.893 ;
      RECT 77.545 2.665 77.555 2.898 ;
      RECT 77.375 2.667 77.4 2.9 ;
      RECT 77.325 2.674 77.375 2.9 ;
      RECT 77.32 2.679 77.325 2.9 ;
      RECT 77.281 2.684 77.32 2.901 ;
      RECT 77.195 2.696 77.281 2.902 ;
      RECT 77.186 2.706 77.195 2.902 ;
      RECT 77.1 2.715 77.186 2.904 ;
      RECT 77.076 2.725 77.1 2.906 ;
      RECT 76.99 2.736 77.076 2.907 ;
      RECT 76.96 2.747 76.99 2.909 ;
      RECT 76.93 2.752 76.96 2.911 ;
      RECT 76.905 2.758 76.93 2.914 ;
      RECT 76.89 2.763 76.905 2.915 ;
      RECT 76.845 2.769 76.89 2.915 ;
      RECT 76.84 2.774 76.845 2.916 ;
      RECT 76.82 2.774 76.84 2.918 ;
      RECT 76.8 2.772 76.82 2.923 ;
      RECT 76.765 2.771 76.8 2.93 ;
      RECT 76.735 2.77 76.765 2.94 ;
      RECT 76.685 2.769 76.735 2.95 ;
      RECT 76.595 2.766 76.68 3.04 ;
      RECT 76.57 2.76 76.595 3.04 ;
      RECT 76.555 2.75 76.57 3.04 ;
      RECT 76.37 2.745 76.42 2.96 ;
      RECT 76.36 2.75 76.37 2.95 ;
      RECT 76.6 3.225 76.86 3.485 ;
      RECT 76.6 3.225 76.89 3.378 ;
      RECT 76.6 3.225 76.925 3.363 ;
      RECT 76.855 3.145 77.045 3.355 ;
      RECT 76.845 3.15 77.055 3.348 ;
      RECT 76.81 3.22 77.055 3.348 ;
      RECT 76.84 3.162 76.86 3.485 ;
      RECT 76.825 3.21 77.055 3.348 ;
      RECT 76.83 3.182 76.86 3.485 ;
      RECT 75.91 2.25 75.98 3.355 ;
      RECT 76.645 2.355 76.905 2.615 ;
      RECT 76.225 2.401 76.24 2.61 ;
      RECT 76.561 2.414 76.645 2.565 ;
      RECT 76.475 2.411 76.561 2.565 ;
      RECT 76.436 2.409 76.475 2.565 ;
      RECT 76.35 2.407 76.436 2.565 ;
      RECT 76.29 2.405 76.35 2.576 ;
      RECT 76.255 2.403 76.29 2.594 ;
      RECT 76.24 2.401 76.255 2.605 ;
      RECT 76.21 2.401 76.225 2.618 ;
      RECT 76.2 2.401 76.21 2.623 ;
      RECT 76.175 2.4 76.2 2.628 ;
      RECT 76.16 2.395 76.175 2.634 ;
      RECT 76.155 2.388 76.16 2.639 ;
      RECT 76.13 2.379 76.155 2.645 ;
      RECT 76.085 2.358 76.13 2.658 ;
      RECT 76.075 2.342 76.085 2.668 ;
      RECT 76.06 2.335 76.075 2.678 ;
      RECT 76.05 2.328 76.06 2.695 ;
      RECT 76.045 2.325 76.05 2.725 ;
      RECT 76.04 2.323 76.045 2.755 ;
      RECT 76.035 2.321 76.04 2.792 ;
      RECT 76.02 2.317 76.035 2.859 ;
      RECT 76.02 3.15 76.03 3.35 ;
      RECT 76.015 2.313 76.02 2.985 ;
      RECT 76.015 3.137 76.02 3.355 ;
      RECT 76.01 2.311 76.015 3.07 ;
      RECT 76.01 3.127 76.015 3.355 ;
      RECT 75.995 2.282 76.01 3.355 ;
      RECT 75.98 2.255 75.995 3.355 ;
      RECT 75.905 2.25 75.91 2.605 ;
      RECT 75.905 2.66 75.91 3.355 ;
      RECT 75.89 2.25 75.905 2.583 ;
      RECT 75.9 2.682 75.905 3.355 ;
      RECT 75.89 2.722 75.9 3.355 ;
      RECT 75.855 2.25 75.89 2.525 ;
      RECT 75.885 2.757 75.89 3.355 ;
      RECT 75.87 2.812 75.885 3.355 ;
      RECT 75.865 2.877 75.87 3.355 ;
      RECT 75.85 2.925 75.865 3.355 ;
      RECT 75.825 2.25 75.855 2.48 ;
      RECT 75.845 2.98 75.85 3.355 ;
      RECT 75.83 3.04 75.845 3.355 ;
      RECT 75.825 3.088 75.83 3.353 ;
      RECT 75.82 2.25 75.825 2.473 ;
      RECT 75.82 3.12 75.825 3.348 ;
      RECT 75.795 2.25 75.82 2.465 ;
      RECT 75.785 2.255 75.795 2.455 ;
      RECT 76 3.53 76.02 3.77 ;
      RECT 75.23 3.46 75.235 3.67 ;
      RECT 76.51 3.533 76.52 3.728 ;
      RECT 76.505 3.523 76.51 3.731 ;
      RECT 76.425 3.52 76.505 3.754 ;
      RECT 76.421 3.52 76.425 3.776 ;
      RECT 76.335 3.52 76.421 3.786 ;
      RECT 76.32 3.52 76.335 3.794 ;
      RECT 76.291 3.521 76.32 3.792 ;
      RECT 76.205 3.526 76.291 3.788 ;
      RECT 76.192 3.53 76.205 3.784 ;
      RECT 76.106 3.53 76.192 3.78 ;
      RECT 76.02 3.53 76.106 3.774 ;
      RECT 75.936 3.53 76 3.768 ;
      RECT 75.85 3.53 75.936 3.763 ;
      RECT 75.83 3.53 75.85 3.759 ;
      RECT 75.77 3.525 75.83 3.756 ;
      RECT 75.742 3.519 75.77 3.753 ;
      RECT 75.656 3.514 75.742 3.749 ;
      RECT 75.57 3.508 75.656 3.743 ;
      RECT 75.495 3.49 75.57 3.738 ;
      RECT 75.46 3.467 75.495 3.734 ;
      RECT 75.45 3.457 75.46 3.733 ;
      RECT 75.395 3.455 75.45 3.732 ;
      RECT 75.32 3.455 75.395 3.728 ;
      RECT 75.31 3.455 75.32 3.723 ;
      RECT 75.295 3.455 75.31 3.715 ;
      RECT 75.245 3.457 75.295 3.693 ;
      RECT 75.235 3.46 75.245 3.673 ;
      RECT 75.225 3.465 75.23 3.668 ;
      RECT 75.22 3.47 75.225 3.663 ;
      RECT 75.345 2.635 75.605 2.895 ;
      RECT 75.345 2.65 75.625 2.86 ;
      RECT 75.345 2.655 75.635 2.855 ;
      RECT 73.33 2.115 73.59 2.375 ;
      RECT 73.32 2.145 73.59 2.355 ;
      RECT 75.24 2.06 75.5 2.32 ;
      RECT 75.235 2.135 75.24 2.321 ;
      RECT 75.21 2.14 75.235 2.323 ;
      RECT 75.195 2.147 75.21 2.326 ;
      RECT 75.135 2.165 75.195 2.331 ;
      RECT 75.105 2.185 75.135 2.338 ;
      RECT 75.08 2.193 75.105 2.343 ;
      RECT 75.055 2.201 75.08 2.345 ;
      RECT 75.037 2.205 75.055 2.344 ;
      RECT 74.951 2.203 75.037 2.344 ;
      RECT 74.865 2.201 74.951 2.344 ;
      RECT 74.779 2.199 74.865 2.343 ;
      RECT 74.693 2.197 74.779 2.343 ;
      RECT 74.607 2.195 74.693 2.343 ;
      RECT 74.521 2.193 74.607 2.343 ;
      RECT 74.435 2.191 74.521 2.342 ;
      RECT 74.417 2.19 74.435 2.342 ;
      RECT 74.331 2.189 74.417 2.342 ;
      RECT 74.245 2.187 74.331 2.342 ;
      RECT 74.159 2.186 74.245 2.341 ;
      RECT 74.073 2.185 74.159 2.341 ;
      RECT 73.987 2.183 74.073 2.341 ;
      RECT 73.901 2.182 73.987 2.341 ;
      RECT 73.815 2.18 73.901 2.34 ;
      RECT 73.791 2.178 73.815 2.34 ;
      RECT 73.705 2.171 73.791 2.34 ;
      RECT 73.676 2.163 73.705 2.34 ;
      RECT 73.59 2.155 73.676 2.34 ;
      RECT 73.31 2.152 73.32 2.35 ;
      RECT 74.815 3.115 74.82 3.465 ;
      RECT 74.585 3.205 74.725 3.465 ;
      RECT 75.06 2.89 75.105 3.1 ;
      RECT 75.115 2.901 75.125 3.095 ;
      RECT 75.105 2.893 75.115 3.1 ;
      RECT 75.04 2.89 75.06 3.105 ;
      RECT 75.01 2.89 75.04 3.128 ;
      RECT 75 2.89 75.01 3.153 ;
      RECT 74.995 2.89 75 3.163 ;
      RECT 74.94 2.89 74.995 3.203 ;
      RECT 74.935 2.89 74.94 3.243 ;
      RECT 74.93 2.892 74.935 3.248 ;
      RECT 74.915 2.902 74.93 3.259 ;
      RECT 74.87 2.96 74.915 3.295 ;
      RECT 74.86 3.015 74.87 3.329 ;
      RECT 74.845 3.042 74.86 3.345 ;
      RECT 74.835 3.069 74.845 3.465 ;
      RECT 74.82 3.092 74.835 3.465 ;
      RECT 74.81 3.132 74.815 3.465 ;
      RECT 74.805 3.142 74.81 3.465 ;
      RECT 74.8 3.157 74.805 3.465 ;
      RECT 74.79 3.162 74.8 3.465 ;
      RECT 74.725 3.185 74.79 3.465 ;
      RECT 74.225 2.68 74.415 2.89 ;
      RECT 72.8 2.605 73.06 2.865 ;
      RECT 73.15 2.6 73.245 2.81 ;
      RECT 73.125 2.615 73.135 2.81 ;
      RECT 74.415 2.687 74.425 2.885 ;
      RECT 74.215 2.687 74.225 2.885 ;
      RECT 74.2 2.702 74.215 2.875 ;
      RECT 74.195 2.71 74.2 2.868 ;
      RECT 74.185 2.713 74.195 2.865 ;
      RECT 74.15 2.712 74.185 2.863 ;
      RECT 74.121 2.708 74.15 2.86 ;
      RECT 74.035 2.703 74.121 2.857 ;
      RECT 73.975 2.697 74.035 2.853 ;
      RECT 73.946 2.693 73.975 2.85 ;
      RECT 73.86 2.685 73.946 2.847 ;
      RECT 73.851 2.679 73.86 2.845 ;
      RECT 73.765 2.674 73.851 2.843 ;
      RECT 73.742 2.669 73.765 2.84 ;
      RECT 73.656 2.663 73.742 2.837 ;
      RECT 73.57 2.654 73.656 2.832 ;
      RECT 73.56 2.649 73.57 2.83 ;
      RECT 73.541 2.648 73.56 2.829 ;
      RECT 73.455 2.643 73.541 2.825 ;
      RECT 73.435 2.638 73.455 2.821 ;
      RECT 73.375 2.633 73.435 2.818 ;
      RECT 73.35 2.623 73.375 2.816 ;
      RECT 73.345 2.616 73.35 2.815 ;
      RECT 73.335 2.607 73.345 2.814 ;
      RECT 73.331 2.6 73.335 2.814 ;
      RECT 73.245 2.6 73.331 2.812 ;
      RECT 73.135 2.607 73.15 2.81 ;
      RECT 73.12 2.617 73.125 2.81 ;
      RECT 73.1 2.62 73.12 2.807 ;
      RECT 73.07 2.62 73.1 2.803 ;
      RECT 73.06 2.62 73.07 2.803 ;
      RECT 73.975 3.115 74.235 3.375 ;
      RECT 73.905 3.125 74.235 3.335 ;
      RECT 73.895 3.132 74.235 3.33 ;
      RECT 73.315 3.12 73.575 3.38 ;
      RECT 73.315 3.16 73.68 3.37 ;
      RECT 73.315 3.162 73.685 3.369 ;
      RECT 73.315 3.17 73.69 3.366 ;
      RECT 72.24 2.245 72.34 3.77 ;
      RECT 72.43 3.385 72.48 3.645 ;
      RECT 72.425 2.258 72.43 2.445 ;
      RECT 72.42 3.366 72.43 3.645 ;
      RECT 72.42 2.255 72.425 2.453 ;
      RECT 72.405 2.249 72.42 2.46 ;
      RECT 72.415 3.354 72.42 3.728 ;
      RECT 72.405 3.342 72.415 3.765 ;
      RECT 72.395 2.245 72.405 2.467 ;
      RECT 72.395 3.327 72.405 3.77 ;
      RECT 72.39 2.245 72.395 2.475 ;
      RECT 72.37 3.297 72.395 3.77 ;
      RECT 72.35 2.245 72.39 2.523 ;
      RECT 72.36 3.257 72.37 3.77 ;
      RECT 72.35 3.212 72.36 3.77 ;
      RECT 72.345 2.245 72.35 2.593 ;
      RECT 72.345 3.17 72.35 3.77 ;
      RECT 72.34 2.245 72.345 3.07 ;
      RECT 72.34 3.152 72.345 3.77 ;
      RECT 72.23 2.248 72.24 3.77 ;
      RECT 72.215 2.255 72.23 3.766 ;
      RECT 72.21 2.265 72.215 3.761 ;
      RECT 72.205 2.465 72.21 3.653 ;
      RECT 72.2 2.55 72.205 3.205 ;
      RECT 71.085 2.365 71.375 2.595 ;
      RECT 71.145 0.885 71.315 2.595 ;
      RECT 71.145 0.885 71.325 1.45 ;
      RECT 71.12 1.095 71.47 1.445 ;
      RECT 71.085 0.885 71.375 1.115 ;
      RECT 71.085 7.765 71.375 7.995 ;
      RECT 71.145 6.285 71.315 7.995 ;
      RECT 71.085 6.285 71.375 6.515 ;
      RECT 70.675 2.735 71.005 2.965 ;
      RECT 70.675 2.765 71.175 2.935 ;
      RECT 70.675 2.395 70.865 2.965 ;
      RECT 70.095 2.365 70.385 2.595 ;
      RECT 70.095 2.395 70.865 2.565 ;
      RECT 70.155 0.885 70.325 2.595 ;
      RECT 70.095 0.885 70.385 1.115 ;
      RECT 70.095 7.765 70.385 7.995 ;
      RECT 70.155 6.285 70.325 7.995 ;
      RECT 70.095 6.285 70.385 6.515 ;
      RECT 70.095 6.325 70.945 6.485 ;
      RECT 70.775 5.915 70.945 6.485 ;
      RECT 70.095 6.32 70.485 6.485 ;
      RECT 70.715 5.915 71.005 6.145 ;
      RECT 70.715 5.945 71.175 6.115 ;
      RECT 69.725 2.735 70.015 2.965 ;
      RECT 69.725 2.765 70.185 2.935 ;
      RECT 69.785 1.655 69.95 2.965 ;
      RECT 68.3 1.625 68.59 1.855 ;
      RECT 68.3 1.655 69.95 1.825 ;
      RECT 68.36 0.885 68.53 1.855 ;
      RECT 68.3 0.885 68.59 1.115 ;
      RECT 68.3 7.765 68.59 7.995 ;
      RECT 68.36 7.025 68.53 7.995 ;
      RECT 68.36 7.12 69.95 7.29 ;
      RECT 69.78 5.915 69.95 7.29 ;
      RECT 68.3 7.025 68.59 7.255 ;
      RECT 69.725 5.915 70.015 6.145 ;
      RECT 69.725 5.945 70.185 6.115 ;
      RECT 68.73 1.965 69.08 2.315 ;
      RECT 68.56 2.025 69.08 2.195 ;
      RECT 68.755 6.655 69.08 6.98 ;
      RECT 68.73 6.655 69.08 6.885 ;
      RECT 68.56 6.685 69.08 6.855 ;
      RECT 66.335 3.43 66.685 3.78 ;
      RECT 66.425 2.395 66.595 3.78 ;
      RECT 67.955 2.365 68.275 2.685 ;
      RECT 67.925 2.365 68.275 2.595 ;
      RECT 66.425 2.395 68.275 2.565 ;
      RECT 67.955 6.28 68.275 6.605 ;
      RECT 67.925 6.285 68.275 6.515 ;
      RECT 67.755 6.315 68.275 6.485 ;
      RECT 66.91 2.705 67.26 3.055 ;
      RECT 66.91 2.765 67.39 2.935 ;
      RECT 66.9 5.84 67.25 6.19 ;
      RECT 66.9 5.945 67.39 6.115 ;
      RECT 63.735 3.665 63.775 3.925 ;
      RECT 63.775 3.645 63.78 3.655 ;
      RECT 65.115 2.735 65.27 3.055 ;
      RECT 65.035 2.735 65.115 3.22 ;
      RECT 65.025 2.735 65.035 3.363 ;
      RECT 65 2.735 65.025 3.41 ;
      RECT 64.975 2.735 65 3.488 ;
      RECT 64.955 2.735 64.975 3.558 ;
      RECT 64.95 2.735 64.955 3.588 ;
      RECT 64.93 2.885 64.95 3.6 ;
      RECT 64.92 2.885 64.93 3.618 ;
      RECT 64.91 2.887 64.92 3.626 ;
      RECT 64.905 2.892 64.91 3.083 ;
      RECT 64.905 3.092 64.91 3.627 ;
      RECT 64.9 3.137 64.905 3.628 ;
      RECT 64.89 3.202 64.9 3.629 ;
      RECT 64.88 3.297 64.89 3.631 ;
      RECT 64.875 3.35 64.88 3.633 ;
      RECT 64.87 3.37 64.875 3.634 ;
      RECT 64.815 3.395 64.87 3.64 ;
      RECT 64.775 3.43 64.815 3.649 ;
      RECT 64.765 3.447 64.775 3.654 ;
      RECT 64.756 3.453 64.765 3.656 ;
      RECT 64.67 3.491 64.756 3.667 ;
      RECT 64.665 3.53 64.67 3.677 ;
      RECT 64.59 3.537 64.665 3.687 ;
      RECT 64.57 3.547 64.59 3.698 ;
      RECT 64.54 3.554 64.57 3.706 ;
      RECT 64.515 3.561 64.54 3.713 ;
      RECT 64.491 3.567 64.515 3.718 ;
      RECT 64.405 3.58 64.491 3.73 ;
      RECT 64.327 3.587 64.405 3.748 ;
      RECT 64.241 3.582 64.327 3.766 ;
      RECT 64.155 3.577 64.241 3.786 ;
      RECT 64.075 3.571 64.155 3.803 ;
      RECT 64.01 3.567 64.075 3.832 ;
      RECT 64.005 3.281 64.01 3.305 ;
      RECT 63.995 3.557 64.01 3.86 ;
      RECT 64 3.275 64.005 3.345 ;
      RECT 63.995 3.269 64 3.415 ;
      RECT 63.99 3.263 63.995 3.493 ;
      RECT 63.99 3.54 63.995 3.925 ;
      RECT 63.982 3.26 63.99 3.925 ;
      RECT 63.896 3.258 63.982 3.925 ;
      RECT 63.81 3.256 63.896 3.925 ;
      RECT 63.8 3.257 63.81 3.925 ;
      RECT 63.795 3.262 63.8 3.925 ;
      RECT 63.785 3.275 63.795 3.925 ;
      RECT 63.78 3.297 63.785 3.925 ;
      RECT 63.775 3.657 63.78 3.925 ;
      RECT 64.405 3.125 64.41 3.345 ;
      RECT 64.91 2.16 64.945 2.42 ;
      RECT 64.895 2.16 64.91 2.428 ;
      RECT 64.866 2.16 64.895 2.45 ;
      RECT 64.78 2.16 64.866 2.51 ;
      RECT 64.76 2.16 64.78 2.575 ;
      RECT 64.7 2.16 64.76 2.74 ;
      RECT 64.695 2.16 64.7 2.888 ;
      RECT 64.69 2.16 64.695 2.9 ;
      RECT 64.685 2.16 64.69 2.926 ;
      RECT 64.655 2.346 64.685 3.006 ;
      RECT 64.65 2.394 64.655 3.095 ;
      RECT 64.645 2.408 64.65 3.11 ;
      RECT 64.64 2.427 64.645 3.14 ;
      RECT 64.635 2.442 64.64 3.156 ;
      RECT 64.63 2.457 64.635 3.178 ;
      RECT 64.625 2.477 64.63 3.2 ;
      RECT 64.615 2.497 64.625 3.233 ;
      RECT 64.6 2.539 64.615 3.295 ;
      RECT 64.595 2.57 64.6 3.335 ;
      RECT 64.59 2.582 64.595 3.34 ;
      RECT 64.585 2.594 64.59 3.345 ;
      RECT 64.58 2.607 64.585 3.345 ;
      RECT 64.575 2.625 64.58 3.345 ;
      RECT 64.57 2.645 64.575 3.345 ;
      RECT 64.565 2.657 64.57 3.345 ;
      RECT 64.56 2.67 64.565 3.345 ;
      RECT 64.54 2.705 64.56 3.345 ;
      RECT 64.49 2.807 64.54 3.345 ;
      RECT 64.485 2.892 64.49 3.345 ;
      RECT 64.48 2.9 64.485 3.345 ;
      RECT 64.475 2.917 64.48 3.345 ;
      RECT 64.47 2.932 64.475 3.345 ;
      RECT 64.435 2.997 64.47 3.345 ;
      RECT 64.42 3.062 64.435 3.345 ;
      RECT 64.415 3.092 64.42 3.345 ;
      RECT 64.41 3.117 64.415 3.345 ;
      RECT 64.395 3.127 64.405 3.345 ;
      RECT 64.38 3.14 64.395 3.338 ;
      RECT 64.125 2.73 64.195 2.94 ;
      RECT 63.915 2.707 63.92 2.9 ;
      RECT 61.37 2.635 61.63 2.895 ;
      RECT 64.205 2.917 64.21 2.92 ;
      RECT 64.195 2.735 64.205 2.935 ;
      RECT 64.096 2.728 64.125 2.94 ;
      RECT 64.01 2.72 64.096 2.94 ;
      RECT 63.995 2.714 64.01 2.938 ;
      RECT 63.975 2.713 63.995 2.925 ;
      RECT 63.97 2.712 63.975 2.908 ;
      RECT 63.92 2.709 63.97 2.903 ;
      RECT 63.89 2.706 63.915 2.898 ;
      RECT 63.87 2.704 63.89 2.893 ;
      RECT 63.855 2.702 63.87 2.89 ;
      RECT 63.825 2.7 63.855 2.888 ;
      RECT 63.76 2.696 63.825 2.88 ;
      RECT 63.73 2.691 63.76 2.875 ;
      RECT 63.71 2.689 63.73 2.873 ;
      RECT 63.68 2.686 63.71 2.868 ;
      RECT 63.62 2.682 63.68 2.86 ;
      RECT 63.615 2.679 63.62 2.855 ;
      RECT 63.545 2.677 63.615 2.85 ;
      RECT 63.516 2.673 63.545 2.843 ;
      RECT 63.43 2.668 63.516 2.835 ;
      RECT 63.396 2.663 63.43 2.827 ;
      RECT 63.31 2.655 63.396 2.819 ;
      RECT 63.271 2.648 63.31 2.811 ;
      RECT 63.185 2.643 63.271 2.803 ;
      RECT 63.12 2.637 63.185 2.793 ;
      RECT 63.1 2.632 63.12 2.788 ;
      RECT 63.091 2.629 63.1 2.787 ;
      RECT 63.005 2.625 63.091 2.781 ;
      RECT 62.965 2.621 63.005 2.773 ;
      RECT 62.945 2.617 62.965 2.771 ;
      RECT 62.885 2.617 62.945 2.768 ;
      RECT 62.865 2.62 62.885 2.766 ;
      RECT 62.844 2.62 62.865 2.766 ;
      RECT 62.758 2.622 62.844 2.77 ;
      RECT 62.672 2.624 62.758 2.776 ;
      RECT 62.586 2.626 62.672 2.783 ;
      RECT 62.5 2.629 62.586 2.789 ;
      RECT 62.466 2.63 62.5 2.794 ;
      RECT 62.38 2.633 62.466 2.799 ;
      RECT 62.351 2.64 62.38 2.804 ;
      RECT 62.265 2.64 62.351 2.809 ;
      RECT 62.232 2.64 62.265 2.814 ;
      RECT 62.146 2.642 62.232 2.819 ;
      RECT 62.06 2.644 62.146 2.826 ;
      RECT 61.996 2.646 62.06 2.832 ;
      RECT 61.91 2.648 61.996 2.838 ;
      RECT 61.907 2.65 61.91 2.841 ;
      RECT 61.821 2.651 61.907 2.845 ;
      RECT 61.735 2.654 61.821 2.852 ;
      RECT 61.716 2.656 61.735 2.856 ;
      RECT 61.63 2.658 61.716 2.861 ;
      RECT 61.36 2.67 61.37 2.865 ;
      RECT 63.595 2.25 63.78 2.46 ;
      RECT 63.59 2.251 63.785 2.458 ;
      RECT 63.585 2.256 63.795 2.453 ;
      RECT 63.58 2.232 63.585 2.45 ;
      RECT 63.55 2.229 63.58 2.443 ;
      RECT 63.545 2.225 63.55 2.434 ;
      RECT 63.51 2.256 63.795 2.429 ;
      RECT 63.285 2.165 63.545 2.425 ;
      RECT 63.585 2.234 63.59 2.453 ;
      RECT 63.59 2.235 63.595 2.458 ;
      RECT 63.285 2.247 63.665 2.425 ;
      RECT 63.285 2.245 63.65 2.425 ;
      RECT 63.285 2.24 63.64 2.425 ;
      RECT 63.24 3.155 63.29 3.44 ;
      RECT 63.185 3.125 63.19 3.44 ;
      RECT 63.155 3.105 63.16 3.44 ;
      RECT 63.305 3.155 63.365 3.415 ;
      RECT 63.3 3.155 63.305 3.423 ;
      RECT 63.29 3.155 63.3 3.435 ;
      RECT 63.205 3.145 63.24 3.44 ;
      RECT 63.2 3.132 63.205 3.44 ;
      RECT 63.19 3.127 63.2 3.44 ;
      RECT 63.17 3.117 63.185 3.44 ;
      RECT 63.16 3.11 63.17 3.44 ;
      RECT 63.15 3.102 63.155 3.44 ;
      RECT 63.12 3.092 63.15 3.44 ;
      RECT 63.105 3.08 63.12 3.44 ;
      RECT 63.09 3.07 63.105 3.435 ;
      RECT 63.07 3.06 63.09 3.41 ;
      RECT 63.06 3.052 63.07 3.387 ;
      RECT 63.03 3.035 63.06 3.377 ;
      RECT 63.025 3.012 63.03 3.368 ;
      RECT 63.02 2.999 63.025 3.366 ;
      RECT 63.005 2.975 63.02 3.36 ;
      RECT 63 2.951 63.005 3.354 ;
      RECT 62.99 2.94 63 3.349 ;
      RECT 62.985 2.93 62.99 3.345 ;
      RECT 62.98 2.922 62.985 3.342 ;
      RECT 62.97 2.917 62.98 3.338 ;
      RECT 62.965 2.912 62.97 3.334 ;
      RECT 62.88 2.91 62.965 3.309 ;
      RECT 62.85 2.91 62.88 3.275 ;
      RECT 62.835 2.91 62.85 3.258 ;
      RECT 62.78 2.91 62.835 3.203 ;
      RECT 62.775 2.915 62.78 3.152 ;
      RECT 62.765 2.92 62.775 3.142 ;
      RECT 62.76 2.93 62.765 3.128 ;
      RECT 62.71 3.67 62.97 3.93 ;
      RECT 62.63 3.685 62.97 3.906 ;
      RECT 62.61 3.685 62.97 3.901 ;
      RECT 62.586 3.685 62.97 3.899 ;
      RECT 62.5 3.685 62.97 3.894 ;
      RECT 62.35 3.625 62.61 3.89 ;
      RECT 62.305 3.685 62.97 3.885 ;
      RECT 62.3 3.692 62.97 3.88 ;
      RECT 62.315 3.68 62.63 3.89 ;
      RECT 62.205 2.115 62.465 2.375 ;
      RECT 62.205 2.172 62.47 2.368 ;
      RECT 62.205 2.202 62.475 2.3 ;
      RECT 62.265 2.633 62.38 2.635 ;
      RECT 62.351 2.63 62.38 2.635 ;
      RECT 61.375 3.634 61.4 3.874 ;
      RECT 61.36 3.637 61.45 3.868 ;
      RECT 61.355 3.642 61.536 3.863 ;
      RECT 61.35 3.65 61.6 3.861 ;
      RECT 61.35 3.65 61.61 3.86 ;
      RECT 61.345 3.657 61.62 3.853 ;
      RECT 61.345 3.657 61.706 3.842 ;
      RECT 61.34 3.692 61.706 3.838 ;
      RECT 61.34 3.692 61.715 3.827 ;
      RECT 61.62 3.565 61.88 3.825 ;
      RECT 61.33 3.742 61.88 3.823 ;
      RECT 61.6 3.61 61.62 3.858 ;
      RECT 61.536 3.613 61.6 3.862 ;
      RECT 61.45 3.618 61.536 3.867 ;
      RECT 61.38 3.629 61.88 3.825 ;
      RECT 61.4 3.623 61.45 3.872 ;
      RECT 61.525 2.1 61.535 2.362 ;
      RECT 61.515 2.157 61.525 2.365 ;
      RECT 61.49 2.162 61.515 2.371 ;
      RECT 61.465 2.166 61.49 2.383 ;
      RECT 61.455 2.169 61.465 2.393 ;
      RECT 61.45 2.17 61.455 2.398 ;
      RECT 61.445 2.171 61.45 2.403 ;
      RECT 61.44 2.172 61.445 2.405 ;
      RECT 61.415 2.175 61.44 2.408 ;
      RECT 61.385 2.181 61.415 2.411 ;
      RECT 61.32 2.192 61.385 2.414 ;
      RECT 61.275 2.2 61.32 2.418 ;
      RECT 61.26 2.2 61.275 2.426 ;
      RECT 61.255 2.201 61.26 2.433 ;
      RECT 61.25 2.203 61.255 2.436 ;
      RECT 61.245 2.207 61.25 2.439 ;
      RECT 61.235 2.215 61.245 2.443 ;
      RECT 61.23 2.228 61.235 2.448 ;
      RECT 61.225 2.236 61.23 2.45 ;
      RECT 61.22 2.242 61.225 2.45 ;
      RECT 61.215 2.246 61.22 2.453 ;
      RECT 61.21 2.248 61.215 2.456 ;
      RECT 61.205 2.251 61.21 2.459 ;
      RECT 61.195 2.256 61.205 2.463 ;
      RECT 61.19 2.262 61.195 2.468 ;
      RECT 61.18 2.268 61.19 2.472 ;
      RECT 61.165 2.275 61.18 2.478 ;
      RECT 61.136 2.289 61.165 2.488 ;
      RECT 61.05 2.324 61.136 2.52 ;
      RECT 61.03 2.357 61.05 2.549 ;
      RECT 61.01 2.37 61.03 2.56 ;
      RECT 60.99 2.382 61.01 2.571 ;
      RECT 60.94 2.404 60.99 2.591 ;
      RECT 60.925 2.422 60.94 2.608 ;
      RECT 60.92 2.428 60.925 2.611 ;
      RECT 60.915 2.432 60.92 2.614 ;
      RECT 60.91 2.436 60.915 2.618 ;
      RECT 60.905 2.438 60.91 2.621 ;
      RECT 60.895 2.445 60.905 2.624 ;
      RECT 60.89 2.45 60.895 2.628 ;
      RECT 60.885 2.452 60.89 2.631 ;
      RECT 60.88 2.456 60.885 2.634 ;
      RECT 60.875 2.458 60.88 2.638 ;
      RECT 60.86 2.463 60.875 2.643 ;
      RECT 60.855 2.468 60.86 2.646 ;
      RECT 60.85 2.476 60.855 2.649 ;
      RECT 60.845 2.478 60.85 2.652 ;
      RECT 60.84 2.48 60.845 2.655 ;
      RECT 60.83 2.482 60.84 2.661 ;
      RECT 60.795 2.496 60.83 2.673 ;
      RECT 60.785 2.511 60.795 2.683 ;
      RECT 60.71 2.54 60.785 2.707 ;
      RECT 60.705 2.565 60.71 2.73 ;
      RECT 60.69 2.569 60.705 2.736 ;
      RECT 60.68 2.577 60.69 2.741 ;
      RECT 60.65 2.59 60.68 2.745 ;
      RECT 60.64 2.605 60.65 2.75 ;
      RECT 60.63 2.61 60.64 2.753 ;
      RECT 60.625 2.612 60.63 2.755 ;
      RECT 60.61 2.615 60.625 2.758 ;
      RECT 60.605 2.617 60.61 2.761 ;
      RECT 60.585 2.622 60.605 2.765 ;
      RECT 60.555 2.627 60.585 2.773 ;
      RECT 60.53 2.634 60.555 2.781 ;
      RECT 60.525 2.639 60.53 2.786 ;
      RECT 60.495 2.642 60.525 2.79 ;
      RECT 60.455 2.645 60.495 2.8 ;
      RECT 60.42 2.642 60.455 2.812 ;
      RECT 60.41 2.638 60.42 2.819 ;
      RECT 60.385 2.634 60.41 2.825 ;
      RECT 60.38 2.63 60.385 2.83 ;
      RECT 60.34 2.627 60.38 2.83 ;
      RECT 60.325 2.612 60.34 2.831 ;
      RECT 60.302 2.6 60.325 2.831 ;
      RECT 60.216 2.6 60.302 2.832 ;
      RECT 60.13 2.6 60.216 2.834 ;
      RECT 60.11 2.6 60.13 2.831 ;
      RECT 60.105 2.605 60.11 2.826 ;
      RECT 60.1 2.61 60.105 2.824 ;
      RECT 60.09 2.62 60.1 2.822 ;
      RECT 60.085 2.626 60.09 2.815 ;
      RECT 60.08 2.628 60.085 2.8 ;
      RECT 60.075 2.632 60.08 2.79 ;
      RECT 61.535 2.1 61.785 2.36 ;
      RECT 59.26 3.635 59.52 3.895 ;
      RECT 61.555 3.125 61.56 3.335 ;
      RECT 61.56 3.13 61.57 3.33 ;
      RECT 61.51 3.125 61.555 3.35 ;
      RECT 61.5 3.125 61.51 3.37 ;
      RECT 61.481 3.125 61.5 3.375 ;
      RECT 61.395 3.125 61.481 3.372 ;
      RECT 61.365 3.127 61.395 3.37 ;
      RECT 61.31 3.137 61.365 3.368 ;
      RECT 61.245 3.151 61.31 3.366 ;
      RECT 61.24 3.159 61.245 3.365 ;
      RECT 61.225 3.162 61.24 3.363 ;
      RECT 61.16 3.172 61.225 3.359 ;
      RECT 61.112 3.186 61.16 3.36 ;
      RECT 61.026 3.203 61.112 3.374 ;
      RECT 60.94 3.224 61.026 3.391 ;
      RECT 60.92 3.237 60.94 3.401 ;
      RECT 60.875 3.245 60.92 3.408 ;
      RECT 60.84 3.253 60.875 3.416 ;
      RECT 60.806 3.261 60.84 3.424 ;
      RECT 60.72 3.275 60.806 3.436 ;
      RECT 60.685 3.292 60.72 3.448 ;
      RECT 60.676 3.301 60.685 3.452 ;
      RECT 60.59 3.319 60.676 3.469 ;
      RECT 60.531 3.346 60.59 3.496 ;
      RECT 60.445 3.373 60.531 3.524 ;
      RECT 60.425 3.395 60.445 3.544 ;
      RECT 60.365 3.41 60.425 3.56 ;
      RECT 60.355 3.422 60.365 3.573 ;
      RECT 60.35 3.427 60.355 3.576 ;
      RECT 60.34 3.43 60.35 3.579 ;
      RECT 60.335 3.432 60.34 3.582 ;
      RECT 60.305 3.44 60.335 3.589 ;
      RECT 60.29 3.447 60.305 3.597 ;
      RECT 60.28 3.452 60.29 3.601 ;
      RECT 60.275 3.455 60.28 3.604 ;
      RECT 60.265 3.457 60.275 3.607 ;
      RECT 60.23 3.467 60.265 3.616 ;
      RECT 60.155 3.49 60.23 3.638 ;
      RECT 60.135 3.508 60.155 3.656 ;
      RECT 60.105 3.515 60.135 3.666 ;
      RECT 60.085 3.523 60.105 3.676 ;
      RECT 60.075 3.529 60.085 3.683 ;
      RECT 60.056 3.534 60.075 3.689 ;
      RECT 59.97 3.554 60.056 3.709 ;
      RECT 59.955 3.574 59.97 3.728 ;
      RECT 59.91 3.586 59.955 3.739 ;
      RECT 59.845 3.607 59.91 3.762 ;
      RECT 59.805 3.627 59.845 3.783 ;
      RECT 59.795 3.637 59.805 3.793 ;
      RECT 59.745 3.649 59.795 3.804 ;
      RECT 59.725 3.665 59.745 3.816 ;
      RECT 59.695 3.675 59.725 3.822 ;
      RECT 59.685 3.68 59.695 3.824 ;
      RECT 59.616 3.681 59.685 3.83 ;
      RECT 59.53 3.683 59.616 3.84 ;
      RECT 59.52 3.684 59.53 3.845 ;
      RECT 60.79 3.71 60.98 3.92 ;
      RECT 60.78 3.715 60.99 3.913 ;
      RECT 60.765 3.715 60.99 3.878 ;
      RECT 60.685 3.6 60.945 3.86 ;
      RECT 59.6 3.13 59.785 3.425 ;
      RECT 59.59 3.13 59.785 3.423 ;
      RECT 59.575 3.13 59.79 3.418 ;
      RECT 59.575 3.13 59.795 3.415 ;
      RECT 59.57 3.13 59.795 3.413 ;
      RECT 59.565 3.385 59.795 3.403 ;
      RECT 59.57 3.13 59.83 3.39 ;
      RECT 59.53 2.165 59.79 2.425 ;
      RECT 59.34 2.09 59.426 2.423 ;
      RECT 59.315 2.094 59.47 2.419 ;
      RECT 59.426 2.086 59.47 2.419 ;
      RECT 59.426 2.087 59.475 2.418 ;
      RECT 59.34 2.092 59.49 2.417 ;
      RECT 59.315 2.1 59.53 2.416 ;
      RECT 59.31 2.095 59.49 2.411 ;
      RECT 59.3 2.11 59.53 2.318 ;
      RECT 59.3 2.162 59.73 2.318 ;
      RECT 59.3 2.155 59.71 2.318 ;
      RECT 59.3 2.142 59.68 2.318 ;
      RECT 59.3 2.13 59.62 2.318 ;
      RECT 59.3 2.115 59.595 2.318 ;
      RECT 58.5 2.745 58.635 3.04 ;
      RECT 58.76 2.768 58.765 2.955 ;
      RECT 59.48 2.665 59.625 2.9 ;
      RECT 59.64 2.665 59.645 2.89 ;
      RECT 59.675 2.676 59.68 2.87 ;
      RECT 59.67 2.668 59.675 2.875 ;
      RECT 59.65 2.665 59.67 2.88 ;
      RECT 59.645 2.665 59.65 2.888 ;
      RECT 59.635 2.665 59.64 2.893 ;
      RECT 59.625 2.665 59.635 2.898 ;
      RECT 59.455 2.667 59.48 2.9 ;
      RECT 59.405 2.674 59.455 2.9 ;
      RECT 59.4 2.679 59.405 2.9 ;
      RECT 59.361 2.684 59.4 2.901 ;
      RECT 59.275 2.696 59.361 2.902 ;
      RECT 59.266 2.706 59.275 2.902 ;
      RECT 59.18 2.715 59.266 2.904 ;
      RECT 59.156 2.725 59.18 2.906 ;
      RECT 59.07 2.736 59.156 2.907 ;
      RECT 59.04 2.747 59.07 2.909 ;
      RECT 59.01 2.752 59.04 2.911 ;
      RECT 58.985 2.758 59.01 2.914 ;
      RECT 58.97 2.763 58.985 2.915 ;
      RECT 58.925 2.769 58.97 2.915 ;
      RECT 58.92 2.774 58.925 2.916 ;
      RECT 58.9 2.774 58.92 2.918 ;
      RECT 58.88 2.772 58.9 2.923 ;
      RECT 58.845 2.771 58.88 2.93 ;
      RECT 58.815 2.77 58.845 2.94 ;
      RECT 58.765 2.769 58.815 2.95 ;
      RECT 58.675 2.766 58.76 3.04 ;
      RECT 58.65 2.76 58.675 3.04 ;
      RECT 58.635 2.75 58.65 3.04 ;
      RECT 58.45 2.745 58.5 2.96 ;
      RECT 58.44 2.75 58.45 2.95 ;
      RECT 58.68 3.225 58.94 3.485 ;
      RECT 58.68 3.225 58.97 3.378 ;
      RECT 58.68 3.225 59.005 3.363 ;
      RECT 58.935 3.145 59.125 3.355 ;
      RECT 58.925 3.15 59.135 3.348 ;
      RECT 58.89 3.22 59.135 3.348 ;
      RECT 58.92 3.162 58.94 3.485 ;
      RECT 58.905 3.21 59.135 3.348 ;
      RECT 58.91 3.182 58.94 3.485 ;
      RECT 57.99 2.25 58.06 3.355 ;
      RECT 58.725 2.355 58.985 2.615 ;
      RECT 58.305 2.401 58.32 2.61 ;
      RECT 58.641 2.414 58.725 2.565 ;
      RECT 58.555 2.411 58.641 2.565 ;
      RECT 58.516 2.409 58.555 2.565 ;
      RECT 58.43 2.407 58.516 2.565 ;
      RECT 58.37 2.405 58.43 2.576 ;
      RECT 58.335 2.403 58.37 2.594 ;
      RECT 58.32 2.401 58.335 2.605 ;
      RECT 58.29 2.401 58.305 2.618 ;
      RECT 58.28 2.401 58.29 2.623 ;
      RECT 58.255 2.4 58.28 2.628 ;
      RECT 58.24 2.395 58.255 2.634 ;
      RECT 58.235 2.388 58.24 2.639 ;
      RECT 58.21 2.379 58.235 2.645 ;
      RECT 58.165 2.358 58.21 2.658 ;
      RECT 58.155 2.342 58.165 2.668 ;
      RECT 58.14 2.335 58.155 2.678 ;
      RECT 58.13 2.328 58.14 2.695 ;
      RECT 58.125 2.325 58.13 2.725 ;
      RECT 58.12 2.323 58.125 2.755 ;
      RECT 58.115 2.321 58.12 2.792 ;
      RECT 58.1 2.317 58.115 2.859 ;
      RECT 58.1 3.15 58.11 3.35 ;
      RECT 58.095 2.313 58.1 2.985 ;
      RECT 58.095 3.137 58.1 3.355 ;
      RECT 58.09 2.311 58.095 3.07 ;
      RECT 58.09 3.127 58.095 3.355 ;
      RECT 58.075 2.282 58.09 3.355 ;
      RECT 58.06 2.255 58.075 3.355 ;
      RECT 57.985 2.25 57.99 2.605 ;
      RECT 57.985 2.66 57.99 3.355 ;
      RECT 57.97 2.25 57.985 2.583 ;
      RECT 57.98 2.682 57.985 3.355 ;
      RECT 57.97 2.722 57.98 3.355 ;
      RECT 57.935 2.25 57.97 2.525 ;
      RECT 57.965 2.757 57.97 3.355 ;
      RECT 57.95 2.812 57.965 3.355 ;
      RECT 57.945 2.877 57.95 3.355 ;
      RECT 57.93 2.925 57.945 3.355 ;
      RECT 57.905 2.25 57.935 2.48 ;
      RECT 57.925 2.98 57.93 3.355 ;
      RECT 57.91 3.04 57.925 3.355 ;
      RECT 57.905 3.088 57.91 3.353 ;
      RECT 57.9 2.25 57.905 2.473 ;
      RECT 57.9 3.12 57.905 3.348 ;
      RECT 57.875 2.25 57.9 2.465 ;
      RECT 57.865 2.255 57.875 2.455 ;
      RECT 58.08 3.53 58.1 3.77 ;
      RECT 57.31 3.46 57.315 3.67 ;
      RECT 58.59 3.533 58.6 3.728 ;
      RECT 58.585 3.523 58.59 3.731 ;
      RECT 58.505 3.52 58.585 3.754 ;
      RECT 58.501 3.52 58.505 3.776 ;
      RECT 58.415 3.52 58.501 3.786 ;
      RECT 58.4 3.52 58.415 3.794 ;
      RECT 58.371 3.521 58.4 3.792 ;
      RECT 58.285 3.526 58.371 3.788 ;
      RECT 58.272 3.53 58.285 3.784 ;
      RECT 58.186 3.53 58.272 3.78 ;
      RECT 58.1 3.53 58.186 3.774 ;
      RECT 58.016 3.53 58.08 3.768 ;
      RECT 57.93 3.53 58.016 3.763 ;
      RECT 57.91 3.53 57.93 3.759 ;
      RECT 57.85 3.525 57.91 3.756 ;
      RECT 57.822 3.519 57.85 3.753 ;
      RECT 57.736 3.514 57.822 3.749 ;
      RECT 57.65 3.508 57.736 3.743 ;
      RECT 57.575 3.49 57.65 3.738 ;
      RECT 57.54 3.467 57.575 3.734 ;
      RECT 57.53 3.457 57.54 3.733 ;
      RECT 57.475 3.455 57.53 3.732 ;
      RECT 57.4 3.455 57.475 3.728 ;
      RECT 57.39 3.455 57.4 3.723 ;
      RECT 57.375 3.455 57.39 3.715 ;
      RECT 57.325 3.457 57.375 3.693 ;
      RECT 57.315 3.46 57.325 3.673 ;
      RECT 57.305 3.465 57.31 3.668 ;
      RECT 57.3 3.47 57.305 3.663 ;
      RECT 57.425 2.635 57.685 2.895 ;
      RECT 57.425 2.65 57.705 2.86 ;
      RECT 57.425 2.655 57.715 2.855 ;
      RECT 55.41 2.115 55.67 2.375 ;
      RECT 55.4 2.145 55.67 2.355 ;
      RECT 57.32 2.06 57.58 2.32 ;
      RECT 57.315 2.135 57.32 2.321 ;
      RECT 57.29 2.14 57.315 2.323 ;
      RECT 57.275 2.147 57.29 2.326 ;
      RECT 57.215 2.165 57.275 2.331 ;
      RECT 57.185 2.185 57.215 2.338 ;
      RECT 57.16 2.193 57.185 2.343 ;
      RECT 57.135 2.201 57.16 2.345 ;
      RECT 57.117 2.205 57.135 2.344 ;
      RECT 57.031 2.203 57.117 2.344 ;
      RECT 56.945 2.201 57.031 2.344 ;
      RECT 56.859 2.199 56.945 2.343 ;
      RECT 56.773 2.197 56.859 2.343 ;
      RECT 56.687 2.195 56.773 2.343 ;
      RECT 56.601 2.193 56.687 2.343 ;
      RECT 56.515 2.191 56.601 2.342 ;
      RECT 56.497 2.19 56.515 2.342 ;
      RECT 56.411 2.189 56.497 2.342 ;
      RECT 56.325 2.187 56.411 2.342 ;
      RECT 56.239 2.186 56.325 2.341 ;
      RECT 56.153 2.185 56.239 2.341 ;
      RECT 56.067 2.183 56.153 2.341 ;
      RECT 55.981 2.182 56.067 2.341 ;
      RECT 55.895 2.18 55.981 2.34 ;
      RECT 55.871 2.178 55.895 2.34 ;
      RECT 55.785 2.171 55.871 2.34 ;
      RECT 55.756 2.163 55.785 2.34 ;
      RECT 55.67 2.155 55.756 2.34 ;
      RECT 55.39 2.152 55.4 2.35 ;
      RECT 56.895 3.115 56.9 3.465 ;
      RECT 56.665 3.205 56.805 3.465 ;
      RECT 57.14 2.89 57.185 3.1 ;
      RECT 57.195 2.901 57.205 3.095 ;
      RECT 57.185 2.893 57.195 3.1 ;
      RECT 57.12 2.89 57.14 3.105 ;
      RECT 57.09 2.89 57.12 3.128 ;
      RECT 57.08 2.89 57.09 3.153 ;
      RECT 57.075 2.89 57.08 3.163 ;
      RECT 57.02 2.89 57.075 3.203 ;
      RECT 57.015 2.89 57.02 3.243 ;
      RECT 57.01 2.892 57.015 3.248 ;
      RECT 56.995 2.902 57.01 3.259 ;
      RECT 56.95 2.96 56.995 3.295 ;
      RECT 56.94 3.015 56.95 3.329 ;
      RECT 56.925 3.042 56.94 3.345 ;
      RECT 56.915 3.069 56.925 3.465 ;
      RECT 56.9 3.092 56.915 3.465 ;
      RECT 56.89 3.132 56.895 3.465 ;
      RECT 56.885 3.142 56.89 3.465 ;
      RECT 56.88 3.157 56.885 3.465 ;
      RECT 56.87 3.162 56.88 3.465 ;
      RECT 56.805 3.185 56.87 3.465 ;
      RECT 56.305 2.68 56.495 2.89 ;
      RECT 54.88 2.605 55.14 2.865 ;
      RECT 55.23 2.6 55.325 2.81 ;
      RECT 55.205 2.615 55.215 2.81 ;
      RECT 56.495 2.687 56.505 2.885 ;
      RECT 56.295 2.687 56.305 2.885 ;
      RECT 56.28 2.702 56.295 2.875 ;
      RECT 56.275 2.71 56.28 2.868 ;
      RECT 56.265 2.713 56.275 2.865 ;
      RECT 56.23 2.712 56.265 2.863 ;
      RECT 56.201 2.708 56.23 2.86 ;
      RECT 56.115 2.703 56.201 2.857 ;
      RECT 56.055 2.697 56.115 2.853 ;
      RECT 56.026 2.693 56.055 2.85 ;
      RECT 55.94 2.685 56.026 2.847 ;
      RECT 55.931 2.679 55.94 2.845 ;
      RECT 55.845 2.674 55.931 2.843 ;
      RECT 55.822 2.669 55.845 2.84 ;
      RECT 55.736 2.663 55.822 2.837 ;
      RECT 55.65 2.654 55.736 2.832 ;
      RECT 55.64 2.649 55.65 2.83 ;
      RECT 55.621 2.648 55.64 2.829 ;
      RECT 55.535 2.643 55.621 2.825 ;
      RECT 55.515 2.638 55.535 2.821 ;
      RECT 55.455 2.633 55.515 2.818 ;
      RECT 55.43 2.623 55.455 2.816 ;
      RECT 55.425 2.616 55.43 2.815 ;
      RECT 55.415 2.607 55.425 2.814 ;
      RECT 55.411 2.6 55.415 2.814 ;
      RECT 55.325 2.6 55.411 2.812 ;
      RECT 55.215 2.607 55.23 2.81 ;
      RECT 55.2 2.617 55.205 2.81 ;
      RECT 55.18 2.62 55.2 2.807 ;
      RECT 55.15 2.62 55.18 2.803 ;
      RECT 55.14 2.62 55.15 2.803 ;
      RECT 56.055 3.115 56.315 3.375 ;
      RECT 55.985 3.125 56.315 3.335 ;
      RECT 55.975 3.132 56.315 3.33 ;
      RECT 55.395 3.12 55.655 3.38 ;
      RECT 55.395 3.16 55.76 3.37 ;
      RECT 55.395 3.162 55.765 3.369 ;
      RECT 55.395 3.17 55.77 3.366 ;
      RECT 54.32 2.245 54.42 3.77 ;
      RECT 54.51 3.385 54.56 3.645 ;
      RECT 54.505 2.258 54.51 2.445 ;
      RECT 54.5 3.366 54.51 3.645 ;
      RECT 54.5 2.255 54.505 2.453 ;
      RECT 54.485 2.249 54.5 2.46 ;
      RECT 54.495 3.354 54.5 3.728 ;
      RECT 54.485 3.342 54.495 3.765 ;
      RECT 54.475 2.245 54.485 2.467 ;
      RECT 54.475 3.327 54.485 3.77 ;
      RECT 54.47 2.245 54.475 2.475 ;
      RECT 54.45 3.297 54.475 3.77 ;
      RECT 54.43 2.245 54.47 2.523 ;
      RECT 54.44 3.257 54.45 3.77 ;
      RECT 54.43 3.212 54.44 3.77 ;
      RECT 54.425 2.245 54.43 2.593 ;
      RECT 54.425 3.17 54.43 3.77 ;
      RECT 54.42 2.245 54.425 3.07 ;
      RECT 54.42 3.152 54.425 3.77 ;
      RECT 54.31 2.248 54.32 3.77 ;
      RECT 54.295 2.255 54.31 3.766 ;
      RECT 54.29 2.265 54.295 3.761 ;
      RECT 54.285 2.465 54.29 3.653 ;
      RECT 54.28 2.55 54.285 3.205 ;
      RECT 53.165 2.365 53.455 2.595 ;
      RECT 53.225 0.885 53.395 2.595 ;
      RECT 53.225 0.885 53.4 1.455 ;
      RECT 53.195 1.1 53.545 1.45 ;
      RECT 53.165 0.885 53.455 1.115 ;
      RECT 53.165 7.765 53.455 7.995 ;
      RECT 53.225 6.285 53.395 7.995 ;
      RECT 53.165 6.285 53.455 6.515 ;
      RECT 52.755 2.735 53.085 2.965 ;
      RECT 52.755 2.765 53.255 2.935 ;
      RECT 52.755 2.395 52.945 2.965 ;
      RECT 52.175 2.365 52.465 2.595 ;
      RECT 52.175 2.395 52.945 2.565 ;
      RECT 52.235 0.885 52.405 2.595 ;
      RECT 52.175 0.885 52.465 1.115 ;
      RECT 52.175 7.765 52.465 7.995 ;
      RECT 52.235 6.285 52.405 7.995 ;
      RECT 52.175 6.285 52.465 6.515 ;
      RECT 52.175 6.325 53.025 6.485 ;
      RECT 52.855 5.915 53.025 6.485 ;
      RECT 52.175 6.32 52.565 6.485 ;
      RECT 52.795 5.915 53.085 6.145 ;
      RECT 52.795 5.945 53.255 6.115 ;
      RECT 51.805 2.735 52.095 2.965 ;
      RECT 51.805 2.765 52.265 2.935 ;
      RECT 51.865 1.655 52.03 2.965 ;
      RECT 50.38 1.625 50.67 1.855 ;
      RECT 50.38 1.655 52.03 1.825 ;
      RECT 50.44 0.885 50.61 1.855 ;
      RECT 50.38 0.885 50.67 1.115 ;
      RECT 50.38 7.765 50.67 7.995 ;
      RECT 50.44 7.025 50.61 7.995 ;
      RECT 50.44 7.12 52.03 7.29 ;
      RECT 51.86 5.915 52.03 7.29 ;
      RECT 50.38 7.025 50.67 7.255 ;
      RECT 51.805 5.915 52.095 6.145 ;
      RECT 51.805 5.945 52.265 6.115 ;
      RECT 50.81 1.965 51.16 2.315 ;
      RECT 50.64 2.025 51.16 2.195 ;
      RECT 50.835 6.655 51.16 6.98 ;
      RECT 50.81 6.655 51.16 6.885 ;
      RECT 50.64 6.685 51.16 6.855 ;
      RECT 48.415 3.43 48.765 3.78 ;
      RECT 48.505 2.395 48.675 3.78 ;
      RECT 50.035 2.365 50.355 2.685 ;
      RECT 50.005 2.365 50.355 2.595 ;
      RECT 48.505 2.395 50.355 2.565 ;
      RECT 50.035 6.28 50.355 6.605 ;
      RECT 50.005 6.285 50.355 6.515 ;
      RECT 49.835 6.315 50.355 6.485 ;
      RECT 48.99 2.705 49.34 3.055 ;
      RECT 48.99 2.765 49.47 2.935 ;
      RECT 48.98 5.84 49.33 6.19 ;
      RECT 48.98 5.945 49.47 6.115 ;
      RECT 45.815 3.665 45.855 3.925 ;
      RECT 45.855 3.645 45.86 3.655 ;
      RECT 47.195 2.735 47.35 3.055 ;
      RECT 47.115 2.735 47.195 3.22 ;
      RECT 47.105 2.735 47.115 3.363 ;
      RECT 47.08 2.735 47.105 3.41 ;
      RECT 47.055 2.735 47.08 3.488 ;
      RECT 47.035 2.735 47.055 3.558 ;
      RECT 47.03 2.735 47.035 3.588 ;
      RECT 47.01 2.885 47.03 3.6 ;
      RECT 47 2.885 47.01 3.618 ;
      RECT 46.99 2.887 47 3.626 ;
      RECT 46.985 2.892 46.99 3.083 ;
      RECT 46.985 3.092 46.99 3.627 ;
      RECT 46.98 3.137 46.985 3.628 ;
      RECT 46.97 3.202 46.98 3.629 ;
      RECT 46.96 3.297 46.97 3.631 ;
      RECT 46.955 3.35 46.96 3.633 ;
      RECT 46.95 3.37 46.955 3.634 ;
      RECT 46.895 3.395 46.95 3.64 ;
      RECT 46.855 3.43 46.895 3.649 ;
      RECT 46.845 3.447 46.855 3.654 ;
      RECT 46.836 3.453 46.845 3.656 ;
      RECT 46.75 3.491 46.836 3.667 ;
      RECT 46.745 3.53 46.75 3.677 ;
      RECT 46.67 3.537 46.745 3.687 ;
      RECT 46.65 3.547 46.67 3.698 ;
      RECT 46.62 3.554 46.65 3.706 ;
      RECT 46.595 3.561 46.62 3.713 ;
      RECT 46.571 3.567 46.595 3.718 ;
      RECT 46.485 3.58 46.571 3.73 ;
      RECT 46.407 3.587 46.485 3.748 ;
      RECT 46.321 3.582 46.407 3.766 ;
      RECT 46.235 3.577 46.321 3.786 ;
      RECT 46.155 3.571 46.235 3.803 ;
      RECT 46.09 3.567 46.155 3.832 ;
      RECT 46.085 3.281 46.09 3.305 ;
      RECT 46.075 3.557 46.09 3.86 ;
      RECT 46.08 3.275 46.085 3.345 ;
      RECT 46.075 3.269 46.08 3.415 ;
      RECT 46.07 3.263 46.075 3.493 ;
      RECT 46.07 3.54 46.075 3.925 ;
      RECT 46.062 3.26 46.07 3.925 ;
      RECT 45.976 3.258 46.062 3.925 ;
      RECT 45.89 3.256 45.976 3.925 ;
      RECT 45.88 3.257 45.89 3.925 ;
      RECT 45.875 3.262 45.88 3.925 ;
      RECT 45.865 3.275 45.875 3.925 ;
      RECT 45.86 3.297 45.865 3.925 ;
      RECT 45.855 3.657 45.86 3.925 ;
      RECT 46.485 3.125 46.49 3.345 ;
      RECT 46.99 2.16 47.025 2.42 ;
      RECT 46.975 2.16 46.99 2.428 ;
      RECT 46.946 2.16 46.975 2.45 ;
      RECT 46.86 2.16 46.946 2.51 ;
      RECT 46.84 2.16 46.86 2.575 ;
      RECT 46.78 2.16 46.84 2.74 ;
      RECT 46.775 2.16 46.78 2.888 ;
      RECT 46.77 2.16 46.775 2.9 ;
      RECT 46.765 2.16 46.77 2.926 ;
      RECT 46.735 2.346 46.765 3.006 ;
      RECT 46.73 2.394 46.735 3.095 ;
      RECT 46.725 2.408 46.73 3.11 ;
      RECT 46.72 2.427 46.725 3.14 ;
      RECT 46.715 2.442 46.72 3.156 ;
      RECT 46.71 2.457 46.715 3.178 ;
      RECT 46.705 2.477 46.71 3.2 ;
      RECT 46.695 2.497 46.705 3.233 ;
      RECT 46.68 2.539 46.695 3.295 ;
      RECT 46.675 2.57 46.68 3.335 ;
      RECT 46.67 2.582 46.675 3.34 ;
      RECT 46.665 2.594 46.67 3.345 ;
      RECT 46.66 2.607 46.665 3.345 ;
      RECT 46.655 2.625 46.66 3.345 ;
      RECT 46.65 2.645 46.655 3.345 ;
      RECT 46.645 2.657 46.65 3.345 ;
      RECT 46.64 2.67 46.645 3.345 ;
      RECT 46.62 2.705 46.64 3.345 ;
      RECT 46.57 2.807 46.62 3.345 ;
      RECT 46.565 2.892 46.57 3.345 ;
      RECT 46.56 2.9 46.565 3.345 ;
      RECT 46.555 2.917 46.56 3.345 ;
      RECT 46.55 2.932 46.555 3.345 ;
      RECT 46.515 2.997 46.55 3.345 ;
      RECT 46.5 3.062 46.515 3.345 ;
      RECT 46.495 3.092 46.5 3.345 ;
      RECT 46.49 3.117 46.495 3.345 ;
      RECT 46.475 3.127 46.485 3.345 ;
      RECT 46.46 3.14 46.475 3.338 ;
      RECT 46.205 2.73 46.275 2.94 ;
      RECT 45.995 2.707 46 2.9 ;
      RECT 43.45 2.635 43.71 2.895 ;
      RECT 46.285 2.917 46.29 2.92 ;
      RECT 46.275 2.735 46.285 2.935 ;
      RECT 46.176 2.728 46.205 2.94 ;
      RECT 46.09 2.72 46.176 2.94 ;
      RECT 46.075 2.714 46.09 2.938 ;
      RECT 46.055 2.713 46.075 2.925 ;
      RECT 46.05 2.712 46.055 2.908 ;
      RECT 46 2.709 46.05 2.903 ;
      RECT 45.97 2.706 45.995 2.898 ;
      RECT 45.95 2.704 45.97 2.893 ;
      RECT 45.935 2.702 45.95 2.89 ;
      RECT 45.905 2.7 45.935 2.888 ;
      RECT 45.84 2.696 45.905 2.88 ;
      RECT 45.81 2.691 45.84 2.875 ;
      RECT 45.79 2.689 45.81 2.873 ;
      RECT 45.76 2.686 45.79 2.868 ;
      RECT 45.7 2.682 45.76 2.86 ;
      RECT 45.695 2.679 45.7 2.855 ;
      RECT 45.625 2.677 45.695 2.85 ;
      RECT 45.596 2.673 45.625 2.843 ;
      RECT 45.51 2.668 45.596 2.835 ;
      RECT 45.476 2.663 45.51 2.827 ;
      RECT 45.39 2.655 45.476 2.819 ;
      RECT 45.351 2.648 45.39 2.811 ;
      RECT 45.265 2.643 45.351 2.803 ;
      RECT 45.2 2.637 45.265 2.793 ;
      RECT 45.18 2.632 45.2 2.788 ;
      RECT 45.171 2.629 45.18 2.787 ;
      RECT 45.085 2.625 45.171 2.781 ;
      RECT 45.045 2.621 45.085 2.773 ;
      RECT 45.025 2.617 45.045 2.771 ;
      RECT 44.965 2.617 45.025 2.768 ;
      RECT 44.945 2.62 44.965 2.766 ;
      RECT 44.924 2.62 44.945 2.766 ;
      RECT 44.838 2.622 44.924 2.77 ;
      RECT 44.752 2.624 44.838 2.776 ;
      RECT 44.666 2.626 44.752 2.783 ;
      RECT 44.58 2.629 44.666 2.789 ;
      RECT 44.546 2.63 44.58 2.794 ;
      RECT 44.46 2.633 44.546 2.799 ;
      RECT 44.431 2.64 44.46 2.804 ;
      RECT 44.345 2.64 44.431 2.809 ;
      RECT 44.312 2.64 44.345 2.814 ;
      RECT 44.226 2.642 44.312 2.819 ;
      RECT 44.14 2.644 44.226 2.826 ;
      RECT 44.076 2.646 44.14 2.832 ;
      RECT 43.99 2.648 44.076 2.838 ;
      RECT 43.987 2.65 43.99 2.841 ;
      RECT 43.901 2.651 43.987 2.845 ;
      RECT 43.815 2.654 43.901 2.852 ;
      RECT 43.796 2.656 43.815 2.856 ;
      RECT 43.71 2.658 43.796 2.861 ;
      RECT 43.44 2.67 43.45 2.865 ;
      RECT 45.675 2.25 45.86 2.46 ;
      RECT 45.67 2.251 45.865 2.458 ;
      RECT 45.665 2.256 45.875 2.453 ;
      RECT 45.66 2.232 45.665 2.45 ;
      RECT 45.63 2.229 45.66 2.443 ;
      RECT 45.625 2.225 45.63 2.434 ;
      RECT 45.59 2.256 45.875 2.429 ;
      RECT 45.365 2.165 45.625 2.425 ;
      RECT 45.665 2.234 45.67 2.453 ;
      RECT 45.67 2.235 45.675 2.458 ;
      RECT 45.365 2.247 45.745 2.425 ;
      RECT 45.365 2.245 45.73 2.425 ;
      RECT 45.365 2.24 45.72 2.425 ;
      RECT 45.32 3.155 45.37 3.44 ;
      RECT 45.265 3.125 45.27 3.44 ;
      RECT 45.235 3.105 45.24 3.44 ;
      RECT 45.385 3.155 45.445 3.415 ;
      RECT 45.38 3.155 45.385 3.423 ;
      RECT 45.37 3.155 45.38 3.435 ;
      RECT 45.285 3.145 45.32 3.44 ;
      RECT 45.28 3.132 45.285 3.44 ;
      RECT 45.27 3.127 45.28 3.44 ;
      RECT 45.25 3.117 45.265 3.44 ;
      RECT 45.24 3.11 45.25 3.44 ;
      RECT 45.23 3.102 45.235 3.44 ;
      RECT 45.2 3.092 45.23 3.44 ;
      RECT 45.185 3.08 45.2 3.44 ;
      RECT 45.17 3.07 45.185 3.435 ;
      RECT 45.15 3.06 45.17 3.41 ;
      RECT 45.14 3.052 45.15 3.387 ;
      RECT 45.11 3.035 45.14 3.377 ;
      RECT 45.105 3.012 45.11 3.368 ;
      RECT 45.1 2.999 45.105 3.366 ;
      RECT 45.085 2.975 45.1 3.36 ;
      RECT 45.08 2.951 45.085 3.354 ;
      RECT 45.07 2.94 45.08 3.349 ;
      RECT 45.065 2.93 45.07 3.345 ;
      RECT 45.06 2.922 45.065 3.342 ;
      RECT 45.05 2.917 45.06 3.338 ;
      RECT 45.045 2.912 45.05 3.334 ;
      RECT 44.96 2.91 45.045 3.309 ;
      RECT 44.93 2.91 44.96 3.275 ;
      RECT 44.915 2.91 44.93 3.258 ;
      RECT 44.86 2.91 44.915 3.203 ;
      RECT 44.855 2.915 44.86 3.152 ;
      RECT 44.845 2.92 44.855 3.142 ;
      RECT 44.84 2.93 44.845 3.128 ;
      RECT 44.79 3.67 45.05 3.93 ;
      RECT 44.71 3.685 45.05 3.906 ;
      RECT 44.69 3.685 45.05 3.901 ;
      RECT 44.666 3.685 45.05 3.899 ;
      RECT 44.58 3.685 45.05 3.894 ;
      RECT 44.43 3.625 44.69 3.89 ;
      RECT 44.385 3.685 45.05 3.885 ;
      RECT 44.38 3.692 45.05 3.88 ;
      RECT 44.395 3.68 44.71 3.89 ;
      RECT 44.285 2.115 44.545 2.375 ;
      RECT 44.285 2.172 44.55 2.368 ;
      RECT 44.285 2.202 44.555 2.3 ;
      RECT 44.345 2.633 44.46 2.635 ;
      RECT 44.431 2.63 44.46 2.635 ;
      RECT 43.455 3.634 43.48 3.874 ;
      RECT 43.44 3.637 43.53 3.868 ;
      RECT 43.435 3.642 43.616 3.863 ;
      RECT 43.43 3.65 43.68 3.861 ;
      RECT 43.43 3.65 43.69 3.86 ;
      RECT 43.425 3.657 43.7 3.853 ;
      RECT 43.425 3.657 43.786 3.842 ;
      RECT 43.42 3.692 43.786 3.838 ;
      RECT 43.42 3.692 43.795 3.827 ;
      RECT 43.7 3.565 43.96 3.825 ;
      RECT 43.41 3.742 43.96 3.823 ;
      RECT 43.68 3.61 43.7 3.858 ;
      RECT 43.616 3.613 43.68 3.862 ;
      RECT 43.53 3.618 43.616 3.867 ;
      RECT 43.46 3.629 43.96 3.825 ;
      RECT 43.48 3.623 43.53 3.872 ;
      RECT 43.605 2.1 43.615 2.362 ;
      RECT 43.595 2.157 43.605 2.365 ;
      RECT 43.57 2.162 43.595 2.371 ;
      RECT 43.545 2.166 43.57 2.383 ;
      RECT 43.535 2.169 43.545 2.393 ;
      RECT 43.53 2.17 43.535 2.398 ;
      RECT 43.525 2.171 43.53 2.403 ;
      RECT 43.52 2.172 43.525 2.405 ;
      RECT 43.495 2.175 43.52 2.408 ;
      RECT 43.465 2.181 43.495 2.411 ;
      RECT 43.4 2.192 43.465 2.414 ;
      RECT 43.355 2.2 43.4 2.418 ;
      RECT 43.34 2.2 43.355 2.426 ;
      RECT 43.335 2.201 43.34 2.433 ;
      RECT 43.33 2.203 43.335 2.436 ;
      RECT 43.325 2.207 43.33 2.439 ;
      RECT 43.315 2.215 43.325 2.443 ;
      RECT 43.31 2.228 43.315 2.448 ;
      RECT 43.305 2.236 43.31 2.45 ;
      RECT 43.3 2.242 43.305 2.45 ;
      RECT 43.295 2.246 43.3 2.453 ;
      RECT 43.29 2.248 43.295 2.456 ;
      RECT 43.285 2.251 43.29 2.459 ;
      RECT 43.275 2.256 43.285 2.463 ;
      RECT 43.27 2.262 43.275 2.468 ;
      RECT 43.26 2.268 43.27 2.472 ;
      RECT 43.245 2.275 43.26 2.478 ;
      RECT 43.216 2.289 43.245 2.488 ;
      RECT 43.13 2.324 43.216 2.52 ;
      RECT 43.11 2.357 43.13 2.549 ;
      RECT 43.09 2.37 43.11 2.56 ;
      RECT 43.07 2.382 43.09 2.571 ;
      RECT 43.02 2.404 43.07 2.591 ;
      RECT 43.005 2.422 43.02 2.608 ;
      RECT 43 2.428 43.005 2.611 ;
      RECT 42.995 2.432 43 2.614 ;
      RECT 42.99 2.436 42.995 2.618 ;
      RECT 42.985 2.438 42.99 2.621 ;
      RECT 42.975 2.445 42.985 2.624 ;
      RECT 42.97 2.45 42.975 2.628 ;
      RECT 42.965 2.452 42.97 2.631 ;
      RECT 42.96 2.456 42.965 2.634 ;
      RECT 42.955 2.458 42.96 2.638 ;
      RECT 42.94 2.463 42.955 2.643 ;
      RECT 42.935 2.468 42.94 2.646 ;
      RECT 42.93 2.476 42.935 2.649 ;
      RECT 42.925 2.478 42.93 2.652 ;
      RECT 42.92 2.48 42.925 2.655 ;
      RECT 42.91 2.482 42.92 2.661 ;
      RECT 42.875 2.496 42.91 2.673 ;
      RECT 42.865 2.511 42.875 2.683 ;
      RECT 42.79 2.54 42.865 2.707 ;
      RECT 42.785 2.565 42.79 2.73 ;
      RECT 42.77 2.569 42.785 2.736 ;
      RECT 42.76 2.577 42.77 2.741 ;
      RECT 42.73 2.59 42.76 2.745 ;
      RECT 42.72 2.605 42.73 2.75 ;
      RECT 42.71 2.61 42.72 2.753 ;
      RECT 42.705 2.612 42.71 2.755 ;
      RECT 42.69 2.615 42.705 2.758 ;
      RECT 42.685 2.617 42.69 2.761 ;
      RECT 42.665 2.622 42.685 2.765 ;
      RECT 42.635 2.627 42.665 2.773 ;
      RECT 42.61 2.634 42.635 2.781 ;
      RECT 42.605 2.639 42.61 2.786 ;
      RECT 42.575 2.642 42.605 2.79 ;
      RECT 42.535 2.645 42.575 2.8 ;
      RECT 42.5 2.642 42.535 2.812 ;
      RECT 42.49 2.638 42.5 2.819 ;
      RECT 42.465 2.634 42.49 2.825 ;
      RECT 42.46 2.63 42.465 2.83 ;
      RECT 42.42 2.627 42.46 2.83 ;
      RECT 42.405 2.612 42.42 2.831 ;
      RECT 42.382 2.6 42.405 2.831 ;
      RECT 42.296 2.6 42.382 2.832 ;
      RECT 42.21 2.6 42.296 2.834 ;
      RECT 42.19 2.6 42.21 2.831 ;
      RECT 42.185 2.605 42.19 2.826 ;
      RECT 42.18 2.61 42.185 2.824 ;
      RECT 42.17 2.62 42.18 2.822 ;
      RECT 42.165 2.626 42.17 2.815 ;
      RECT 42.16 2.628 42.165 2.8 ;
      RECT 42.155 2.632 42.16 2.79 ;
      RECT 43.615 2.1 43.865 2.36 ;
      RECT 41.34 3.635 41.6 3.895 ;
      RECT 43.635 3.125 43.64 3.335 ;
      RECT 43.64 3.13 43.65 3.33 ;
      RECT 43.59 3.125 43.635 3.35 ;
      RECT 43.58 3.125 43.59 3.37 ;
      RECT 43.561 3.125 43.58 3.375 ;
      RECT 43.475 3.125 43.561 3.372 ;
      RECT 43.445 3.127 43.475 3.37 ;
      RECT 43.39 3.137 43.445 3.368 ;
      RECT 43.325 3.151 43.39 3.366 ;
      RECT 43.32 3.159 43.325 3.365 ;
      RECT 43.305 3.162 43.32 3.363 ;
      RECT 43.24 3.172 43.305 3.359 ;
      RECT 43.192 3.186 43.24 3.36 ;
      RECT 43.106 3.203 43.192 3.374 ;
      RECT 43.02 3.224 43.106 3.391 ;
      RECT 43 3.237 43.02 3.401 ;
      RECT 42.955 3.245 43 3.408 ;
      RECT 42.92 3.253 42.955 3.416 ;
      RECT 42.886 3.261 42.92 3.424 ;
      RECT 42.8 3.275 42.886 3.436 ;
      RECT 42.765 3.292 42.8 3.448 ;
      RECT 42.756 3.301 42.765 3.452 ;
      RECT 42.67 3.319 42.756 3.469 ;
      RECT 42.611 3.346 42.67 3.496 ;
      RECT 42.525 3.373 42.611 3.524 ;
      RECT 42.505 3.395 42.525 3.544 ;
      RECT 42.445 3.41 42.505 3.56 ;
      RECT 42.435 3.422 42.445 3.573 ;
      RECT 42.43 3.427 42.435 3.576 ;
      RECT 42.42 3.43 42.43 3.579 ;
      RECT 42.415 3.432 42.42 3.582 ;
      RECT 42.385 3.44 42.415 3.589 ;
      RECT 42.37 3.447 42.385 3.597 ;
      RECT 42.36 3.452 42.37 3.601 ;
      RECT 42.355 3.455 42.36 3.604 ;
      RECT 42.345 3.457 42.355 3.607 ;
      RECT 42.31 3.467 42.345 3.616 ;
      RECT 42.235 3.49 42.31 3.638 ;
      RECT 42.215 3.508 42.235 3.656 ;
      RECT 42.185 3.515 42.215 3.666 ;
      RECT 42.165 3.523 42.185 3.676 ;
      RECT 42.155 3.529 42.165 3.683 ;
      RECT 42.136 3.534 42.155 3.689 ;
      RECT 42.05 3.554 42.136 3.709 ;
      RECT 42.035 3.574 42.05 3.728 ;
      RECT 41.99 3.586 42.035 3.739 ;
      RECT 41.925 3.607 41.99 3.762 ;
      RECT 41.885 3.627 41.925 3.783 ;
      RECT 41.875 3.637 41.885 3.793 ;
      RECT 41.825 3.649 41.875 3.804 ;
      RECT 41.805 3.665 41.825 3.816 ;
      RECT 41.775 3.675 41.805 3.822 ;
      RECT 41.765 3.68 41.775 3.824 ;
      RECT 41.696 3.681 41.765 3.83 ;
      RECT 41.61 3.683 41.696 3.84 ;
      RECT 41.6 3.684 41.61 3.845 ;
      RECT 42.87 3.71 43.06 3.92 ;
      RECT 42.86 3.715 43.07 3.913 ;
      RECT 42.845 3.715 43.07 3.878 ;
      RECT 42.765 3.6 43.025 3.86 ;
      RECT 41.68 3.13 41.865 3.425 ;
      RECT 41.67 3.13 41.865 3.423 ;
      RECT 41.655 3.13 41.87 3.418 ;
      RECT 41.655 3.13 41.875 3.415 ;
      RECT 41.65 3.13 41.875 3.413 ;
      RECT 41.645 3.385 41.875 3.403 ;
      RECT 41.65 3.13 41.91 3.39 ;
      RECT 41.61 2.165 41.87 2.425 ;
      RECT 41.42 2.09 41.506 2.423 ;
      RECT 41.395 2.094 41.55 2.419 ;
      RECT 41.506 2.086 41.55 2.419 ;
      RECT 41.506 2.087 41.555 2.418 ;
      RECT 41.42 2.092 41.57 2.417 ;
      RECT 41.395 2.1 41.61 2.416 ;
      RECT 41.39 2.095 41.57 2.411 ;
      RECT 41.38 2.11 41.61 2.318 ;
      RECT 41.38 2.162 41.81 2.318 ;
      RECT 41.38 2.155 41.79 2.318 ;
      RECT 41.38 2.142 41.76 2.318 ;
      RECT 41.38 2.13 41.7 2.318 ;
      RECT 41.38 2.115 41.675 2.318 ;
      RECT 40.58 2.745 40.715 3.04 ;
      RECT 40.84 2.768 40.845 2.955 ;
      RECT 41.56 2.665 41.705 2.9 ;
      RECT 41.72 2.665 41.725 2.89 ;
      RECT 41.755 2.676 41.76 2.87 ;
      RECT 41.75 2.668 41.755 2.875 ;
      RECT 41.73 2.665 41.75 2.88 ;
      RECT 41.725 2.665 41.73 2.888 ;
      RECT 41.715 2.665 41.72 2.893 ;
      RECT 41.705 2.665 41.715 2.898 ;
      RECT 41.535 2.667 41.56 2.9 ;
      RECT 41.485 2.674 41.535 2.9 ;
      RECT 41.48 2.679 41.485 2.9 ;
      RECT 41.441 2.684 41.48 2.901 ;
      RECT 41.355 2.696 41.441 2.902 ;
      RECT 41.346 2.706 41.355 2.902 ;
      RECT 41.26 2.715 41.346 2.904 ;
      RECT 41.236 2.725 41.26 2.906 ;
      RECT 41.15 2.736 41.236 2.907 ;
      RECT 41.12 2.747 41.15 2.909 ;
      RECT 41.09 2.752 41.12 2.911 ;
      RECT 41.065 2.758 41.09 2.914 ;
      RECT 41.05 2.763 41.065 2.915 ;
      RECT 41.005 2.769 41.05 2.915 ;
      RECT 41 2.774 41.005 2.916 ;
      RECT 40.98 2.774 41 2.918 ;
      RECT 40.96 2.772 40.98 2.923 ;
      RECT 40.925 2.771 40.96 2.93 ;
      RECT 40.895 2.77 40.925 2.94 ;
      RECT 40.845 2.769 40.895 2.95 ;
      RECT 40.755 2.766 40.84 3.04 ;
      RECT 40.73 2.76 40.755 3.04 ;
      RECT 40.715 2.75 40.73 3.04 ;
      RECT 40.53 2.745 40.58 2.96 ;
      RECT 40.52 2.75 40.53 2.95 ;
      RECT 40.76 3.225 41.02 3.485 ;
      RECT 40.76 3.225 41.05 3.378 ;
      RECT 40.76 3.225 41.085 3.363 ;
      RECT 41.015 3.145 41.205 3.355 ;
      RECT 41.005 3.15 41.215 3.348 ;
      RECT 40.97 3.22 41.215 3.348 ;
      RECT 41 3.162 41.02 3.485 ;
      RECT 40.985 3.21 41.215 3.348 ;
      RECT 40.99 3.182 41.02 3.485 ;
      RECT 40.07 2.25 40.14 3.355 ;
      RECT 40.805 2.355 41.065 2.615 ;
      RECT 40.385 2.401 40.4 2.61 ;
      RECT 40.721 2.414 40.805 2.565 ;
      RECT 40.635 2.411 40.721 2.565 ;
      RECT 40.596 2.409 40.635 2.565 ;
      RECT 40.51 2.407 40.596 2.565 ;
      RECT 40.45 2.405 40.51 2.576 ;
      RECT 40.415 2.403 40.45 2.594 ;
      RECT 40.4 2.401 40.415 2.605 ;
      RECT 40.37 2.401 40.385 2.618 ;
      RECT 40.36 2.401 40.37 2.623 ;
      RECT 40.335 2.4 40.36 2.628 ;
      RECT 40.32 2.395 40.335 2.634 ;
      RECT 40.315 2.388 40.32 2.639 ;
      RECT 40.29 2.379 40.315 2.645 ;
      RECT 40.245 2.358 40.29 2.658 ;
      RECT 40.235 2.342 40.245 2.668 ;
      RECT 40.22 2.335 40.235 2.678 ;
      RECT 40.21 2.328 40.22 2.695 ;
      RECT 40.205 2.325 40.21 2.725 ;
      RECT 40.2 2.323 40.205 2.755 ;
      RECT 40.195 2.321 40.2 2.792 ;
      RECT 40.18 2.317 40.195 2.859 ;
      RECT 40.18 3.15 40.19 3.35 ;
      RECT 40.175 2.313 40.18 2.985 ;
      RECT 40.175 3.137 40.18 3.355 ;
      RECT 40.17 2.311 40.175 3.07 ;
      RECT 40.17 3.127 40.175 3.355 ;
      RECT 40.155 2.282 40.17 3.355 ;
      RECT 40.14 2.255 40.155 3.355 ;
      RECT 40.065 2.25 40.07 2.605 ;
      RECT 40.065 2.66 40.07 3.355 ;
      RECT 40.05 2.25 40.065 2.583 ;
      RECT 40.06 2.682 40.065 3.355 ;
      RECT 40.05 2.722 40.06 3.355 ;
      RECT 40.015 2.25 40.05 2.525 ;
      RECT 40.045 2.757 40.05 3.355 ;
      RECT 40.03 2.812 40.045 3.355 ;
      RECT 40.025 2.877 40.03 3.355 ;
      RECT 40.01 2.925 40.025 3.355 ;
      RECT 39.985 2.25 40.015 2.48 ;
      RECT 40.005 2.98 40.01 3.355 ;
      RECT 39.99 3.04 40.005 3.355 ;
      RECT 39.985 3.088 39.99 3.353 ;
      RECT 39.98 2.25 39.985 2.473 ;
      RECT 39.98 3.12 39.985 3.348 ;
      RECT 39.955 2.25 39.98 2.465 ;
      RECT 39.945 2.255 39.955 2.455 ;
      RECT 40.16 3.53 40.18 3.77 ;
      RECT 39.39 3.46 39.395 3.67 ;
      RECT 40.67 3.533 40.68 3.728 ;
      RECT 40.665 3.523 40.67 3.731 ;
      RECT 40.585 3.52 40.665 3.754 ;
      RECT 40.581 3.52 40.585 3.776 ;
      RECT 40.495 3.52 40.581 3.786 ;
      RECT 40.48 3.52 40.495 3.794 ;
      RECT 40.451 3.521 40.48 3.792 ;
      RECT 40.365 3.526 40.451 3.788 ;
      RECT 40.352 3.53 40.365 3.784 ;
      RECT 40.266 3.53 40.352 3.78 ;
      RECT 40.18 3.53 40.266 3.774 ;
      RECT 40.096 3.53 40.16 3.768 ;
      RECT 40.01 3.53 40.096 3.763 ;
      RECT 39.99 3.53 40.01 3.759 ;
      RECT 39.93 3.525 39.99 3.756 ;
      RECT 39.902 3.519 39.93 3.753 ;
      RECT 39.816 3.514 39.902 3.749 ;
      RECT 39.73 3.508 39.816 3.743 ;
      RECT 39.655 3.49 39.73 3.738 ;
      RECT 39.62 3.467 39.655 3.734 ;
      RECT 39.61 3.457 39.62 3.733 ;
      RECT 39.555 3.455 39.61 3.732 ;
      RECT 39.48 3.455 39.555 3.728 ;
      RECT 39.47 3.455 39.48 3.723 ;
      RECT 39.455 3.455 39.47 3.715 ;
      RECT 39.405 3.457 39.455 3.693 ;
      RECT 39.395 3.46 39.405 3.673 ;
      RECT 39.385 3.465 39.39 3.668 ;
      RECT 39.38 3.47 39.385 3.663 ;
      RECT 39.505 2.635 39.765 2.895 ;
      RECT 39.505 2.65 39.785 2.86 ;
      RECT 39.505 2.655 39.795 2.855 ;
      RECT 37.49 2.115 37.75 2.375 ;
      RECT 37.48 2.145 37.75 2.355 ;
      RECT 39.4 2.06 39.66 2.32 ;
      RECT 39.395 2.135 39.4 2.321 ;
      RECT 39.37 2.14 39.395 2.323 ;
      RECT 39.355 2.147 39.37 2.326 ;
      RECT 39.295 2.165 39.355 2.331 ;
      RECT 39.265 2.185 39.295 2.338 ;
      RECT 39.24 2.193 39.265 2.343 ;
      RECT 39.215 2.201 39.24 2.345 ;
      RECT 39.197 2.205 39.215 2.344 ;
      RECT 39.111 2.203 39.197 2.344 ;
      RECT 39.025 2.201 39.111 2.344 ;
      RECT 38.939 2.199 39.025 2.343 ;
      RECT 38.853 2.197 38.939 2.343 ;
      RECT 38.767 2.195 38.853 2.343 ;
      RECT 38.681 2.193 38.767 2.343 ;
      RECT 38.595 2.191 38.681 2.342 ;
      RECT 38.577 2.19 38.595 2.342 ;
      RECT 38.491 2.189 38.577 2.342 ;
      RECT 38.405 2.187 38.491 2.342 ;
      RECT 38.319 2.186 38.405 2.341 ;
      RECT 38.233 2.185 38.319 2.341 ;
      RECT 38.147 2.183 38.233 2.341 ;
      RECT 38.061 2.182 38.147 2.341 ;
      RECT 37.975 2.18 38.061 2.34 ;
      RECT 37.951 2.178 37.975 2.34 ;
      RECT 37.865 2.171 37.951 2.34 ;
      RECT 37.836 2.163 37.865 2.34 ;
      RECT 37.75 2.155 37.836 2.34 ;
      RECT 37.47 2.152 37.48 2.35 ;
      RECT 38.975 3.115 38.98 3.465 ;
      RECT 38.745 3.205 38.885 3.465 ;
      RECT 39.22 2.89 39.265 3.1 ;
      RECT 39.275 2.901 39.285 3.095 ;
      RECT 39.265 2.893 39.275 3.1 ;
      RECT 39.2 2.89 39.22 3.105 ;
      RECT 39.17 2.89 39.2 3.128 ;
      RECT 39.16 2.89 39.17 3.153 ;
      RECT 39.155 2.89 39.16 3.163 ;
      RECT 39.1 2.89 39.155 3.203 ;
      RECT 39.095 2.89 39.1 3.243 ;
      RECT 39.09 2.892 39.095 3.248 ;
      RECT 39.075 2.902 39.09 3.259 ;
      RECT 39.03 2.96 39.075 3.295 ;
      RECT 39.02 3.015 39.03 3.329 ;
      RECT 39.005 3.042 39.02 3.345 ;
      RECT 38.995 3.069 39.005 3.465 ;
      RECT 38.98 3.092 38.995 3.465 ;
      RECT 38.97 3.132 38.975 3.465 ;
      RECT 38.965 3.142 38.97 3.465 ;
      RECT 38.96 3.157 38.965 3.465 ;
      RECT 38.95 3.162 38.96 3.465 ;
      RECT 38.885 3.185 38.95 3.465 ;
      RECT 38.385 2.68 38.575 2.89 ;
      RECT 36.96 2.605 37.22 2.865 ;
      RECT 37.31 2.6 37.405 2.81 ;
      RECT 37.285 2.615 37.295 2.81 ;
      RECT 38.575 2.687 38.585 2.885 ;
      RECT 38.375 2.687 38.385 2.885 ;
      RECT 38.36 2.702 38.375 2.875 ;
      RECT 38.355 2.71 38.36 2.868 ;
      RECT 38.345 2.713 38.355 2.865 ;
      RECT 38.31 2.712 38.345 2.863 ;
      RECT 38.281 2.708 38.31 2.86 ;
      RECT 38.195 2.703 38.281 2.857 ;
      RECT 38.135 2.697 38.195 2.853 ;
      RECT 38.106 2.693 38.135 2.85 ;
      RECT 38.02 2.685 38.106 2.847 ;
      RECT 38.011 2.679 38.02 2.845 ;
      RECT 37.925 2.674 38.011 2.843 ;
      RECT 37.902 2.669 37.925 2.84 ;
      RECT 37.816 2.663 37.902 2.837 ;
      RECT 37.73 2.654 37.816 2.832 ;
      RECT 37.72 2.649 37.73 2.83 ;
      RECT 37.701 2.648 37.72 2.829 ;
      RECT 37.615 2.643 37.701 2.825 ;
      RECT 37.595 2.638 37.615 2.821 ;
      RECT 37.535 2.633 37.595 2.818 ;
      RECT 37.51 2.623 37.535 2.816 ;
      RECT 37.505 2.616 37.51 2.815 ;
      RECT 37.495 2.607 37.505 2.814 ;
      RECT 37.491 2.6 37.495 2.814 ;
      RECT 37.405 2.6 37.491 2.812 ;
      RECT 37.295 2.607 37.31 2.81 ;
      RECT 37.28 2.617 37.285 2.81 ;
      RECT 37.26 2.62 37.28 2.807 ;
      RECT 37.23 2.62 37.26 2.803 ;
      RECT 37.22 2.62 37.23 2.803 ;
      RECT 38.135 3.115 38.395 3.375 ;
      RECT 38.065 3.125 38.395 3.335 ;
      RECT 38.055 3.132 38.395 3.33 ;
      RECT 37.475 3.12 37.735 3.38 ;
      RECT 37.475 3.16 37.84 3.37 ;
      RECT 37.475 3.162 37.845 3.369 ;
      RECT 37.475 3.17 37.85 3.366 ;
      RECT 36.4 2.245 36.5 3.77 ;
      RECT 36.59 3.385 36.64 3.645 ;
      RECT 36.585 2.258 36.59 2.445 ;
      RECT 36.58 3.366 36.59 3.645 ;
      RECT 36.58 2.255 36.585 2.453 ;
      RECT 36.565 2.249 36.58 2.46 ;
      RECT 36.575 3.354 36.58 3.728 ;
      RECT 36.565 3.342 36.575 3.765 ;
      RECT 36.555 2.245 36.565 2.467 ;
      RECT 36.555 3.327 36.565 3.77 ;
      RECT 36.55 2.245 36.555 2.475 ;
      RECT 36.53 3.297 36.555 3.77 ;
      RECT 36.51 2.245 36.55 2.523 ;
      RECT 36.52 3.257 36.53 3.77 ;
      RECT 36.51 3.212 36.52 3.77 ;
      RECT 36.505 2.245 36.51 2.593 ;
      RECT 36.505 3.17 36.51 3.77 ;
      RECT 36.5 2.245 36.505 3.07 ;
      RECT 36.5 3.152 36.505 3.77 ;
      RECT 36.39 2.248 36.4 3.77 ;
      RECT 36.375 2.255 36.39 3.766 ;
      RECT 36.37 2.265 36.375 3.761 ;
      RECT 36.365 2.465 36.37 3.653 ;
      RECT 36.36 2.55 36.365 3.205 ;
      RECT 35.25 2.365 35.54 2.595 ;
      RECT 35.31 0.885 35.48 2.595 ;
      RECT 35.275 1.095 35.625 1.445 ;
      RECT 35.25 0.885 35.54 1.115 ;
      RECT 35.25 7.765 35.54 7.995 ;
      RECT 35.31 6.285 35.48 7.995 ;
      RECT 35.25 6.285 35.54 6.515 ;
      RECT 34.84 2.735 35.17 2.965 ;
      RECT 34.84 2.765 35.34 2.935 ;
      RECT 34.84 2.395 35.03 2.965 ;
      RECT 34.26 2.365 34.55 2.595 ;
      RECT 34.26 2.395 35.03 2.565 ;
      RECT 34.32 0.885 34.49 2.595 ;
      RECT 34.26 0.885 34.55 1.115 ;
      RECT 34.26 7.765 34.55 7.995 ;
      RECT 34.32 6.285 34.49 7.995 ;
      RECT 34.26 6.285 34.55 6.515 ;
      RECT 34.26 6.325 35.11 6.485 ;
      RECT 34.94 5.915 35.11 6.485 ;
      RECT 34.26 6.32 34.65 6.485 ;
      RECT 34.88 5.915 35.17 6.145 ;
      RECT 34.88 5.945 35.34 6.115 ;
      RECT 33.89 2.735 34.18 2.965 ;
      RECT 33.89 2.765 34.35 2.935 ;
      RECT 33.95 1.655 34.115 2.965 ;
      RECT 32.465 1.625 32.755 1.855 ;
      RECT 32.465 1.655 34.115 1.825 ;
      RECT 32.525 0.885 32.695 1.855 ;
      RECT 32.465 0.885 32.755 1.115 ;
      RECT 32.465 7.765 32.755 7.995 ;
      RECT 32.525 7.025 32.695 7.995 ;
      RECT 32.525 7.12 34.115 7.29 ;
      RECT 33.945 5.915 34.115 7.29 ;
      RECT 32.465 7.025 32.755 7.255 ;
      RECT 33.89 5.915 34.18 6.145 ;
      RECT 33.89 5.945 34.35 6.115 ;
      RECT 32.895 1.965 33.245 2.315 ;
      RECT 32.725 2.025 33.245 2.195 ;
      RECT 32.92 6.655 33.245 6.98 ;
      RECT 32.895 6.655 33.245 6.885 ;
      RECT 32.725 6.685 33.245 6.855 ;
      RECT 30.5 3.43 30.85 3.78 ;
      RECT 30.59 2.395 30.76 3.78 ;
      RECT 32.12 2.365 32.44 2.685 ;
      RECT 32.09 2.365 32.44 2.595 ;
      RECT 30.59 2.395 32.44 2.565 ;
      RECT 32.12 6.28 32.44 6.605 ;
      RECT 32.09 6.285 32.44 6.515 ;
      RECT 31.92 6.315 32.44 6.485 ;
      RECT 31.075 2.705 31.425 3.055 ;
      RECT 31.075 2.765 31.555 2.935 ;
      RECT 31.065 5.84 31.415 6.19 ;
      RECT 31.065 5.945 31.555 6.115 ;
      RECT 27.9 3.665 27.94 3.925 ;
      RECT 27.94 3.645 27.945 3.655 ;
      RECT 29.28 2.735 29.435 3.055 ;
      RECT 29.2 2.735 29.28 3.22 ;
      RECT 29.19 2.735 29.2 3.363 ;
      RECT 29.165 2.735 29.19 3.41 ;
      RECT 29.14 2.735 29.165 3.488 ;
      RECT 29.12 2.735 29.14 3.558 ;
      RECT 29.115 2.735 29.12 3.588 ;
      RECT 29.095 2.885 29.115 3.6 ;
      RECT 29.085 2.885 29.095 3.618 ;
      RECT 29.075 2.887 29.085 3.626 ;
      RECT 29.07 2.892 29.075 3.083 ;
      RECT 29.07 3.092 29.075 3.627 ;
      RECT 29.065 3.137 29.07 3.628 ;
      RECT 29.055 3.202 29.065 3.629 ;
      RECT 29.045 3.297 29.055 3.631 ;
      RECT 29.04 3.35 29.045 3.633 ;
      RECT 29.035 3.37 29.04 3.634 ;
      RECT 28.98 3.395 29.035 3.64 ;
      RECT 28.94 3.43 28.98 3.649 ;
      RECT 28.93 3.447 28.94 3.654 ;
      RECT 28.921 3.453 28.93 3.656 ;
      RECT 28.835 3.491 28.921 3.667 ;
      RECT 28.83 3.53 28.835 3.677 ;
      RECT 28.755 3.537 28.83 3.687 ;
      RECT 28.735 3.547 28.755 3.698 ;
      RECT 28.705 3.554 28.735 3.706 ;
      RECT 28.68 3.561 28.705 3.713 ;
      RECT 28.656 3.567 28.68 3.718 ;
      RECT 28.57 3.58 28.656 3.73 ;
      RECT 28.492 3.587 28.57 3.748 ;
      RECT 28.406 3.582 28.492 3.766 ;
      RECT 28.32 3.577 28.406 3.786 ;
      RECT 28.24 3.571 28.32 3.803 ;
      RECT 28.175 3.567 28.24 3.832 ;
      RECT 28.17 3.281 28.175 3.305 ;
      RECT 28.16 3.557 28.175 3.86 ;
      RECT 28.165 3.275 28.17 3.345 ;
      RECT 28.16 3.269 28.165 3.415 ;
      RECT 28.155 3.263 28.16 3.493 ;
      RECT 28.155 3.54 28.16 3.925 ;
      RECT 28.147 3.26 28.155 3.925 ;
      RECT 28.061 3.258 28.147 3.925 ;
      RECT 27.975 3.256 28.061 3.925 ;
      RECT 27.965 3.257 27.975 3.925 ;
      RECT 27.96 3.262 27.965 3.925 ;
      RECT 27.95 3.275 27.96 3.925 ;
      RECT 27.945 3.297 27.95 3.925 ;
      RECT 27.94 3.657 27.945 3.925 ;
      RECT 28.57 3.125 28.575 3.345 ;
      RECT 29.075 2.16 29.11 2.42 ;
      RECT 29.06 2.16 29.075 2.428 ;
      RECT 29.031 2.16 29.06 2.45 ;
      RECT 28.945 2.16 29.031 2.51 ;
      RECT 28.925 2.16 28.945 2.575 ;
      RECT 28.865 2.16 28.925 2.74 ;
      RECT 28.86 2.16 28.865 2.888 ;
      RECT 28.855 2.16 28.86 2.9 ;
      RECT 28.85 2.16 28.855 2.926 ;
      RECT 28.82 2.346 28.85 3.006 ;
      RECT 28.815 2.394 28.82 3.095 ;
      RECT 28.81 2.408 28.815 3.11 ;
      RECT 28.805 2.427 28.81 3.14 ;
      RECT 28.8 2.442 28.805 3.156 ;
      RECT 28.795 2.457 28.8 3.178 ;
      RECT 28.79 2.477 28.795 3.2 ;
      RECT 28.78 2.497 28.79 3.233 ;
      RECT 28.765 2.539 28.78 3.295 ;
      RECT 28.76 2.57 28.765 3.335 ;
      RECT 28.755 2.582 28.76 3.34 ;
      RECT 28.75 2.594 28.755 3.345 ;
      RECT 28.745 2.607 28.75 3.345 ;
      RECT 28.74 2.625 28.745 3.345 ;
      RECT 28.735 2.645 28.74 3.345 ;
      RECT 28.73 2.657 28.735 3.345 ;
      RECT 28.725 2.67 28.73 3.345 ;
      RECT 28.705 2.705 28.725 3.345 ;
      RECT 28.655 2.807 28.705 3.345 ;
      RECT 28.65 2.892 28.655 3.345 ;
      RECT 28.645 2.9 28.65 3.345 ;
      RECT 28.64 2.917 28.645 3.345 ;
      RECT 28.635 2.932 28.64 3.345 ;
      RECT 28.6 2.997 28.635 3.345 ;
      RECT 28.585 3.062 28.6 3.345 ;
      RECT 28.58 3.092 28.585 3.345 ;
      RECT 28.575 3.117 28.58 3.345 ;
      RECT 28.56 3.127 28.57 3.345 ;
      RECT 28.545 3.14 28.56 3.338 ;
      RECT 28.29 2.73 28.36 2.94 ;
      RECT 28.08 2.707 28.085 2.9 ;
      RECT 25.535 2.635 25.795 2.895 ;
      RECT 28.37 2.917 28.375 2.92 ;
      RECT 28.36 2.735 28.37 2.935 ;
      RECT 28.261 2.728 28.29 2.94 ;
      RECT 28.175 2.72 28.261 2.94 ;
      RECT 28.16 2.714 28.175 2.938 ;
      RECT 28.14 2.713 28.16 2.925 ;
      RECT 28.135 2.712 28.14 2.908 ;
      RECT 28.085 2.709 28.135 2.903 ;
      RECT 28.055 2.706 28.08 2.898 ;
      RECT 28.035 2.704 28.055 2.893 ;
      RECT 28.02 2.702 28.035 2.89 ;
      RECT 27.99 2.7 28.02 2.888 ;
      RECT 27.925 2.696 27.99 2.88 ;
      RECT 27.895 2.691 27.925 2.875 ;
      RECT 27.875 2.689 27.895 2.873 ;
      RECT 27.845 2.686 27.875 2.868 ;
      RECT 27.785 2.682 27.845 2.86 ;
      RECT 27.78 2.679 27.785 2.855 ;
      RECT 27.71 2.677 27.78 2.85 ;
      RECT 27.681 2.673 27.71 2.843 ;
      RECT 27.595 2.668 27.681 2.835 ;
      RECT 27.561 2.663 27.595 2.827 ;
      RECT 27.475 2.655 27.561 2.819 ;
      RECT 27.436 2.648 27.475 2.811 ;
      RECT 27.35 2.643 27.436 2.803 ;
      RECT 27.285 2.637 27.35 2.793 ;
      RECT 27.265 2.632 27.285 2.788 ;
      RECT 27.256 2.629 27.265 2.787 ;
      RECT 27.17 2.625 27.256 2.781 ;
      RECT 27.13 2.621 27.17 2.773 ;
      RECT 27.11 2.617 27.13 2.771 ;
      RECT 27.05 2.617 27.11 2.768 ;
      RECT 27.03 2.62 27.05 2.766 ;
      RECT 27.009 2.62 27.03 2.766 ;
      RECT 26.923 2.622 27.009 2.77 ;
      RECT 26.837 2.624 26.923 2.776 ;
      RECT 26.751 2.626 26.837 2.783 ;
      RECT 26.665 2.629 26.751 2.789 ;
      RECT 26.631 2.63 26.665 2.794 ;
      RECT 26.545 2.633 26.631 2.799 ;
      RECT 26.516 2.64 26.545 2.804 ;
      RECT 26.43 2.64 26.516 2.809 ;
      RECT 26.397 2.64 26.43 2.814 ;
      RECT 26.311 2.642 26.397 2.819 ;
      RECT 26.225 2.644 26.311 2.826 ;
      RECT 26.161 2.646 26.225 2.832 ;
      RECT 26.075 2.648 26.161 2.838 ;
      RECT 26.072 2.65 26.075 2.841 ;
      RECT 25.986 2.651 26.072 2.845 ;
      RECT 25.9 2.654 25.986 2.852 ;
      RECT 25.881 2.656 25.9 2.856 ;
      RECT 25.795 2.658 25.881 2.861 ;
      RECT 25.525 2.67 25.535 2.865 ;
      RECT 27.76 2.25 27.945 2.46 ;
      RECT 27.755 2.251 27.95 2.458 ;
      RECT 27.75 2.256 27.96 2.453 ;
      RECT 27.745 2.232 27.75 2.45 ;
      RECT 27.715 2.229 27.745 2.443 ;
      RECT 27.71 2.225 27.715 2.434 ;
      RECT 27.675 2.256 27.96 2.429 ;
      RECT 27.45 2.165 27.71 2.425 ;
      RECT 27.75 2.234 27.755 2.453 ;
      RECT 27.755 2.235 27.76 2.458 ;
      RECT 27.45 2.247 27.83 2.425 ;
      RECT 27.45 2.245 27.815 2.425 ;
      RECT 27.45 2.24 27.805 2.425 ;
      RECT 27.405 3.155 27.455 3.44 ;
      RECT 27.35 3.125 27.355 3.44 ;
      RECT 27.32 3.105 27.325 3.44 ;
      RECT 27.47 3.155 27.53 3.415 ;
      RECT 27.465 3.155 27.47 3.423 ;
      RECT 27.455 3.155 27.465 3.435 ;
      RECT 27.37 3.145 27.405 3.44 ;
      RECT 27.365 3.132 27.37 3.44 ;
      RECT 27.355 3.127 27.365 3.44 ;
      RECT 27.335 3.117 27.35 3.44 ;
      RECT 27.325 3.11 27.335 3.44 ;
      RECT 27.315 3.102 27.32 3.44 ;
      RECT 27.285 3.092 27.315 3.44 ;
      RECT 27.27 3.08 27.285 3.44 ;
      RECT 27.255 3.07 27.27 3.435 ;
      RECT 27.235 3.06 27.255 3.41 ;
      RECT 27.225 3.052 27.235 3.387 ;
      RECT 27.195 3.035 27.225 3.377 ;
      RECT 27.19 3.012 27.195 3.368 ;
      RECT 27.185 2.999 27.19 3.366 ;
      RECT 27.17 2.975 27.185 3.36 ;
      RECT 27.165 2.951 27.17 3.354 ;
      RECT 27.155 2.94 27.165 3.349 ;
      RECT 27.15 2.93 27.155 3.345 ;
      RECT 27.145 2.922 27.15 3.342 ;
      RECT 27.135 2.917 27.145 3.338 ;
      RECT 27.13 2.912 27.135 3.334 ;
      RECT 27.045 2.91 27.13 3.309 ;
      RECT 27.015 2.91 27.045 3.275 ;
      RECT 27 2.91 27.015 3.258 ;
      RECT 26.945 2.91 27 3.203 ;
      RECT 26.94 2.915 26.945 3.152 ;
      RECT 26.93 2.92 26.94 3.142 ;
      RECT 26.925 2.93 26.93 3.128 ;
      RECT 26.875 3.67 27.135 3.93 ;
      RECT 26.795 3.685 27.135 3.906 ;
      RECT 26.775 3.685 27.135 3.901 ;
      RECT 26.751 3.685 27.135 3.899 ;
      RECT 26.665 3.685 27.135 3.894 ;
      RECT 26.515 3.625 26.775 3.89 ;
      RECT 26.47 3.685 27.135 3.885 ;
      RECT 26.465 3.692 27.135 3.88 ;
      RECT 26.48 3.68 26.795 3.89 ;
      RECT 26.37 2.115 26.63 2.375 ;
      RECT 26.37 2.172 26.635 2.368 ;
      RECT 26.37 2.202 26.64 2.3 ;
      RECT 26.43 2.633 26.545 2.635 ;
      RECT 26.516 2.63 26.545 2.635 ;
      RECT 25.54 3.634 25.565 3.874 ;
      RECT 25.525 3.637 25.615 3.868 ;
      RECT 25.52 3.642 25.701 3.863 ;
      RECT 25.515 3.65 25.765 3.861 ;
      RECT 25.515 3.65 25.775 3.86 ;
      RECT 25.51 3.657 25.785 3.853 ;
      RECT 25.51 3.657 25.871 3.842 ;
      RECT 25.505 3.692 25.871 3.838 ;
      RECT 25.505 3.692 25.88 3.827 ;
      RECT 25.785 3.565 26.045 3.825 ;
      RECT 25.495 3.742 26.045 3.823 ;
      RECT 25.765 3.61 25.785 3.858 ;
      RECT 25.701 3.613 25.765 3.862 ;
      RECT 25.615 3.618 25.701 3.867 ;
      RECT 25.545 3.629 26.045 3.825 ;
      RECT 25.565 3.623 25.615 3.872 ;
      RECT 25.69 2.1 25.7 2.362 ;
      RECT 25.68 2.157 25.69 2.365 ;
      RECT 25.655 2.162 25.68 2.371 ;
      RECT 25.63 2.166 25.655 2.383 ;
      RECT 25.62 2.169 25.63 2.393 ;
      RECT 25.615 2.17 25.62 2.398 ;
      RECT 25.61 2.171 25.615 2.403 ;
      RECT 25.605 2.172 25.61 2.405 ;
      RECT 25.58 2.175 25.605 2.408 ;
      RECT 25.55 2.181 25.58 2.411 ;
      RECT 25.485 2.192 25.55 2.414 ;
      RECT 25.44 2.2 25.485 2.418 ;
      RECT 25.425 2.2 25.44 2.426 ;
      RECT 25.42 2.201 25.425 2.433 ;
      RECT 25.415 2.203 25.42 2.436 ;
      RECT 25.41 2.207 25.415 2.439 ;
      RECT 25.4 2.215 25.41 2.443 ;
      RECT 25.395 2.228 25.4 2.448 ;
      RECT 25.39 2.236 25.395 2.45 ;
      RECT 25.385 2.242 25.39 2.45 ;
      RECT 25.38 2.246 25.385 2.453 ;
      RECT 25.375 2.248 25.38 2.456 ;
      RECT 25.37 2.251 25.375 2.459 ;
      RECT 25.36 2.256 25.37 2.463 ;
      RECT 25.355 2.262 25.36 2.468 ;
      RECT 25.345 2.268 25.355 2.472 ;
      RECT 25.33 2.275 25.345 2.478 ;
      RECT 25.301 2.289 25.33 2.488 ;
      RECT 25.215 2.324 25.301 2.52 ;
      RECT 25.195 2.357 25.215 2.549 ;
      RECT 25.175 2.37 25.195 2.56 ;
      RECT 25.155 2.382 25.175 2.571 ;
      RECT 25.105 2.404 25.155 2.591 ;
      RECT 25.09 2.422 25.105 2.608 ;
      RECT 25.085 2.428 25.09 2.611 ;
      RECT 25.08 2.432 25.085 2.614 ;
      RECT 25.075 2.436 25.08 2.618 ;
      RECT 25.07 2.438 25.075 2.621 ;
      RECT 25.06 2.445 25.07 2.624 ;
      RECT 25.055 2.45 25.06 2.628 ;
      RECT 25.05 2.452 25.055 2.631 ;
      RECT 25.045 2.456 25.05 2.634 ;
      RECT 25.04 2.458 25.045 2.638 ;
      RECT 25.025 2.463 25.04 2.643 ;
      RECT 25.02 2.468 25.025 2.646 ;
      RECT 25.015 2.476 25.02 2.649 ;
      RECT 25.01 2.478 25.015 2.652 ;
      RECT 25.005 2.48 25.01 2.655 ;
      RECT 24.995 2.482 25.005 2.661 ;
      RECT 24.96 2.496 24.995 2.673 ;
      RECT 24.95 2.511 24.96 2.683 ;
      RECT 24.875 2.54 24.95 2.707 ;
      RECT 24.87 2.565 24.875 2.73 ;
      RECT 24.855 2.569 24.87 2.736 ;
      RECT 24.845 2.577 24.855 2.741 ;
      RECT 24.815 2.59 24.845 2.745 ;
      RECT 24.805 2.605 24.815 2.75 ;
      RECT 24.795 2.61 24.805 2.753 ;
      RECT 24.79 2.612 24.795 2.755 ;
      RECT 24.775 2.615 24.79 2.758 ;
      RECT 24.77 2.617 24.775 2.761 ;
      RECT 24.75 2.622 24.77 2.765 ;
      RECT 24.72 2.627 24.75 2.773 ;
      RECT 24.695 2.634 24.72 2.781 ;
      RECT 24.69 2.639 24.695 2.786 ;
      RECT 24.66 2.642 24.69 2.79 ;
      RECT 24.62 2.645 24.66 2.8 ;
      RECT 24.585 2.642 24.62 2.812 ;
      RECT 24.575 2.638 24.585 2.819 ;
      RECT 24.55 2.634 24.575 2.825 ;
      RECT 24.545 2.63 24.55 2.83 ;
      RECT 24.505 2.627 24.545 2.83 ;
      RECT 24.49 2.612 24.505 2.831 ;
      RECT 24.467 2.6 24.49 2.831 ;
      RECT 24.381 2.6 24.467 2.832 ;
      RECT 24.295 2.6 24.381 2.834 ;
      RECT 24.275 2.6 24.295 2.831 ;
      RECT 24.27 2.605 24.275 2.826 ;
      RECT 24.265 2.61 24.27 2.824 ;
      RECT 24.255 2.62 24.265 2.822 ;
      RECT 24.25 2.626 24.255 2.815 ;
      RECT 24.245 2.628 24.25 2.8 ;
      RECT 24.24 2.632 24.245 2.79 ;
      RECT 25.7 2.1 25.95 2.36 ;
      RECT 23.425 3.635 23.685 3.895 ;
      RECT 25.72 3.125 25.725 3.335 ;
      RECT 25.725 3.13 25.735 3.33 ;
      RECT 25.675 3.125 25.72 3.35 ;
      RECT 25.665 3.125 25.675 3.37 ;
      RECT 25.646 3.125 25.665 3.375 ;
      RECT 25.56 3.125 25.646 3.372 ;
      RECT 25.53 3.127 25.56 3.37 ;
      RECT 25.475 3.137 25.53 3.368 ;
      RECT 25.41 3.151 25.475 3.366 ;
      RECT 25.405 3.159 25.41 3.365 ;
      RECT 25.39 3.162 25.405 3.363 ;
      RECT 25.325 3.172 25.39 3.359 ;
      RECT 25.277 3.186 25.325 3.36 ;
      RECT 25.191 3.203 25.277 3.374 ;
      RECT 25.105 3.224 25.191 3.391 ;
      RECT 25.085 3.237 25.105 3.401 ;
      RECT 25.04 3.245 25.085 3.408 ;
      RECT 25.005 3.253 25.04 3.416 ;
      RECT 24.971 3.261 25.005 3.424 ;
      RECT 24.885 3.275 24.971 3.436 ;
      RECT 24.85 3.292 24.885 3.448 ;
      RECT 24.841 3.301 24.85 3.452 ;
      RECT 24.755 3.319 24.841 3.469 ;
      RECT 24.696 3.346 24.755 3.496 ;
      RECT 24.61 3.373 24.696 3.524 ;
      RECT 24.59 3.395 24.61 3.544 ;
      RECT 24.53 3.41 24.59 3.56 ;
      RECT 24.52 3.422 24.53 3.573 ;
      RECT 24.515 3.427 24.52 3.576 ;
      RECT 24.505 3.43 24.515 3.579 ;
      RECT 24.5 3.432 24.505 3.582 ;
      RECT 24.47 3.44 24.5 3.589 ;
      RECT 24.455 3.447 24.47 3.597 ;
      RECT 24.445 3.452 24.455 3.601 ;
      RECT 24.44 3.455 24.445 3.604 ;
      RECT 24.43 3.457 24.44 3.607 ;
      RECT 24.395 3.467 24.43 3.616 ;
      RECT 24.32 3.49 24.395 3.638 ;
      RECT 24.3 3.508 24.32 3.656 ;
      RECT 24.27 3.515 24.3 3.666 ;
      RECT 24.25 3.523 24.27 3.676 ;
      RECT 24.24 3.529 24.25 3.683 ;
      RECT 24.221 3.534 24.24 3.689 ;
      RECT 24.135 3.554 24.221 3.709 ;
      RECT 24.12 3.574 24.135 3.728 ;
      RECT 24.075 3.586 24.12 3.739 ;
      RECT 24.01 3.607 24.075 3.762 ;
      RECT 23.97 3.627 24.01 3.783 ;
      RECT 23.96 3.637 23.97 3.793 ;
      RECT 23.91 3.649 23.96 3.804 ;
      RECT 23.89 3.665 23.91 3.816 ;
      RECT 23.86 3.675 23.89 3.822 ;
      RECT 23.85 3.68 23.86 3.824 ;
      RECT 23.781 3.681 23.85 3.83 ;
      RECT 23.695 3.683 23.781 3.84 ;
      RECT 23.685 3.684 23.695 3.845 ;
      RECT 24.955 3.71 25.145 3.92 ;
      RECT 24.945 3.715 25.155 3.913 ;
      RECT 24.93 3.715 25.155 3.878 ;
      RECT 24.85 3.6 25.11 3.86 ;
      RECT 23.765 3.13 23.95 3.425 ;
      RECT 23.755 3.13 23.95 3.423 ;
      RECT 23.74 3.13 23.955 3.418 ;
      RECT 23.74 3.13 23.96 3.415 ;
      RECT 23.735 3.13 23.96 3.413 ;
      RECT 23.73 3.385 23.96 3.403 ;
      RECT 23.735 3.13 23.995 3.39 ;
      RECT 23.695 2.165 23.955 2.425 ;
      RECT 23.505 2.09 23.591 2.423 ;
      RECT 23.48 2.094 23.635 2.419 ;
      RECT 23.591 2.086 23.635 2.419 ;
      RECT 23.591 2.087 23.64 2.418 ;
      RECT 23.505 2.092 23.655 2.417 ;
      RECT 23.48 2.1 23.695 2.416 ;
      RECT 23.475 2.095 23.655 2.411 ;
      RECT 23.465 2.11 23.695 2.318 ;
      RECT 23.465 2.162 23.895 2.318 ;
      RECT 23.465 2.155 23.875 2.318 ;
      RECT 23.465 2.142 23.845 2.318 ;
      RECT 23.465 2.13 23.785 2.318 ;
      RECT 23.465 2.115 23.76 2.318 ;
      RECT 22.665 2.745 22.8 3.04 ;
      RECT 22.925 2.768 22.93 2.955 ;
      RECT 23.645 2.665 23.79 2.9 ;
      RECT 23.805 2.665 23.81 2.89 ;
      RECT 23.84 2.676 23.845 2.87 ;
      RECT 23.835 2.668 23.84 2.875 ;
      RECT 23.815 2.665 23.835 2.88 ;
      RECT 23.81 2.665 23.815 2.888 ;
      RECT 23.8 2.665 23.805 2.893 ;
      RECT 23.79 2.665 23.8 2.898 ;
      RECT 23.62 2.667 23.645 2.9 ;
      RECT 23.57 2.674 23.62 2.9 ;
      RECT 23.565 2.679 23.57 2.9 ;
      RECT 23.526 2.684 23.565 2.901 ;
      RECT 23.44 2.696 23.526 2.902 ;
      RECT 23.431 2.706 23.44 2.902 ;
      RECT 23.345 2.715 23.431 2.904 ;
      RECT 23.321 2.725 23.345 2.906 ;
      RECT 23.235 2.736 23.321 2.907 ;
      RECT 23.205 2.747 23.235 2.909 ;
      RECT 23.175 2.752 23.205 2.911 ;
      RECT 23.15 2.758 23.175 2.914 ;
      RECT 23.135 2.763 23.15 2.915 ;
      RECT 23.09 2.769 23.135 2.915 ;
      RECT 23.085 2.774 23.09 2.916 ;
      RECT 23.065 2.774 23.085 2.918 ;
      RECT 23.045 2.772 23.065 2.923 ;
      RECT 23.01 2.771 23.045 2.93 ;
      RECT 22.98 2.77 23.01 2.94 ;
      RECT 22.93 2.769 22.98 2.95 ;
      RECT 22.84 2.766 22.925 3.04 ;
      RECT 22.815 2.76 22.84 3.04 ;
      RECT 22.8 2.75 22.815 3.04 ;
      RECT 22.615 2.745 22.665 2.96 ;
      RECT 22.605 2.75 22.615 2.95 ;
      RECT 22.845 3.225 23.105 3.485 ;
      RECT 22.845 3.225 23.135 3.378 ;
      RECT 22.845 3.225 23.17 3.363 ;
      RECT 23.1 3.145 23.29 3.355 ;
      RECT 23.09 3.15 23.3 3.348 ;
      RECT 23.055 3.22 23.3 3.348 ;
      RECT 23.085 3.162 23.105 3.485 ;
      RECT 23.07 3.21 23.3 3.348 ;
      RECT 23.075 3.182 23.105 3.485 ;
      RECT 22.155 2.25 22.225 3.355 ;
      RECT 22.89 2.355 23.15 2.615 ;
      RECT 22.47 2.401 22.485 2.61 ;
      RECT 22.806 2.414 22.89 2.565 ;
      RECT 22.72 2.411 22.806 2.565 ;
      RECT 22.681 2.409 22.72 2.565 ;
      RECT 22.595 2.407 22.681 2.565 ;
      RECT 22.535 2.405 22.595 2.576 ;
      RECT 22.5 2.403 22.535 2.594 ;
      RECT 22.485 2.401 22.5 2.605 ;
      RECT 22.455 2.401 22.47 2.618 ;
      RECT 22.445 2.401 22.455 2.623 ;
      RECT 22.42 2.4 22.445 2.628 ;
      RECT 22.405 2.395 22.42 2.634 ;
      RECT 22.4 2.388 22.405 2.639 ;
      RECT 22.375 2.379 22.4 2.645 ;
      RECT 22.33 2.358 22.375 2.658 ;
      RECT 22.32 2.342 22.33 2.668 ;
      RECT 22.305 2.335 22.32 2.678 ;
      RECT 22.295 2.328 22.305 2.695 ;
      RECT 22.29 2.325 22.295 2.725 ;
      RECT 22.285 2.323 22.29 2.755 ;
      RECT 22.28 2.321 22.285 2.792 ;
      RECT 22.265 2.317 22.28 2.859 ;
      RECT 22.265 3.15 22.275 3.35 ;
      RECT 22.26 2.313 22.265 2.985 ;
      RECT 22.26 3.137 22.265 3.355 ;
      RECT 22.255 2.311 22.26 3.07 ;
      RECT 22.255 3.127 22.26 3.355 ;
      RECT 22.24 2.282 22.255 3.355 ;
      RECT 22.225 2.255 22.24 3.355 ;
      RECT 22.15 2.25 22.155 2.605 ;
      RECT 22.15 2.66 22.155 3.355 ;
      RECT 22.135 2.25 22.15 2.583 ;
      RECT 22.145 2.682 22.15 3.355 ;
      RECT 22.135 2.722 22.145 3.355 ;
      RECT 22.1 2.25 22.135 2.525 ;
      RECT 22.13 2.757 22.135 3.355 ;
      RECT 22.115 2.812 22.13 3.355 ;
      RECT 22.11 2.877 22.115 3.355 ;
      RECT 22.095 2.925 22.11 3.355 ;
      RECT 22.07 2.25 22.1 2.48 ;
      RECT 22.09 2.98 22.095 3.355 ;
      RECT 22.075 3.04 22.09 3.355 ;
      RECT 22.07 3.088 22.075 3.353 ;
      RECT 22.065 2.25 22.07 2.473 ;
      RECT 22.065 3.12 22.07 3.348 ;
      RECT 22.04 2.25 22.065 2.465 ;
      RECT 22.03 2.255 22.04 2.455 ;
      RECT 22.245 3.53 22.265 3.77 ;
      RECT 21.475 3.46 21.48 3.67 ;
      RECT 22.755 3.533 22.765 3.728 ;
      RECT 22.75 3.523 22.755 3.731 ;
      RECT 22.67 3.52 22.75 3.754 ;
      RECT 22.666 3.52 22.67 3.776 ;
      RECT 22.58 3.52 22.666 3.786 ;
      RECT 22.565 3.52 22.58 3.794 ;
      RECT 22.536 3.521 22.565 3.792 ;
      RECT 22.45 3.526 22.536 3.788 ;
      RECT 22.437 3.53 22.45 3.784 ;
      RECT 22.351 3.53 22.437 3.78 ;
      RECT 22.265 3.53 22.351 3.774 ;
      RECT 22.181 3.53 22.245 3.768 ;
      RECT 22.095 3.53 22.181 3.763 ;
      RECT 22.075 3.53 22.095 3.759 ;
      RECT 22.015 3.525 22.075 3.756 ;
      RECT 21.987 3.519 22.015 3.753 ;
      RECT 21.901 3.514 21.987 3.749 ;
      RECT 21.815 3.508 21.901 3.743 ;
      RECT 21.74 3.49 21.815 3.738 ;
      RECT 21.705 3.467 21.74 3.734 ;
      RECT 21.695 3.457 21.705 3.733 ;
      RECT 21.64 3.455 21.695 3.732 ;
      RECT 21.565 3.455 21.64 3.728 ;
      RECT 21.555 3.455 21.565 3.723 ;
      RECT 21.54 3.455 21.555 3.715 ;
      RECT 21.49 3.457 21.54 3.693 ;
      RECT 21.48 3.46 21.49 3.673 ;
      RECT 21.47 3.465 21.475 3.668 ;
      RECT 21.465 3.47 21.47 3.663 ;
      RECT 21.59 2.635 21.85 2.895 ;
      RECT 21.59 2.65 21.87 2.86 ;
      RECT 21.59 2.655 21.88 2.855 ;
      RECT 19.575 2.115 19.835 2.375 ;
      RECT 19.565 2.145 19.835 2.355 ;
      RECT 21.485 2.06 21.745 2.32 ;
      RECT 21.48 2.135 21.485 2.321 ;
      RECT 21.455 2.14 21.48 2.323 ;
      RECT 21.44 2.147 21.455 2.326 ;
      RECT 21.38 2.165 21.44 2.331 ;
      RECT 21.35 2.185 21.38 2.338 ;
      RECT 21.325 2.193 21.35 2.343 ;
      RECT 21.3 2.201 21.325 2.345 ;
      RECT 21.282 2.205 21.3 2.344 ;
      RECT 21.196 2.203 21.282 2.344 ;
      RECT 21.11 2.201 21.196 2.344 ;
      RECT 21.024 2.199 21.11 2.343 ;
      RECT 20.938 2.197 21.024 2.343 ;
      RECT 20.852 2.195 20.938 2.343 ;
      RECT 20.766 2.193 20.852 2.343 ;
      RECT 20.68 2.191 20.766 2.342 ;
      RECT 20.662 2.19 20.68 2.342 ;
      RECT 20.576 2.189 20.662 2.342 ;
      RECT 20.49 2.187 20.576 2.342 ;
      RECT 20.404 2.186 20.49 2.341 ;
      RECT 20.318 2.185 20.404 2.341 ;
      RECT 20.232 2.183 20.318 2.341 ;
      RECT 20.146 2.182 20.232 2.341 ;
      RECT 20.06 2.18 20.146 2.34 ;
      RECT 20.036 2.178 20.06 2.34 ;
      RECT 19.95 2.171 20.036 2.34 ;
      RECT 19.921 2.163 19.95 2.34 ;
      RECT 19.835 2.155 19.921 2.34 ;
      RECT 19.555 2.152 19.565 2.35 ;
      RECT 21.06 3.115 21.065 3.465 ;
      RECT 20.83 3.205 20.97 3.465 ;
      RECT 21.305 2.89 21.35 3.1 ;
      RECT 21.36 2.901 21.37 3.095 ;
      RECT 21.35 2.893 21.36 3.1 ;
      RECT 21.285 2.89 21.305 3.105 ;
      RECT 21.255 2.89 21.285 3.128 ;
      RECT 21.245 2.89 21.255 3.153 ;
      RECT 21.24 2.89 21.245 3.163 ;
      RECT 21.185 2.89 21.24 3.203 ;
      RECT 21.18 2.89 21.185 3.243 ;
      RECT 21.175 2.892 21.18 3.248 ;
      RECT 21.16 2.902 21.175 3.259 ;
      RECT 21.115 2.96 21.16 3.295 ;
      RECT 21.105 3.015 21.115 3.329 ;
      RECT 21.09 3.042 21.105 3.345 ;
      RECT 21.08 3.069 21.09 3.465 ;
      RECT 21.065 3.092 21.08 3.465 ;
      RECT 21.055 3.132 21.06 3.465 ;
      RECT 21.05 3.142 21.055 3.465 ;
      RECT 21.045 3.157 21.05 3.465 ;
      RECT 21.035 3.162 21.045 3.465 ;
      RECT 20.97 3.185 21.035 3.465 ;
      RECT 20.47 2.68 20.66 2.89 ;
      RECT 19.045 2.605 19.305 2.865 ;
      RECT 19.395 2.6 19.49 2.81 ;
      RECT 19.37 2.615 19.38 2.81 ;
      RECT 20.66 2.687 20.67 2.885 ;
      RECT 20.46 2.687 20.47 2.885 ;
      RECT 20.445 2.702 20.46 2.875 ;
      RECT 20.44 2.71 20.445 2.868 ;
      RECT 20.43 2.713 20.44 2.865 ;
      RECT 20.395 2.712 20.43 2.863 ;
      RECT 20.366 2.708 20.395 2.86 ;
      RECT 20.28 2.703 20.366 2.857 ;
      RECT 20.22 2.697 20.28 2.853 ;
      RECT 20.191 2.693 20.22 2.85 ;
      RECT 20.105 2.685 20.191 2.847 ;
      RECT 20.096 2.679 20.105 2.845 ;
      RECT 20.01 2.674 20.096 2.843 ;
      RECT 19.987 2.669 20.01 2.84 ;
      RECT 19.901 2.663 19.987 2.837 ;
      RECT 19.815 2.654 19.901 2.832 ;
      RECT 19.805 2.649 19.815 2.83 ;
      RECT 19.786 2.648 19.805 2.829 ;
      RECT 19.7 2.643 19.786 2.825 ;
      RECT 19.68 2.638 19.7 2.821 ;
      RECT 19.62 2.633 19.68 2.818 ;
      RECT 19.595 2.623 19.62 2.816 ;
      RECT 19.59 2.616 19.595 2.815 ;
      RECT 19.58 2.607 19.59 2.814 ;
      RECT 19.576 2.6 19.58 2.814 ;
      RECT 19.49 2.6 19.576 2.812 ;
      RECT 19.38 2.607 19.395 2.81 ;
      RECT 19.365 2.617 19.37 2.81 ;
      RECT 19.345 2.62 19.365 2.807 ;
      RECT 19.315 2.62 19.345 2.803 ;
      RECT 19.305 2.62 19.315 2.803 ;
      RECT 20.22 3.115 20.48 3.375 ;
      RECT 20.15 3.125 20.48 3.335 ;
      RECT 20.14 3.132 20.48 3.33 ;
      RECT 19.56 3.12 19.82 3.38 ;
      RECT 19.56 3.16 19.925 3.37 ;
      RECT 19.56 3.162 19.93 3.369 ;
      RECT 19.56 3.17 19.935 3.366 ;
      RECT 18.485 2.245 18.585 3.77 ;
      RECT 18.675 3.385 18.725 3.645 ;
      RECT 18.67 2.258 18.675 2.445 ;
      RECT 18.665 3.366 18.675 3.645 ;
      RECT 18.665 2.255 18.67 2.453 ;
      RECT 18.65 2.249 18.665 2.46 ;
      RECT 18.66 3.354 18.665 3.728 ;
      RECT 18.65 3.342 18.66 3.765 ;
      RECT 18.64 2.245 18.65 2.467 ;
      RECT 18.64 3.327 18.65 3.77 ;
      RECT 18.635 2.245 18.64 2.475 ;
      RECT 18.615 3.297 18.64 3.77 ;
      RECT 18.595 2.245 18.635 2.523 ;
      RECT 18.605 3.257 18.615 3.77 ;
      RECT 18.595 3.212 18.605 3.77 ;
      RECT 18.59 2.245 18.595 2.593 ;
      RECT 18.59 3.17 18.595 3.77 ;
      RECT 18.585 2.245 18.59 3.07 ;
      RECT 18.585 3.152 18.59 3.77 ;
      RECT 18.475 2.248 18.485 3.77 ;
      RECT 18.46 2.255 18.475 3.766 ;
      RECT 18.455 2.265 18.46 3.761 ;
      RECT 18.45 2.465 18.455 3.653 ;
      RECT 18.445 2.55 18.45 3.205 ;
      RECT 17.33 2.365 17.62 2.595 ;
      RECT 17.39 0.885 17.56 2.595 ;
      RECT 17.305 1.095 17.655 1.445 ;
      RECT 17.33 0.885 17.62 1.445 ;
      RECT 17.33 7.765 17.62 7.995 ;
      RECT 17.39 6.285 17.56 7.995 ;
      RECT 17.33 6.285 17.62 6.515 ;
      RECT 16.92 2.735 17.25 2.965 ;
      RECT 16.92 2.765 17.42 2.935 ;
      RECT 16.92 2.395 17.11 2.965 ;
      RECT 16.34 2.365 16.63 2.595 ;
      RECT 16.34 2.395 17.11 2.565 ;
      RECT 16.4 0.885 16.57 2.595 ;
      RECT 16.34 0.885 16.63 1.115 ;
      RECT 16.34 7.765 16.63 7.995 ;
      RECT 16.4 6.285 16.57 7.995 ;
      RECT 16.34 6.285 16.63 6.515 ;
      RECT 16.34 6.325 17.19 6.485 ;
      RECT 17.02 5.915 17.19 6.485 ;
      RECT 16.34 6.32 16.73 6.485 ;
      RECT 16.96 5.915 17.25 6.145 ;
      RECT 16.96 5.945 17.42 6.115 ;
      RECT 15.97 2.735 16.26 2.965 ;
      RECT 15.97 2.765 16.43 2.935 ;
      RECT 16.03 1.655 16.195 2.965 ;
      RECT 14.545 1.625 14.835 1.855 ;
      RECT 14.545 1.655 16.195 1.825 ;
      RECT 14.605 0.885 14.775 1.855 ;
      RECT 14.545 0.885 14.835 1.115 ;
      RECT 14.545 7.765 14.835 7.995 ;
      RECT 14.605 7.025 14.775 7.995 ;
      RECT 14.605 7.12 16.195 7.29 ;
      RECT 16.025 5.915 16.195 7.29 ;
      RECT 14.545 7.025 14.835 7.255 ;
      RECT 15.97 5.915 16.26 6.145 ;
      RECT 15.97 5.945 16.43 6.115 ;
      RECT 14.975 1.965 15.325 2.315 ;
      RECT 14.805 2.025 15.325 2.195 ;
      RECT 15 6.655 15.325 6.98 ;
      RECT 14.975 6.655 15.325 6.885 ;
      RECT 14.805 6.685 15.325 6.855 ;
      RECT 12.58 3.43 12.93 3.78 ;
      RECT 12.67 2.395 12.84 3.78 ;
      RECT 14.2 2.365 14.52 2.685 ;
      RECT 14.17 2.365 14.52 2.595 ;
      RECT 12.67 2.395 14.52 2.565 ;
      RECT 14.2 6.28 14.52 6.605 ;
      RECT 14.17 6.285 14.52 6.515 ;
      RECT 14 6.315 14.52 6.485 ;
      RECT 13.155 2.705 13.505 3.055 ;
      RECT 13.155 2.765 13.635 2.935 ;
      RECT 13.145 5.84 13.495 6.19 ;
      RECT 13.145 5.945 13.635 6.115 ;
      RECT 9.98 3.665 10.02 3.925 ;
      RECT 10.02 3.645 10.025 3.655 ;
      RECT 11.36 2.735 11.515 3.055 ;
      RECT 11.28 2.735 11.36 3.22 ;
      RECT 11.27 2.735 11.28 3.363 ;
      RECT 11.245 2.735 11.27 3.41 ;
      RECT 11.22 2.735 11.245 3.488 ;
      RECT 11.2 2.735 11.22 3.558 ;
      RECT 11.195 2.735 11.2 3.588 ;
      RECT 11.175 2.885 11.195 3.6 ;
      RECT 11.165 2.885 11.175 3.618 ;
      RECT 11.155 2.887 11.165 3.626 ;
      RECT 11.15 2.892 11.155 3.083 ;
      RECT 11.15 3.092 11.155 3.627 ;
      RECT 11.145 3.137 11.15 3.628 ;
      RECT 11.135 3.202 11.145 3.629 ;
      RECT 11.125 3.297 11.135 3.631 ;
      RECT 11.12 3.35 11.125 3.633 ;
      RECT 11.115 3.37 11.12 3.634 ;
      RECT 11.06 3.395 11.115 3.64 ;
      RECT 11.02 3.43 11.06 3.649 ;
      RECT 11.01 3.447 11.02 3.654 ;
      RECT 11.001 3.453 11.01 3.656 ;
      RECT 10.915 3.491 11.001 3.667 ;
      RECT 10.91 3.53 10.915 3.677 ;
      RECT 10.835 3.537 10.91 3.687 ;
      RECT 10.815 3.547 10.835 3.698 ;
      RECT 10.785 3.554 10.815 3.706 ;
      RECT 10.76 3.561 10.785 3.713 ;
      RECT 10.736 3.567 10.76 3.718 ;
      RECT 10.65 3.58 10.736 3.73 ;
      RECT 10.572 3.587 10.65 3.748 ;
      RECT 10.486 3.582 10.572 3.766 ;
      RECT 10.4 3.577 10.486 3.786 ;
      RECT 10.32 3.571 10.4 3.803 ;
      RECT 10.255 3.567 10.32 3.832 ;
      RECT 10.25 3.281 10.255 3.305 ;
      RECT 10.24 3.557 10.255 3.86 ;
      RECT 10.245 3.275 10.25 3.345 ;
      RECT 10.24 3.269 10.245 3.415 ;
      RECT 10.235 3.263 10.24 3.493 ;
      RECT 10.235 3.54 10.24 3.925 ;
      RECT 10.227 3.26 10.235 3.925 ;
      RECT 10.141 3.258 10.227 3.925 ;
      RECT 10.055 3.256 10.141 3.925 ;
      RECT 10.045 3.257 10.055 3.925 ;
      RECT 10.04 3.262 10.045 3.925 ;
      RECT 10.03 3.275 10.04 3.925 ;
      RECT 10.025 3.297 10.03 3.925 ;
      RECT 10.02 3.657 10.025 3.925 ;
      RECT 10.65 3.125 10.655 3.345 ;
      RECT 11.155 2.16 11.19 2.42 ;
      RECT 11.14 2.16 11.155 2.428 ;
      RECT 11.111 2.16 11.14 2.45 ;
      RECT 11.025 2.16 11.111 2.51 ;
      RECT 11.005 2.16 11.025 2.575 ;
      RECT 10.945 2.16 11.005 2.74 ;
      RECT 10.94 2.16 10.945 2.888 ;
      RECT 10.935 2.16 10.94 2.9 ;
      RECT 10.93 2.16 10.935 2.926 ;
      RECT 10.9 2.346 10.93 3.006 ;
      RECT 10.895 2.394 10.9 3.095 ;
      RECT 10.89 2.408 10.895 3.11 ;
      RECT 10.885 2.427 10.89 3.14 ;
      RECT 10.88 2.442 10.885 3.156 ;
      RECT 10.875 2.457 10.88 3.178 ;
      RECT 10.87 2.477 10.875 3.2 ;
      RECT 10.86 2.497 10.87 3.233 ;
      RECT 10.845 2.539 10.86 3.295 ;
      RECT 10.84 2.57 10.845 3.335 ;
      RECT 10.835 2.582 10.84 3.34 ;
      RECT 10.83 2.594 10.835 3.345 ;
      RECT 10.825 2.607 10.83 3.345 ;
      RECT 10.82 2.625 10.825 3.345 ;
      RECT 10.815 2.645 10.82 3.345 ;
      RECT 10.81 2.657 10.815 3.345 ;
      RECT 10.805 2.67 10.81 3.345 ;
      RECT 10.785 2.705 10.805 3.345 ;
      RECT 10.735 2.807 10.785 3.345 ;
      RECT 10.73 2.892 10.735 3.345 ;
      RECT 10.725 2.9 10.73 3.345 ;
      RECT 10.72 2.917 10.725 3.345 ;
      RECT 10.715 2.932 10.72 3.345 ;
      RECT 10.68 2.997 10.715 3.345 ;
      RECT 10.665 3.062 10.68 3.345 ;
      RECT 10.66 3.092 10.665 3.345 ;
      RECT 10.655 3.117 10.66 3.345 ;
      RECT 10.64 3.127 10.65 3.345 ;
      RECT 10.625 3.14 10.64 3.338 ;
      RECT 10.37 2.73 10.44 2.94 ;
      RECT 10.16 2.707 10.165 2.9 ;
      RECT 7.615 2.635 7.875 2.895 ;
      RECT 10.45 2.917 10.455 2.92 ;
      RECT 10.44 2.735 10.45 2.935 ;
      RECT 10.341 2.728 10.37 2.94 ;
      RECT 10.255 2.72 10.341 2.94 ;
      RECT 10.24 2.714 10.255 2.938 ;
      RECT 10.22 2.713 10.24 2.925 ;
      RECT 10.215 2.712 10.22 2.908 ;
      RECT 10.165 2.709 10.215 2.903 ;
      RECT 10.135 2.706 10.16 2.898 ;
      RECT 10.115 2.704 10.135 2.893 ;
      RECT 10.1 2.702 10.115 2.89 ;
      RECT 10.07 2.7 10.1 2.888 ;
      RECT 10.005 2.696 10.07 2.88 ;
      RECT 9.975 2.691 10.005 2.875 ;
      RECT 9.955 2.689 9.975 2.873 ;
      RECT 9.925 2.686 9.955 2.868 ;
      RECT 9.865 2.682 9.925 2.86 ;
      RECT 9.86 2.679 9.865 2.855 ;
      RECT 9.79 2.677 9.86 2.85 ;
      RECT 9.761 2.673 9.79 2.843 ;
      RECT 9.675 2.668 9.761 2.835 ;
      RECT 9.641 2.663 9.675 2.827 ;
      RECT 9.555 2.655 9.641 2.819 ;
      RECT 9.516 2.648 9.555 2.811 ;
      RECT 9.43 2.643 9.516 2.803 ;
      RECT 9.365 2.637 9.43 2.793 ;
      RECT 9.345 2.632 9.365 2.788 ;
      RECT 9.336 2.629 9.345 2.787 ;
      RECT 9.25 2.625 9.336 2.781 ;
      RECT 9.21 2.621 9.25 2.773 ;
      RECT 9.19 2.617 9.21 2.771 ;
      RECT 9.13 2.617 9.19 2.768 ;
      RECT 9.11 2.62 9.13 2.766 ;
      RECT 9.089 2.62 9.11 2.766 ;
      RECT 9.003 2.622 9.089 2.77 ;
      RECT 8.917 2.624 9.003 2.776 ;
      RECT 8.831 2.626 8.917 2.783 ;
      RECT 8.745 2.629 8.831 2.789 ;
      RECT 8.711 2.63 8.745 2.794 ;
      RECT 8.625 2.633 8.711 2.799 ;
      RECT 8.596 2.64 8.625 2.804 ;
      RECT 8.51 2.64 8.596 2.809 ;
      RECT 8.477 2.64 8.51 2.814 ;
      RECT 8.391 2.642 8.477 2.819 ;
      RECT 8.305 2.644 8.391 2.826 ;
      RECT 8.241 2.646 8.305 2.832 ;
      RECT 8.155 2.648 8.241 2.838 ;
      RECT 8.152 2.65 8.155 2.841 ;
      RECT 8.066 2.651 8.152 2.845 ;
      RECT 7.98 2.654 8.066 2.852 ;
      RECT 7.961 2.656 7.98 2.856 ;
      RECT 7.875 2.658 7.961 2.861 ;
      RECT 7.605 2.67 7.615 2.865 ;
      RECT 9.84 2.25 10.025 2.46 ;
      RECT 9.835 2.251 10.03 2.458 ;
      RECT 9.83 2.256 10.04 2.453 ;
      RECT 9.825 2.232 9.83 2.45 ;
      RECT 9.795 2.229 9.825 2.443 ;
      RECT 9.79 2.225 9.795 2.434 ;
      RECT 9.755 2.256 10.04 2.429 ;
      RECT 9.53 2.165 9.79 2.425 ;
      RECT 9.83 2.234 9.835 2.453 ;
      RECT 9.835 2.235 9.84 2.458 ;
      RECT 9.53 2.247 9.91 2.425 ;
      RECT 9.53 2.245 9.895 2.425 ;
      RECT 9.53 2.24 9.885 2.425 ;
      RECT 9.485 3.155 9.535 3.44 ;
      RECT 9.43 3.125 9.435 3.44 ;
      RECT 9.4 3.105 9.405 3.44 ;
      RECT 9.55 3.155 9.61 3.415 ;
      RECT 9.545 3.155 9.55 3.423 ;
      RECT 9.535 3.155 9.545 3.435 ;
      RECT 9.45 3.145 9.485 3.44 ;
      RECT 9.445 3.132 9.45 3.44 ;
      RECT 9.435 3.127 9.445 3.44 ;
      RECT 9.415 3.117 9.43 3.44 ;
      RECT 9.405 3.11 9.415 3.44 ;
      RECT 9.395 3.102 9.4 3.44 ;
      RECT 9.365 3.092 9.395 3.44 ;
      RECT 9.35 3.08 9.365 3.44 ;
      RECT 9.335 3.07 9.35 3.435 ;
      RECT 9.315 3.06 9.335 3.41 ;
      RECT 9.305 3.052 9.315 3.387 ;
      RECT 9.275 3.035 9.305 3.377 ;
      RECT 9.27 3.012 9.275 3.368 ;
      RECT 9.265 2.999 9.27 3.366 ;
      RECT 9.25 2.975 9.265 3.36 ;
      RECT 9.245 2.951 9.25 3.354 ;
      RECT 9.235 2.94 9.245 3.349 ;
      RECT 9.23 2.93 9.235 3.345 ;
      RECT 9.225 2.922 9.23 3.342 ;
      RECT 9.215 2.917 9.225 3.338 ;
      RECT 9.21 2.912 9.215 3.334 ;
      RECT 9.125 2.91 9.21 3.309 ;
      RECT 9.095 2.91 9.125 3.275 ;
      RECT 9.08 2.91 9.095 3.258 ;
      RECT 9.025 2.91 9.08 3.203 ;
      RECT 9.02 2.915 9.025 3.152 ;
      RECT 9.01 2.92 9.02 3.142 ;
      RECT 9.005 2.93 9.01 3.128 ;
      RECT 8.955 3.67 9.215 3.93 ;
      RECT 8.875 3.685 9.215 3.906 ;
      RECT 8.855 3.685 9.215 3.901 ;
      RECT 8.831 3.685 9.215 3.899 ;
      RECT 8.745 3.685 9.215 3.894 ;
      RECT 8.595 3.625 8.855 3.89 ;
      RECT 8.55 3.685 9.215 3.885 ;
      RECT 8.545 3.692 9.215 3.88 ;
      RECT 8.56 3.68 8.875 3.89 ;
      RECT 8.45 2.115 8.71 2.375 ;
      RECT 8.45 2.172 8.715 2.368 ;
      RECT 8.45 2.202 8.72 2.3 ;
      RECT 8.51 2.633 8.625 2.635 ;
      RECT 8.596 2.63 8.625 2.635 ;
      RECT 7.62 3.634 7.645 3.874 ;
      RECT 7.605 3.637 7.695 3.868 ;
      RECT 7.6 3.642 7.781 3.863 ;
      RECT 7.595 3.65 7.845 3.861 ;
      RECT 7.595 3.65 7.855 3.86 ;
      RECT 7.59 3.657 7.865 3.853 ;
      RECT 7.59 3.657 7.951 3.842 ;
      RECT 7.585 3.692 7.951 3.838 ;
      RECT 7.585 3.692 7.96 3.827 ;
      RECT 7.865 3.565 8.125 3.825 ;
      RECT 7.575 3.742 8.125 3.823 ;
      RECT 7.845 3.61 7.865 3.858 ;
      RECT 7.781 3.613 7.845 3.862 ;
      RECT 7.695 3.618 7.781 3.867 ;
      RECT 7.625 3.629 8.125 3.825 ;
      RECT 7.645 3.623 7.695 3.872 ;
      RECT 7.77 2.1 7.78 2.362 ;
      RECT 7.76 2.157 7.77 2.365 ;
      RECT 7.735 2.162 7.76 2.371 ;
      RECT 7.71 2.166 7.735 2.383 ;
      RECT 7.7 2.169 7.71 2.393 ;
      RECT 7.695 2.17 7.7 2.398 ;
      RECT 7.69 2.171 7.695 2.403 ;
      RECT 7.685 2.172 7.69 2.405 ;
      RECT 7.66 2.175 7.685 2.408 ;
      RECT 7.63 2.181 7.66 2.411 ;
      RECT 7.565 2.192 7.63 2.414 ;
      RECT 7.52 2.2 7.565 2.418 ;
      RECT 7.505 2.2 7.52 2.426 ;
      RECT 7.5 2.201 7.505 2.433 ;
      RECT 7.495 2.203 7.5 2.436 ;
      RECT 7.49 2.207 7.495 2.439 ;
      RECT 7.48 2.215 7.49 2.443 ;
      RECT 7.475 2.228 7.48 2.448 ;
      RECT 7.47 2.236 7.475 2.45 ;
      RECT 7.465 2.242 7.47 2.45 ;
      RECT 7.46 2.246 7.465 2.453 ;
      RECT 7.455 2.248 7.46 2.456 ;
      RECT 7.45 2.251 7.455 2.459 ;
      RECT 7.44 2.256 7.45 2.463 ;
      RECT 7.435 2.262 7.44 2.468 ;
      RECT 7.425 2.268 7.435 2.472 ;
      RECT 7.41 2.275 7.425 2.478 ;
      RECT 7.381 2.289 7.41 2.488 ;
      RECT 7.295 2.324 7.381 2.52 ;
      RECT 7.275 2.357 7.295 2.549 ;
      RECT 7.255 2.37 7.275 2.56 ;
      RECT 7.235 2.382 7.255 2.571 ;
      RECT 7.185 2.404 7.235 2.591 ;
      RECT 7.17 2.422 7.185 2.608 ;
      RECT 7.165 2.428 7.17 2.611 ;
      RECT 7.16 2.432 7.165 2.614 ;
      RECT 7.155 2.436 7.16 2.618 ;
      RECT 7.15 2.438 7.155 2.621 ;
      RECT 7.14 2.445 7.15 2.624 ;
      RECT 7.135 2.45 7.14 2.628 ;
      RECT 7.13 2.452 7.135 2.631 ;
      RECT 7.125 2.456 7.13 2.634 ;
      RECT 7.12 2.458 7.125 2.638 ;
      RECT 7.105 2.463 7.12 2.643 ;
      RECT 7.1 2.468 7.105 2.646 ;
      RECT 7.095 2.476 7.1 2.649 ;
      RECT 7.09 2.478 7.095 2.652 ;
      RECT 7.085 2.48 7.09 2.655 ;
      RECT 7.075 2.482 7.085 2.661 ;
      RECT 7.04 2.496 7.075 2.673 ;
      RECT 7.03 2.511 7.04 2.683 ;
      RECT 6.955 2.54 7.03 2.707 ;
      RECT 6.95 2.565 6.955 2.73 ;
      RECT 6.935 2.569 6.95 2.736 ;
      RECT 6.925 2.577 6.935 2.741 ;
      RECT 6.895 2.59 6.925 2.745 ;
      RECT 6.885 2.605 6.895 2.75 ;
      RECT 6.875 2.61 6.885 2.753 ;
      RECT 6.87 2.612 6.875 2.755 ;
      RECT 6.855 2.615 6.87 2.758 ;
      RECT 6.85 2.617 6.855 2.761 ;
      RECT 6.83 2.622 6.85 2.765 ;
      RECT 6.8 2.627 6.83 2.773 ;
      RECT 6.775 2.634 6.8 2.781 ;
      RECT 6.77 2.639 6.775 2.786 ;
      RECT 6.74 2.642 6.77 2.79 ;
      RECT 6.7 2.645 6.74 2.8 ;
      RECT 6.665 2.642 6.7 2.812 ;
      RECT 6.655 2.638 6.665 2.819 ;
      RECT 6.63 2.634 6.655 2.825 ;
      RECT 6.625 2.63 6.63 2.83 ;
      RECT 6.585 2.627 6.625 2.83 ;
      RECT 6.57 2.612 6.585 2.831 ;
      RECT 6.547 2.6 6.57 2.831 ;
      RECT 6.461 2.6 6.547 2.832 ;
      RECT 6.375 2.6 6.461 2.834 ;
      RECT 6.355 2.6 6.375 2.831 ;
      RECT 6.35 2.605 6.355 2.826 ;
      RECT 6.345 2.61 6.35 2.824 ;
      RECT 6.335 2.62 6.345 2.822 ;
      RECT 6.33 2.626 6.335 2.815 ;
      RECT 6.325 2.628 6.33 2.8 ;
      RECT 6.32 2.632 6.325 2.79 ;
      RECT 7.78 2.1 8.03 2.36 ;
      RECT 5.505 3.635 5.765 3.895 ;
      RECT 7.8 3.125 7.805 3.335 ;
      RECT 7.805 3.13 7.815 3.33 ;
      RECT 7.755 3.125 7.8 3.35 ;
      RECT 7.745 3.125 7.755 3.37 ;
      RECT 7.726 3.125 7.745 3.375 ;
      RECT 7.64 3.125 7.726 3.372 ;
      RECT 7.61 3.127 7.64 3.37 ;
      RECT 7.555 3.137 7.61 3.368 ;
      RECT 7.49 3.151 7.555 3.366 ;
      RECT 7.485 3.159 7.49 3.365 ;
      RECT 7.47 3.162 7.485 3.363 ;
      RECT 7.405 3.172 7.47 3.359 ;
      RECT 7.357 3.186 7.405 3.36 ;
      RECT 7.271 3.203 7.357 3.374 ;
      RECT 7.185 3.224 7.271 3.391 ;
      RECT 7.165 3.237 7.185 3.401 ;
      RECT 7.12 3.245 7.165 3.408 ;
      RECT 7.085 3.253 7.12 3.416 ;
      RECT 7.051 3.261 7.085 3.424 ;
      RECT 6.965 3.275 7.051 3.436 ;
      RECT 6.93 3.292 6.965 3.448 ;
      RECT 6.921 3.301 6.93 3.452 ;
      RECT 6.835 3.319 6.921 3.469 ;
      RECT 6.776 3.346 6.835 3.496 ;
      RECT 6.69 3.373 6.776 3.524 ;
      RECT 6.67 3.395 6.69 3.544 ;
      RECT 6.61 3.41 6.67 3.56 ;
      RECT 6.6 3.422 6.61 3.573 ;
      RECT 6.595 3.427 6.6 3.576 ;
      RECT 6.585 3.43 6.595 3.579 ;
      RECT 6.58 3.432 6.585 3.582 ;
      RECT 6.55 3.44 6.58 3.589 ;
      RECT 6.535 3.447 6.55 3.597 ;
      RECT 6.525 3.452 6.535 3.601 ;
      RECT 6.52 3.455 6.525 3.604 ;
      RECT 6.51 3.457 6.52 3.607 ;
      RECT 6.475 3.467 6.51 3.616 ;
      RECT 6.4 3.49 6.475 3.638 ;
      RECT 6.38 3.508 6.4 3.656 ;
      RECT 6.35 3.515 6.38 3.666 ;
      RECT 6.33 3.523 6.35 3.676 ;
      RECT 6.32 3.529 6.33 3.683 ;
      RECT 6.301 3.534 6.32 3.689 ;
      RECT 6.215 3.554 6.301 3.709 ;
      RECT 6.2 3.574 6.215 3.728 ;
      RECT 6.155 3.586 6.2 3.739 ;
      RECT 6.09 3.607 6.155 3.762 ;
      RECT 6.05 3.627 6.09 3.783 ;
      RECT 6.04 3.637 6.05 3.793 ;
      RECT 5.99 3.649 6.04 3.804 ;
      RECT 5.97 3.665 5.99 3.816 ;
      RECT 5.94 3.675 5.97 3.822 ;
      RECT 5.93 3.68 5.94 3.824 ;
      RECT 5.861 3.681 5.93 3.83 ;
      RECT 5.775 3.683 5.861 3.84 ;
      RECT 5.765 3.684 5.775 3.845 ;
      RECT 7.035 3.71 7.225 3.92 ;
      RECT 7.025 3.715 7.235 3.913 ;
      RECT 7.01 3.715 7.235 3.878 ;
      RECT 6.93 3.6 7.19 3.86 ;
      RECT 5.845 3.13 6.03 3.425 ;
      RECT 5.835 3.13 6.03 3.423 ;
      RECT 5.82 3.13 6.035 3.418 ;
      RECT 5.82 3.13 6.04 3.415 ;
      RECT 5.815 3.13 6.04 3.413 ;
      RECT 5.81 3.385 6.04 3.403 ;
      RECT 5.815 3.13 6.075 3.39 ;
      RECT 5.775 2.165 6.035 2.425 ;
      RECT 5.585 2.09 5.671 2.423 ;
      RECT 5.56 2.094 5.715 2.419 ;
      RECT 5.671 2.086 5.715 2.419 ;
      RECT 5.671 2.087 5.72 2.418 ;
      RECT 5.585 2.092 5.735 2.417 ;
      RECT 5.56 2.1 5.775 2.416 ;
      RECT 5.555 2.095 5.735 2.411 ;
      RECT 5.545 2.11 5.775 2.318 ;
      RECT 5.545 2.162 5.975 2.318 ;
      RECT 5.545 2.155 5.955 2.318 ;
      RECT 5.545 2.142 5.925 2.318 ;
      RECT 5.545 2.13 5.865 2.318 ;
      RECT 5.545 2.115 5.84 2.318 ;
      RECT 4.745 2.745 4.88 3.04 ;
      RECT 5.005 2.768 5.01 2.955 ;
      RECT 5.725 2.665 5.87 2.9 ;
      RECT 5.885 2.665 5.89 2.89 ;
      RECT 5.92 2.676 5.925 2.87 ;
      RECT 5.915 2.668 5.92 2.875 ;
      RECT 5.895 2.665 5.915 2.88 ;
      RECT 5.89 2.665 5.895 2.888 ;
      RECT 5.88 2.665 5.885 2.893 ;
      RECT 5.87 2.665 5.88 2.898 ;
      RECT 5.7 2.667 5.725 2.9 ;
      RECT 5.65 2.674 5.7 2.9 ;
      RECT 5.645 2.679 5.65 2.9 ;
      RECT 5.606 2.684 5.645 2.901 ;
      RECT 5.52 2.696 5.606 2.902 ;
      RECT 5.511 2.706 5.52 2.902 ;
      RECT 5.425 2.715 5.511 2.904 ;
      RECT 5.401 2.725 5.425 2.906 ;
      RECT 5.315 2.736 5.401 2.907 ;
      RECT 5.285 2.747 5.315 2.909 ;
      RECT 5.255 2.752 5.285 2.911 ;
      RECT 5.23 2.758 5.255 2.914 ;
      RECT 5.215 2.763 5.23 2.915 ;
      RECT 5.17 2.769 5.215 2.915 ;
      RECT 5.165 2.774 5.17 2.916 ;
      RECT 5.145 2.774 5.165 2.918 ;
      RECT 5.125 2.772 5.145 2.923 ;
      RECT 5.09 2.771 5.125 2.93 ;
      RECT 5.06 2.77 5.09 2.94 ;
      RECT 5.01 2.769 5.06 2.95 ;
      RECT 4.92 2.766 5.005 3.04 ;
      RECT 4.895 2.76 4.92 3.04 ;
      RECT 4.88 2.75 4.895 3.04 ;
      RECT 4.695 2.745 4.745 2.96 ;
      RECT 4.685 2.75 4.695 2.95 ;
      RECT 4.925 3.225 5.185 3.485 ;
      RECT 4.925 3.225 5.215 3.378 ;
      RECT 4.925 3.225 5.25 3.363 ;
      RECT 5.18 3.145 5.37 3.355 ;
      RECT 5.17 3.15 5.38 3.348 ;
      RECT 5.135 3.22 5.38 3.348 ;
      RECT 5.165 3.162 5.185 3.485 ;
      RECT 5.15 3.21 5.38 3.348 ;
      RECT 5.155 3.182 5.185 3.485 ;
      RECT 4.235 2.25 4.305 3.355 ;
      RECT 4.97 2.355 5.23 2.615 ;
      RECT 4.55 2.401 4.565 2.61 ;
      RECT 4.886 2.414 4.97 2.565 ;
      RECT 4.8 2.411 4.886 2.565 ;
      RECT 4.761 2.409 4.8 2.565 ;
      RECT 4.675 2.407 4.761 2.565 ;
      RECT 4.615 2.405 4.675 2.576 ;
      RECT 4.58 2.403 4.615 2.594 ;
      RECT 4.565 2.401 4.58 2.605 ;
      RECT 4.535 2.401 4.55 2.618 ;
      RECT 4.525 2.401 4.535 2.623 ;
      RECT 4.5 2.4 4.525 2.628 ;
      RECT 4.485 2.395 4.5 2.634 ;
      RECT 4.48 2.388 4.485 2.639 ;
      RECT 4.455 2.379 4.48 2.645 ;
      RECT 4.41 2.358 4.455 2.658 ;
      RECT 4.4 2.342 4.41 2.668 ;
      RECT 4.385 2.335 4.4 2.678 ;
      RECT 4.375 2.328 4.385 2.695 ;
      RECT 4.37 2.325 4.375 2.725 ;
      RECT 4.365 2.323 4.37 2.755 ;
      RECT 4.36 2.321 4.365 2.792 ;
      RECT 4.345 2.317 4.36 2.859 ;
      RECT 4.345 3.15 4.355 3.35 ;
      RECT 4.34 2.313 4.345 2.985 ;
      RECT 4.34 3.137 4.345 3.355 ;
      RECT 4.335 2.311 4.34 3.07 ;
      RECT 4.335 3.127 4.34 3.355 ;
      RECT 4.32 2.282 4.335 3.355 ;
      RECT 4.305 2.255 4.32 3.355 ;
      RECT 4.23 2.25 4.235 2.605 ;
      RECT 4.23 2.66 4.235 3.355 ;
      RECT 4.215 2.25 4.23 2.583 ;
      RECT 4.225 2.682 4.23 3.355 ;
      RECT 4.215 2.722 4.225 3.355 ;
      RECT 4.18 2.25 4.215 2.525 ;
      RECT 4.21 2.757 4.215 3.355 ;
      RECT 4.195 2.812 4.21 3.355 ;
      RECT 4.19 2.877 4.195 3.355 ;
      RECT 4.175 2.925 4.19 3.355 ;
      RECT 4.15 2.25 4.18 2.48 ;
      RECT 4.17 2.98 4.175 3.355 ;
      RECT 4.155 3.04 4.17 3.355 ;
      RECT 4.15 3.088 4.155 3.353 ;
      RECT 4.145 2.25 4.15 2.473 ;
      RECT 4.145 3.12 4.15 3.348 ;
      RECT 4.12 2.25 4.145 2.465 ;
      RECT 4.11 2.255 4.12 2.455 ;
      RECT 4.325 3.53 4.345 3.77 ;
      RECT 3.555 3.46 3.56 3.67 ;
      RECT 4.835 3.533 4.845 3.728 ;
      RECT 4.83 3.523 4.835 3.731 ;
      RECT 4.75 3.52 4.83 3.754 ;
      RECT 4.746 3.52 4.75 3.776 ;
      RECT 4.66 3.52 4.746 3.786 ;
      RECT 4.645 3.52 4.66 3.794 ;
      RECT 4.616 3.521 4.645 3.792 ;
      RECT 4.53 3.526 4.616 3.788 ;
      RECT 4.517 3.53 4.53 3.784 ;
      RECT 4.431 3.53 4.517 3.78 ;
      RECT 4.345 3.53 4.431 3.774 ;
      RECT 4.261 3.53 4.325 3.768 ;
      RECT 4.175 3.53 4.261 3.763 ;
      RECT 4.155 3.53 4.175 3.759 ;
      RECT 4.095 3.525 4.155 3.756 ;
      RECT 4.067 3.519 4.095 3.753 ;
      RECT 3.981 3.514 4.067 3.749 ;
      RECT 3.895 3.508 3.981 3.743 ;
      RECT 3.82 3.49 3.895 3.738 ;
      RECT 3.785 3.467 3.82 3.734 ;
      RECT 3.775 3.457 3.785 3.733 ;
      RECT 3.72 3.455 3.775 3.732 ;
      RECT 3.645 3.455 3.72 3.728 ;
      RECT 3.635 3.455 3.645 3.723 ;
      RECT 3.62 3.455 3.635 3.715 ;
      RECT 3.57 3.457 3.62 3.693 ;
      RECT 3.56 3.46 3.57 3.673 ;
      RECT 3.55 3.465 3.555 3.668 ;
      RECT 3.545 3.47 3.55 3.663 ;
      RECT 3.67 2.635 3.93 2.895 ;
      RECT 3.67 2.65 3.95 2.86 ;
      RECT 3.67 2.655 3.96 2.855 ;
      RECT 1.655 2.115 1.915 2.375 ;
      RECT 1.645 2.145 1.915 2.355 ;
      RECT 3.565 2.06 3.825 2.32 ;
      RECT 3.56 2.135 3.565 2.321 ;
      RECT 3.535 2.14 3.56 2.323 ;
      RECT 3.52 2.147 3.535 2.326 ;
      RECT 3.46 2.165 3.52 2.331 ;
      RECT 3.43 2.185 3.46 2.338 ;
      RECT 3.405 2.193 3.43 2.343 ;
      RECT 3.38 2.201 3.405 2.345 ;
      RECT 3.362 2.205 3.38 2.344 ;
      RECT 3.276 2.203 3.362 2.344 ;
      RECT 3.19 2.201 3.276 2.344 ;
      RECT 3.104 2.199 3.19 2.343 ;
      RECT 3.018 2.197 3.104 2.343 ;
      RECT 2.932 2.195 3.018 2.343 ;
      RECT 2.846 2.193 2.932 2.343 ;
      RECT 2.76 2.191 2.846 2.342 ;
      RECT 2.742 2.19 2.76 2.342 ;
      RECT 2.656 2.189 2.742 2.342 ;
      RECT 2.57 2.187 2.656 2.342 ;
      RECT 2.484 2.186 2.57 2.341 ;
      RECT 2.398 2.185 2.484 2.341 ;
      RECT 2.312 2.183 2.398 2.341 ;
      RECT 2.226 2.182 2.312 2.341 ;
      RECT 2.14 2.18 2.226 2.34 ;
      RECT 2.116 2.178 2.14 2.34 ;
      RECT 2.03 2.171 2.116 2.34 ;
      RECT 2.001 2.163 2.03 2.34 ;
      RECT 1.915 2.155 2.001 2.34 ;
      RECT 1.635 2.152 1.645 2.35 ;
      RECT 3.14 3.115 3.145 3.465 ;
      RECT 2.91 3.205 3.05 3.465 ;
      RECT 3.385 2.89 3.43 3.1 ;
      RECT 3.44 2.901 3.45 3.095 ;
      RECT 3.43 2.893 3.44 3.1 ;
      RECT 3.365 2.89 3.385 3.105 ;
      RECT 3.335 2.89 3.365 3.128 ;
      RECT 3.325 2.89 3.335 3.153 ;
      RECT 3.32 2.89 3.325 3.163 ;
      RECT 3.265 2.89 3.32 3.203 ;
      RECT 3.26 2.89 3.265 3.243 ;
      RECT 3.255 2.892 3.26 3.248 ;
      RECT 3.24 2.902 3.255 3.259 ;
      RECT 3.195 2.96 3.24 3.295 ;
      RECT 3.185 3.015 3.195 3.329 ;
      RECT 3.17 3.042 3.185 3.345 ;
      RECT 3.16 3.069 3.17 3.465 ;
      RECT 3.145 3.092 3.16 3.465 ;
      RECT 3.135 3.132 3.14 3.465 ;
      RECT 3.13 3.142 3.135 3.465 ;
      RECT 3.125 3.157 3.13 3.465 ;
      RECT 3.115 3.162 3.125 3.465 ;
      RECT 3.05 3.185 3.115 3.465 ;
      RECT 2.55 2.68 2.74 2.89 ;
      RECT 1.125 2.605 1.385 2.865 ;
      RECT 1.475 2.6 1.57 2.81 ;
      RECT 1.45 2.615 1.46 2.81 ;
      RECT 2.74 2.687 2.75 2.885 ;
      RECT 2.54 2.687 2.55 2.885 ;
      RECT 2.525 2.702 2.54 2.875 ;
      RECT 2.52 2.71 2.525 2.868 ;
      RECT 2.51 2.713 2.52 2.865 ;
      RECT 2.475 2.712 2.51 2.863 ;
      RECT 2.446 2.708 2.475 2.86 ;
      RECT 2.36 2.703 2.446 2.857 ;
      RECT 2.3 2.697 2.36 2.853 ;
      RECT 2.271 2.693 2.3 2.85 ;
      RECT 2.185 2.685 2.271 2.847 ;
      RECT 2.176 2.679 2.185 2.845 ;
      RECT 2.09 2.674 2.176 2.843 ;
      RECT 2.067 2.669 2.09 2.84 ;
      RECT 1.981 2.663 2.067 2.837 ;
      RECT 1.895 2.654 1.981 2.832 ;
      RECT 1.885 2.649 1.895 2.83 ;
      RECT 1.866 2.648 1.885 2.829 ;
      RECT 1.78 2.643 1.866 2.825 ;
      RECT 1.76 2.638 1.78 2.821 ;
      RECT 1.7 2.633 1.76 2.818 ;
      RECT 1.675 2.623 1.7 2.816 ;
      RECT 1.67 2.616 1.675 2.815 ;
      RECT 1.66 2.607 1.67 2.814 ;
      RECT 1.656 2.6 1.66 2.814 ;
      RECT 1.57 2.6 1.656 2.812 ;
      RECT 1.46 2.607 1.475 2.81 ;
      RECT 1.445 2.617 1.45 2.81 ;
      RECT 1.425 2.62 1.445 2.807 ;
      RECT 1.395 2.62 1.425 2.803 ;
      RECT 1.385 2.62 1.395 2.803 ;
      RECT 2.3 3.115 2.56 3.375 ;
      RECT 2.23 3.125 2.56 3.335 ;
      RECT 2.22 3.132 2.56 3.33 ;
      RECT 1.64 3.12 1.9 3.38 ;
      RECT 1.64 3.16 2.005 3.37 ;
      RECT 1.64 3.162 2.01 3.369 ;
      RECT 1.64 3.17 2.015 3.366 ;
      RECT 0.565 2.245 0.665 3.77 ;
      RECT 0.755 3.385 0.805 3.645 ;
      RECT 0.75 2.258 0.755 2.445 ;
      RECT 0.745 3.366 0.755 3.645 ;
      RECT 0.745 2.255 0.75 2.453 ;
      RECT 0.73 2.249 0.745 2.46 ;
      RECT 0.74 3.354 0.745 3.728 ;
      RECT 0.73 3.342 0.74 3.765 ;
      RECT 0.72 2.245 0.73 2.467 ;
      RECT 0.72 3.327 0.73 3.77 ;
      RECT 0.715 2.245 0.72 2.475 ;
      RECT 0.695 3.297 0.72 3.77 ;
      RECT 0.675 2.245 0.715 2.523 ;
      RECT 0.685 3.257 0.695 3.77 ;
      RECT 0.675 3.212 0.685 3.77 ;
      RECT 0.67 2.245 0.675 2.593 ;
      RECT 0.67 3.17 0.675 3.77 ;
      RECT 0.665 2.245 0.67 3.07 ;
      RECT 0.665 3.152 0.67 3.77 ;
      RECT 0.555 2.248 0.565 3.77 ;
      RECT 0.54 2.255 0.555 3.766 ;
      RECT 0.535 2.265 0.54 3.761 ;
      RECT 0.53 2.465 0.535 3.653 ;
      RECT 0.525 2.55 0.53 3.205 ;
      RECT 0.01 8.575 89.605 8.88 ;
      RECT 78.21 2.225 78.47 2.485 ;
      RECT 60.29 2.225 60.55 2.485 ;
      RECT 42.37 2.225 42.63 2.485 ;
      RECT 24.455 2.225 24.715 2.485 ;
      RECT 6.535 2.225 6.795 2.485 ;
    LAYER mcon ;
      RECT 89.065 0.915 89.235 1.085 ;
      RECT 89.065 2.395 89.235 2.565 ;
      RECT 89.065 6.315 89.235 6.485 ;
      RECT 89.065 7.795 89.235 7.965 ;
      RECT 88.715 0.105 88.885 0.275 ;
      RECT 88.715 4.165 88.885 4.335 ;
      RECT 88.715 4.545 88.885 4.715 ;
      RECT 88.715 8.605 88.885 8.775 ;
      RECT 88.695 2.765 88.865 2.935 ;
      RECT 88.695 5.945 88.865 6.115 ;
      RECT 88.075 0.915 88.245 1.085 ;
      RECT 88.075 2.395 88.245 2.565 ;
      RECT 88.075 6.315 88.245 6.485 ;
      RECT 88.075 7.795 88.245 7.965 ;
      RECT 87.725 0.105 87.895 0.275 ;
      RECT 87.725 4.165 87.895 4.335 ;
      RECT 87.725 4.545 87.895 4.715 ;
      RECT 87.725 8.605 87.895 8.775 ;
      RECT 87.705 2.765 87.875 2.935 ;
      RECT 87.705 5.945 87.875 6.115 ;
      RECT 87.02 0.105 87.19 0.275 ;
      RECT 87.02 4.165 87.19 4.335 ;
      RECT 87.02 4.545 87.19 4.715 ;
      RECT 87.02 8.605 87.19 8.775 ;
      RECT 86.71 2.025 86.88 2.195 ;
      RECT 86.71 6.685 86.88 6.855 ;
      RECT 86.34 0.105 86.51 0.275 ;
      RECT 86.34 8.605 86.51 8.775 ;
      RECT 86.28 0.915 86.45 1.085 ;
      RECT 86.28 1.655 86.45 1.825 ;
      RECT 86.28 7.055 86.45 7.225 ;
      RECT 86.28 7.795 86.45 7.965 ;
      RECT 85.905 2.395 86.075 2.565 ;
      RECT 85.905 6.315 86.075 6.485 ;
      RECT 85.66 0.105 85.83 0.275 ;
      RECT 85.66 8.605 85.83 8.775 ;
      RECT 84.98 0.105 85.15 0.275 ;
      RECT 84.98 8.605 85.15 8.775 ;
      RECT 84.91 2.765 85.08 2.935 ;
      RECT 84.91 5.945 85.08 6.115 ;
      RECT 83.7 1.565 83.87 1.735 ;
      RECT 83.7 4.285 83.87 4.455 ;
      RECT 83.24 1.565 83.41 1.735 ;
      RECT 83.24 4.285 83.41 4.455 ;
      RECT 82.845 2.905 83.015 3.075 ;
      RECT 82.78 1.565 82.95 1.735 ;
      RECT 82.78 4.285 82.95 4.455 ;
      RECT 82.635 2.245 82.805 2.415 ;
      RECT 82.32 1.565 82.49 1.735 ;
      RECT 82.32 3.155 82.49 3.325 ;
      RECT 82.32 4.285 82.49 4.455 ;
      RECT 81.935 2.75 82.105 2.92 ;
      RECT 81.86 1.565 82.03 1.735 ;
      RECT 81.86 4.285 82.03 4.455 ;
      RECT 81.72 3.315 81.89 3.485 ;
      RECT 81.7 3.715 81.87 3.885 ;
      RECT 81.525 2.27 81.695 2.44 ;
      RECT 81.4 1.565 81.57 1.735 ;
      RECT 81.4 4.285 81.57 4.455 ;
      RECT 81.03 3.25 81.2 3.42 ;
      RECT 80.94 1.565 81.11 1.735 ;
      RECT 80.94 4.285 81.11 4.455 ;
      RECT 80.705 2.935 80.875 3.105 ;
      RECT 80.64 3.715 80.81 3.885 ;
      RECT 80.48 1.565 80.65 1.735 ;
      RECT 80.48 4.285 80.65 4.455 ;
      RECT 80.24 3.7 80.41 3.87 ;
      RECT 80.2 2.185 80.37 2.355 ;
      RECT 80.02 1.565 80.19 1.735 ;
      RECT 80.02 4.285 80.19 4.455 ;
      RECT 79.56 1.565 79.73 1.735 ;
      RECT 79.56 4.285 79.73 4.455 ;
      RECT 79.3 2.685 79.47 2.855 ;
      RECT 79.3 3.145 79.47 3.315 ;
      RECT 79.3 3.66 79.47 3.83 ;
      RECT 79.185 2.22 79.355 2.39 ;
      RECT 79.1 1.565 79.27 1.735 ;
      RECT 79.1 4.285 79.27 4.455 ;
      RECT 78.72 3.73 78.89 3.9 ;
      RECT 78.64 1.565 78.81 1.735 ;
      RECT 78.64 4.285 78.81 4.455 ;
      RECT 78.24 2.26 78.41 2.43 ;
      RECT 78.18 1.565 78.35 1.735 ;
      RECT 78.18 4.285 78.35 4.455 ;
      RECT 78.025 2.635 78.195 2.805 ;
      RECT 77.72 1.565 77.89 1.735 ;
      RECT 77.72 4.285 77.89 4.455 ;
      RECT 77.525 3.235 77.695 3.405 ;
      RECT 77.41 2.685 77.58 2.855 ;
      RECT 77.26 1.565 77.43 1.735 ;
      RECT 77.26 4.285 77.43 4.455 ;
      RECT 77.24 2.135 77.41 2.305 ;
      RECT 76.865 3.165 77.035 3.335 ;
      RECT 76.8 1.565 76.97 1.735 ;
      RECT 76.8 4.285 76.97 4.455 ;
      RECT 76.38 2.765 76.55 2.935 ;
      RECT 76.34 1.565 76.51 1.735 ;
      RECT 76.34 4.285 76.51 4.455 ;
      RECT 76.33 3.54 76.5 3.71 ;
      RECT 75.88 1.565 76.05 1.735 ;
      RECT 75.88 4.285 76.05 4.455 ;
      RECT 75.84 3.165 76.01 3.335 ;
      RECT 75.805 2.27 75.975 2.44 ;
      RECT 75.445 2.67 75.615 2.84 ;
      RECT 75.42 1.565 75.59 1.735 ;
      RECT 75.42 4.285 75.59 4.455 ;
      RECT 75.24 3.48 75.41 3.65 ;
      RECT 74.96 1.565 75.13 1.735 ;
      RECT 74.96 4.285 75.13 4.455 ;
      RECT 74.935 2.91 75.105 3.08 ;
      RECT 74.5 1.565 74.67 1.735 ;
      RECT 74.5 4.285 74.67 4.455 ;
      RECT 74.235 2.7 74.405 2.87 ;
      RECT 74.04 1.565 74.21 1.735 ;
      RECT 74.04 4.285 74.21 4.455 ;
      RECT 73.915 3.145 74.085 3.315 ;
      RECT 73.58 1.565 73.75 1.735 ;
      RECT 73.58 4.285 73.75 4.455 ;
      RECT 73.5 3.18 73.67 3.35 ;
      RECT 73.33 2.165 73.5 2.335 ;
      RECT 73.155 2.62 73.325 2.79 ;
      RECT 73.12 1.565 73.29 1.735 ;
      RECT 73.12 4.285 73.29 4.455 ;
      RECT 72.66 1.565 72.83 1.735 ;
      RECT 72.66 4.285 72.83 4.455 ;
      RECT 72.235 2.27 72.405 2.44 ;
      RECT 72.23 3.585 72.4 3.755 ;
      RECT 72.2 1.565 72.37 1.735 ;
      RECT 72.2 4.285 72.37 4.455 ;
      RECT 71.145 0.915 71.315 1.085 ;
      RECT 71.145 2.395 71.315 2.565 ;
      RECT 71.145 6.315 71.315 6.485 ;
      RECT 71.145 7.795 71.315 7.965 ;
      RECT 70.795 0.105 70.965 0.275 ;
      RECT 70.795 4.165 70.965 4.335 ;
      RECT 70.795 4.545 70.965 4.715 ;
      RECT 70.795 8.605 70.965 8.775 ;
      RECT 70.775 2.765 70.945 2.935 ;
      RECT 70.775 5.945 70.945 6.115 ;
      RECT 70.155 0.915 70.325 1.085 ;
      RECT 70.155 2.395 70.325 2.565 ;
      RECT 70.155 6.315 70.325 6.485 ;
      RECT 70.155 7.795 70.325 7.965 ;
      RECT 69.805 0.105 69.975 0.275 ;
      RECT 69.805 4.165 69.975 4.335 ;
      RECT 69.805 4.545 69.975 4.715 ;
      RECT 69.805 8.605 69.975 8.775 ;
      RECT 69.785 2.765 69.955 2.935 ;
      RECT 69.785 5.945 69.955 6.115 ;
      RECT 69.1 0.105 69.27 0.275 ;
      RECT 69.1 4.165 69.27 4.335 ;
      RECT 69.1 4.545 69.27 4.715 ;
      RECT 69.1 8.605 69.27 8.775 ;
      RECT 68.79 2.025 68.96 2.195 ;
      RECT 68.79 6.685 68.96 6.855 ;
      RECT 68.42 0.105 68.59 0.275 ;
      RECT 68.42 8.605 68.59 8.775 ;
      RECT 68.36 0.915 68.53 1.085 ;
      RECT 68.36 1.655 68.53 1.825 ;
      RECT 68.36 7.055 68.53 7.225 ;
      RECT 68.36 7.795 68.53 7.965 ;
      RECT 67.985 2.395 68.155 2.565 ;
      RECT 67.985 6.315 68.155 6.485 ;
      RECT 67.74 0.105 67.91 0.275 ;
      RECT 67.74 8.605 67.91 8.775 ;
      RECT 67.06 0.105 67.23 0.275 ;
      RECT 67.06 8.605 67.23 8.775 ;
      RECT 66.99 2.765 67.16 2.935 ;
      RECT 66.99 5.945 67.16 6.115 ;
      RECT 65.78 1.565 65.95 1.735 ;
      RECT 65.78 4.285 65.95 4.455 ;
      RECT 65.32 1.565 65.49 1.735 ;
      RECT 65.32 4.285 65.49 4.455 ;
      RECT 64.925 2.905 65.095 3.075 ;
      RECT 64.86 1.565 65.03 1.735 ;
      RECT 64.86 4.285 65.03 4.455 ;
      RECT 64.715 2.245 64.885 2.415 ;
      RECT 64.4 1.565 64.57 1.735 ;
      RECT 64.4 3.155 64.57 3.325 ;
      RECT 64.4 4.285 64.57 4.455 ;
      RECT 64.015 2.75 64.185 2.92 ;
      RECT 63.94 1.565 64.11 1.735 ;
      RECT 63.94 4.285 64.11 4.455 ;
      RECT 63.8 3.315 63.97 3.485 ;
      RECT 63.78 3.715 63.95 3.885 ;
      RECT 63.605 2.27 63.775 2.44 ;
      RECT 63.48 1.565 63.65 1.735 ;
      RECT 63.48 4.285 63.65 4.455 ;
      RECT 63.11 3.25 63.28 3.42 ;
      RECT 63.02 1.565 63.19 1.735 ;
      RECT 63.02 4.285 63.19 4.455 ;
      RECT 62.785 2.935 62.955 3.105 ;
      RECT 62.72 3.715 62.89 3.885 ;
      RECT 62.56 1.565 62.73 1.735 ;
      RECT 62.56 4.285 62.73 4.455 ;
      RECT 62.32 3.7 62.49 3.87 ;
      RECT 62.28 2.185 62.45 2.355 ;
      RECT 62.1 1.565 62.27 1.735 ;
      RECT 62.1 4.285 62.27 4.455 ;
      RECT 61.64 1.565 61.81 1.735 ;
      RECT 61.64 4.285 61.81 4.455 ;
      RECT 61.38 2.685 61.55 2.855 ;
      RECT 61.38 3.145 61.55 3.315 ;
      RECT 61.38 3.66 61.55 3.83 ;
      RECT 61.265 2.22 61.435 2.39 ;
      RECT 61.18 1.565 61.35 1.735 ;
      RECT 61.18 4.285 61.35 4.455 ;
      RECT 60.8 3.73 60.97 3.9 ;
      RECT 60.72 1.565 60.89 1.735 ;
      RECT 60.72 4.285 60.89 4.455 ;
      RECT 60.32 2.26 60.49 2.43 ;
      RECT 60.26 1.565 60.43 1.735 ;
      RECT 60.26 4.285 60.43 4.455 ;
      RECT 60.105 2.635 60.275 2.805 ;
      RECT 59.8 1.565 59.97 1.735 ;
      RECT 59.8 4.285 59.97 4.455 ;
      RECT 59.605 3.235 59.775 3.405 ;
      RECT 59.49 2.685 59.66 2.855 ;
      RECT 59.34 1.565 59.51 1.735 ;
      RECT 59.34 4.285 59.51 4.455 ;
      RECT 59.32 2.135 59.49 2.305 ;
      RECT 58.945 3.165 59.115 3.335 ;
      RECT 58.88 1.565 59.05 1.735 ;
      RECT 58.88 4.285 59.05 4.455 ;
      RECT 58.46 2.765 58.63 2.935 ;
      RECT 58.42 1.565 58.59 1.735 ;
      RECT 58.42 4.285 58.59 4.455 ;
      RECT 58.41 3.54 58.58 3.71 ;
      RECT 57.96 1.565 58.13 1.735 ;
      RECT 57.96 4.285 58.13 4.455 ;
      RECT 57.92 3.165 58.09 3.335 ;
      RECT 57.885 2.27 58.055 2.44 ;
      RECT 57.525 2.67 57.695 2.84 ;
      RECT 57.5 1.565 57.67 1.735 ;
      RECT 57.5 4.285 57.67 4.455 ;
      RECT 57.32 3.48 57.49 3.65 ;
      RECT 57.04 1.565 57.21 1.735 ;
      RECT 57.04 4.285 57.21 4.455 ;
      RECT 57.015 2.91 57.185 3.08 ;
      RECT 56.58 1.565 56.75 1.735 ;
      RECT 56.58 4.285 56.75 4.455 ;
      RECT 56.315 2.7 56.485 2.87 ;
      RECT 56.12 1.565 56.29 1.735 ;
      RECT 56.12 4.285 56.29 4.455 ;
      RECT 55.995 3.145 56.165 3.315 ;
      RECT 55.66 1.565 55.83 1.735 ;
      RECT 55.66 4.285 55.83 4.455 ;
      RECT 55.58 3.18 55.75 3.35 ;
      RECT 55.41 2.165 55.58 2.335 ;
      RECT 55.235 2.62 55.405 2.79 ;
      RECT 55.2 1.565 55.37 1.735 ;
      RECT 55.2 4.285 55.37 4.455 ;
      RECT 54.74 1.565 54.91 1.735 ;
      RECT 54.74 4.285 54.91 4.455 ;
      RECT 54.315 2.27 54.485 2.44 ;
      RECT 54.31 3.585 54.48 3.755 ;
      RECT 54.28 1.565 54.45 1.735 ;
      RECT 54.28 4.285 54.45 4.455 ;
      RECT 53.225 0.915 53.395 1.085 ;
      RECT 53.225 2.395 53.395 2.565 ;
      RECT 53.225 6.315 53.395 6.485 ;
      RECT 53.225 7.795 53.395 7.965 ;
      RECT 52.875 0.105 53.045 0.275 ;
      RECT 52.875 4.165 53.045 4.335 ;
      RECT 52.875 4.545 53.045 4.715 ;
      RECT 52.875 8.605 53.045 8.775 ;
      RECT 52.855 2.765 53.025 2.935 ;
      RECT 52.855 5.945 53.025 6.115 ;
      RECT 52.235 0.915 52.405 1.085 ;
      RECT 52.235 2.395 52.405 2.565 ;
      RECT 52.235 6.315 52.405 6.485 ;
      RECT 52.235 7.795 52.405 7.965 ;
      RECT 51.885 0.105 52.055 0.275 ;
      RECT 51.885 4.165 52.055 4.335 ;
      RECT 51.885 4.545 52.055 4.715 ;
      RECT 51.885 8.605 52.055 8.775 ;
      RECT 51.865 2.765 52.035 2.935 ;
      RECT 51.865 5.945 52.035 6.115 ;
      RECT 51.18 0.105 51.35 0.275 ;
      RECT 51.18 4.165 51.35 4.335 ;
      RECT 51.18 4.545 51.35 4.715 ;
      RECT 51.18 8.605 51.35 8.775 ;
      RECT 50.87 2.025 51.04 2.195 ;
      RECT 50.87 6.685 51.04 6.855 ;
      RECT 50.5 0.105 50.67 0.275 ;
      RECT 50.5 8.605 50.67 8.775 ;
      RECT 50.44 0.915 50.61 1.085 ;
      RECT 50.44 1.655 50.61 1.825 ;
      RECT 50.44 7.055 50.61 7.225 ;
      RECT 50.44 7.795 50.61 7.965 ;
      RECT 50.065 2.395 50.235 2.565 ;
      RECT 50.065 6.315 50.235 6.485 ;
      RECT 49.82 0.105 49.99 0.275 ;
      RECT 49.82 8.605 49.99 8.775 ;
      RECT 49.14 0.105 49.31 0.275 ;
      RECT 49.14 8.605 49.31 8.775 ;
      RECT 49.07 2.765 49.24 2.935 ;
      RECT 49.07 5.945 49.24 6.115 ;
      RECT 47.86 1.565 48.03 1.735 ;
      RECT 47.86 4.285 48.03 4.455 ;
      RECT 47.4 1.565 47.57 1.735 ;
      RECT 47.4 4.285 47.57 4.455 ;
      RECT 47.005 2.905 47.175 3.075 ;
      RECT 46.94 1.565 47.11 1.735 ;
      RECT 46.94 4.285 47.11 4.455 ;
      RECT 46.795 2.245 46.965 2.415 ;
      RECT 46.48 1.565 46.65 1.735 ;
      RECT 46.48 3.155 46.65 3.325 ;
      RECT 46.48 4.285 46.65 4.455 ;
      RECT 46.095 2.75 46.265 2.92 ;
      RECT 46.02 1.565 46.19 1.735 ;
      RECT 46.02 4.285 46.19 4.455 ;
      RECT 45.88 3.315 46.05 3.485 ;
      RECT 45.86 3.715 46.03 3.885 ;
      RECT 45.685 2.27 45.855 2.44 ;
      RECT 45.56 1.565 45.73 1.735 ;
      RECT 45.56 4.285 45.73 4.455 ;
      RECT 45.19 3.25 45.36 3.42 ;
      RECT 45.1 1.565 45.27 1.735 ;
      RECT 45.1 4.285 45.27 4.455 ;
      RECT 44.865 2.935 45.035 3.105 ;
      RECT 44.8 3.715 44.97 3.885 ;
      RECT 44.64 1.565 44.81 1.735 ;
      RECT 44.64 4.285 44.81 4.455 ;
      RECT 44.4 3.7 44.57 3.87 ;
      RECT 44.36 2.185 44.53 2.355 ;
      RECT 44.18 1.565 44.35 1.735 ;
      RECT 44.18 4.285 44.35 4.455 ;
      RECT 43.72 1.565 43.89 1.735 ;
      RECT 43.72 4.285 43.89 4.455 ;
      RECT 43.46 2.685 43.63 2.855 ;
      RECT 43.46 3.145 43.63 3.315 ;
      RECT 43.46 3.66 43.63 3.83 ;
      RECT 43.345 2.22 43.515 2.39 ;
      RECT 43.26 1.565 43.43 1.735 ;
      RECT 43.26 4.285 43.43 4.455 ;
      RECT 42.88 3.73 43.05 3.9 ;
      RECT 42.8 1.565 42.97 1.735 ;
      RECT 42.8 4.285 42.97 4.455 ;
      RECT 42.4 2.26 42.57 2.43 ;
      RECT 42.34 1.565 42.51 1.735 ;
      RECT 42.34 4.285 42.51 4.455 ;
      RECT 42.185 2.635 42.355 2.805 ;
      RECT 41.88 1.565 42.05 1.735 ;
      RECT 41.88 4.285 42.05 4.455 ;
      RECT 41.685 3.235 41.855 3.405 ;
      RECT 41.57 2.685 41.74 2.855 ;
      RECT 41.42 1.565 41.59 1.735 ;
      RECT 41.42 4.285 41.59 4.455 ;
      RECT 41.4 2.135 41.57 2.305 ;
      RECT 41.025 3.165 41.195 3.335 ;
      RECT 40.96 1.565 41.13 1.735 ;
      RECT 40.96 4.285 41.13 4.455 ;
      RECT 40.54 2.765 40.71 2.935 ;
      RECT 40.5 1.565 40.67 1.735 ;
      RECT 40.5 4.285 40.67 4.455 ;
      RECT 40.49 3.54 40.66 3.71 ;
      RECT 40.04 1.565 40.21 1.735 ;
      RECT 40.04 4.285 40.21 4.455 ;
      RECT 40 3.165 40.17 3.335 ;
      RECT 39.965 2.27 40.135 2.44 ;
      RECT 39.605 2.67 39.775 2.84 ;
      RECT 39.58 1.565 39.75 1.735 ;
      RECT 39.58 4.285 39.75 4.455 ;
      RECT 39.4 3.48 39.57 3.65 ;
      RECT 39.12 1.565 39.29 1.735 ;
      RECT 39.12 4.285 39.29 4.455 ;
      RECT 39.095 2.91 39.265 3.08 ;
      RECT 38.66 1.565 38.83 1.735 ;
      RECT 38.66 4.285 38.83 4.455 ;
      RECT 38.395 2.7 38.565 2.87 ;
      RECT 38.2 1.565 38.37 1.735 ;
      RECT 38.2 4.285 38.37 4.455 ;
      RECT 38.075 3.145 38.245 3.315 ;
      RECT 37.74 1.565 37.91 1.735 ;
      RECT 37.74 4.285 37.91 4.455 ;
      RECT 37.66 3.18 37.83 3.35 ;
      RECT 37.49 2.165 37.66 2.335 ;
      RECT 37.315 2.62 37.485 2.79 ;
      RECT 37.28 1.565 37.45 1.735 ;
      RECT 37.28 4.285 37.45 4.455 ;
      RECT 36.82 1.565 36.99 1.735 ;
      RECT 36.82 4.285 36.99 4.455 ;
      RECT 36.395 2.27 36.565 2.44 ;
      RECT 36.39 3.585 36.56 3.755 ;
      RECT 36.36 1.565 36.53 1.735 ;
      RECT 36.36 4.285 36.53 4.455 ;
      RECT 35.31 0.915 35.48 1.085 ;
      RECT 35.31 2.395 35.48 2.565 ;
      RECT 35.31 6.315 35.48 6.485 ;
      RECT 35.31 7.795 35.48 7.965 ;
      RECT 34.96 0.105 35.13 0.275 ;
      RECT 34.96 4.165 35.13 4.335 ;
      RECT 34.96 4.545 35.13 4.715 ;
      RECT 34.96 8.605 35.13 8.775 ;
      RECT 34.94 2.765 35.11 2.935 ;
      RECT 34.94 5.945 35.11 6.115 ;
      RECT 34.32 0.915 34.49 1.085 ;
      RECT 34.32 2.395 34.49 2.565 ;
      RECT 34.32 6.315 34.49 6.485 ;
      RECT 34.32 7.795 34.49 7.965 ;
      RECT 33.97 0.105 34.14 0.275 ;
      RECT 33.97 4.165 34.14 4.335 ;
      RECT 33.97 4.545 34.14 4.715 ;
      RECT 33.97 8.605 34.14 8.775 ;
      RECT 33.95 2.765 34.12 2.935 ;
      RECT 33.95 5.945 34.12 6.115 ;
      RECT 33.265 0.105 33.435 0.275 ;
      RECT 33.265 4.165 33.435 4.335 ;
      RECT 33.265 4.545 33.435 4.715 ;
      RECT 33.265 8.605 33.435 8.775 ;
      RECT 32.955 2.025 33.125 2.195 ;
      RECT 32.955 6.685 33.125 6.855 ;
      RECT 32.585 0.105 32.755 0.275 ;
      RECT 32.585 8.605 32.755 8.775 ;
      RECT 32.525 0.915 32.695 1.085 ;
      RECT 32.525 1.655 32.695 1.825 ;
      RECT 32.525 7.055 32.695 7.225 ;
      RECT 32.525 7.795 32.695 7.965 ;
      RECT 32.15 2.395 32.32 2.565 ;
      RECT 32.15 6.315 32.32 6.485 ;
      RECT 31.905 0.105 32.075 0.275 ;
      RECT 31.905 8.605 32.075 8.775 ;
      RECT 31.225 0.105 31.395 0.275 ;
      RECT 31.225 8.605 31.395 8.775 ;
      RECT 31.155 2.765 31.325 2.935 ;
      RECT 31.155 5.945 31.325 6.115 ;
      RECT 29.945 1.565 30.115 1.735 ;
      RECT 29.945 4.285 30.115 4.455 ;
      RECT 29.485 1.565 29.655 1.735 ;
      RECT 29.485 4.285 29.655 4.455 ;
      RECT 29.09 2.905 29.26 3.075 ;
      RECT 29.025 1.565 29.195 1.735 ;
      RECT 29.025 4.285 29.195 4.455 ;
      RECT 28.88 2.245 29.05 2.415 ;
      RECT 28.565 1.565 28.735 1.735 ;
      RECT 28.565 3.155 28.735 3.325 ;
      RECT 28.565 4.285 28.735 4.455 ;
      RECT 28.18 2.75 28.35 2.92 ;
      RECT 28.105 1.565 28.275 1.735 ;
      RECT 28.105 4.285 28.275 4.455 ;
      RECT 27.965 3.315 28.135 3.485 ;
      RECT 27.945 3.715 28.115 3.885 ;
      RECT 27.77 2.27 27.94 2.44 ;
      RECT 27.645 1.565 27.815 1.735 ;
      RECT 27.645 4.285 27.815 4.455 ;
      RECT 27.275 3.25 27.445 3.42 ;
      RECT 27.185 1.565 27.355 1.735 ;
      RECT 27.185 4.285 27.355 4.455 ;
      RECT 26.95 2.935 27.12 3.105 ;
      RECT 26.885 3.715 27.055 3.885 ;
      RECT 26.725 1.565 26.895 1.735 ;
      RECT 26.725 4.285 26.895 4.455 ;
      RECT 26.485 3.7 26.655 3.87 ;
      RECT 26.445 2.185 26.615 2.355 ;
      RECT 26.265 1.565 26.435 1.735 ;
      RECT 26.265 4.285 26.435 4.455 ;
      RECT 25.805 1.565 25.975 1.735 ;
      RECT 25.805 4.285 25.975 4.455 ;
      RECT 25.545 2.685 25.715 2.855 ;
      RECT 25.545 3.145 25.715 3.315 ;
      RECT 25.545 3.66 25.715 3.83 ;
      RECT 25.43 2.22 25.6 2.39 ;
      RECT 25.345 1.565 25.515 1.735 ;
      RECT 25.345 4.285 25.515 4.455 ;
      RECT 24.965 3.73 25.135 3.9 ;
      RECT 24.885 1.565 25.055 1.735 ;
      RECT 24.885 4.285 25.055 4.455 ;
      RECT 24.485 2.26 24.655 2.43 ;
      RECT 24.425 1.565 24.595 1.735 ;
      RECT 24.425 4.285 24.595 4.455 ;
      RECT 24.27 2.635 24.44 2.805 ;
      RECT 23.965 1.565 24.135 1.735 ;
      RECT 23.965 4.285 24.135 4.455 ;
      RECT 23.77 3.235 23.94 3.405 ;
      RECT 23.655 2.685 23.825 2.855 ;
      RECT 23.505 1.565 23.675 1.735 ;
      RECT 23.505 4.285 23.675 4.455 ;
      RECT 23.485 2.135 23.655 2.305 ;
      RECT 23.11 3.165 23.28 3.335 ;
      RECT 23.045 1.565 23.215 1.735 ;
      RECT 23.045 4.285 23.215 4.455 ;
      RECT 22.625 2.765 22.795 2.935 ;
      RECT 22.585 1.565 22.755 1.735 ;
      RECT 22.585 4.285 22.755 4.455 ;
      RECT 22.575 3.54 22.745 3.71 ;
      RECT 22.125 1.565 22.295 1.735 ;
      RECT 22.125 4.285 22.295 4.455 ;
      RECT 22.085 3.165 22.255 3.335 ;
      RECT 22.05 2.27 22.22 2.44 ;
      RECT 21.69 2.67 21.86 2.84 ;
      RECT 21.665 1.565 21.835 1.735 ;
      RECT 21.665 4.285 21.835 4.455 ;
      RECT 21.485 3.48 21.655 3.65 ;
      RECT 21.205 1.565 21.375 1.735 ;
      RECT 21.205 4.285 21.375 4.455 ;
      RECT 21.18 2.91 21.35 3.08 ;
      RECT 20.745 1.565 20.915 1.735 ;
      RECT 20.745 4.285 20.915 4.455 ;
      RECT 20.48 2.7 20.65 2.87 ;
      RECT 20.285 1.565 20.455 1.735 ;
      RECT 20.285 4.285 20.455 4.455 ;
      RECT 20.16 3.145 20.33 3.315 ;
      RECT 19.825 1.565 19.995 1.735 ;
      RECT 19.825 4.285 19.995 4.455 ;
      RECT 19.745 3.18 19.915 3.35 ;
      RECT 19.575 2.165 19.745 2.335 ;
      RECT 19.4 2.62 19.57 2.79 ;
      RECT 19.365 1.565 19.535 1.735 ;
      RECT 19.365 4.285 19.535 4.455 ;
      RECT 18.905 1.565 19.075 1.735 ;
      RECT 18.905 4.285 19.075 4.455 ;
      RECT 18.48 2.27 18.65 2.44 ;
      RECT 18.475 3.585 18.645 3.755 ;
      RECT 18.445 1.565 18.615 1.735 ;
      RECT 18.445 4.285 18.615 4.455 ;
      RECT 17.39 0.915 17.56 1.085 ;
      RECT 17.39 2.395 17.56 2.565 ;
      RECT 17.39 6.315 17.56 6.485 ;
      RECT 17.39 7.795 17.56 7.965 ;
      RECT 17.04 0.105 17.21 0.275 ;
      RECT 17.04 4.165 17.21 4.335 ;
      RECT 17.04 4.545 17.21 4.715 ;
      RECT 17.04 8.605 17.21 8.775 ;
      RECT 17.02 2.765 17.19 2.935 ;
      RECT 17.02 5.945 17.19 6.115 ;
      RECT 16.4 0.915 16.57 1.085 ;
      RECT 16.4 2.395 16.57 2.565 ;
      RECT 16.4 6.315 16.57 6.485 ;
      RECT 16.4 7.795 16.57 7.965 ;
      RECT 16.05 0.105 16.22 0.275 ;
      RECT 16.05 4.165 16.22 4.335 ;
      RECT 16.05 4.545 16.22 4.715 ;
      RECT 16.05 8.605 16.22 8.775 ;
      RECT 16.03 2.765 16.2 2.935 ;
      RECT 16.03 5.945 16.2 6.115 ;
      RECT 15.345 0.105 15.515 0.275 ;
      RECT 15.345 4.165 15.515 4.335 ;
      RECT 15.345 4.545 15.515 4.715 ;
      RECT 15.345 8.605 15.515 8.775 ;
      RECT 15.035 2.025 15.205 2.195 ;
      RECT 15.035 6.685 15.205 6.855 ;
      RECT 14.665 0.105 14.835 0.275 ;
      RECT 14.665 8.605 14.835 8.775 ;
      RECT 14.605 0.915 14.775 1.085 ;
      RECT 14.605 1.655 14.775 1.825 ;
      RECT 14.605 7.055 14.775 7.225 ;
      RECT 14.605 7.795 14.775 7.965 ;
      RECT 14.23 2.395 14.4 2.565 ;
      RECT 14.23 6.315 14.4 6.485 ;
      RECT 13.985 0.105 14.155 0.275 ;
      RECT 13.985 8.605 14.155 8.775 ;
      RECT 13.305 0.105 13.475 0.275 ;
      RECT 13.305 8.605 13.475 8.775 ;
      RECT 13.235 2.765 13.405 2.935 ;
      RECT 13.235 5.945 13.405 6.115 ;
      RECT 12.025 1.565 12.195 1.735 ;
      RECT 12.025 4.285 12.195 4.455 ;
      RECT 11.565 1.565 11.735 1.735 ;
      RECT 11.565 4.285 11.735 4.455 ;
      RECT 11.17 2.905 11.34 3.075 ;
      RECT 11.105 1.565 11.275 1.735 ;
      RECT 11.105 4.285 11.275 4.455 ;
      RECT 10.96 2.245 11.13 2.415 ;
      RECT 10.645 1.565 10.815 1.735 ;
      RECT 10.645 3.155 10.815 3.325 ;
      RECT 10.645 4.285 10.815 4.455 ;
      RECT 10.26 2.75 10.43 2.92 ;
      RECT 10.185 1.565 10.355 1.735 ;
      RECT 10.185 4.285 10.355 4.455 ;
      RECT 10.045 3.315 10.215 3.485 ;
      RECT 10.025 3.715 10.195 3.885 ;
      RECT 9.85 2.27 10.02 2.44 ;
      RECT 9.725 1.565 9.895 1.735 ;
      RECT 9.725 4.285 9.895 4.455 ;
      RECT 9.355 3.25 9.525 3.42 ;
      RECT 9.265 1.565 9.435 1.735 ;
      RECT 9.265 4.285 9.435 4.455 ;
      RECT 9.03 2.935 9.2 3.105 ;
      RECT 8.965 3.715 9.135 3.885 ;
      RECT 8.805 1.565 8.975 1.735 ;
      RECT 8.805 4.285 8.975 4.455 ;
      RECT 8.565 3.7 8.735 3.87 ;
      RECT 8.525 2.185 8.695 2.355 ;
      RECT 8.345 1.565 8.515 1.735 ;
      RECT 8.345 4.285 8.515 4.455 ;
      RECT 7.885 1.565 8.055 1.735 ;
      RECT 7.885 4.285 8.055 4.455 ;
      RECT 7.625 2.685 7.795 2.855 ;
      RECT 7.625 3.145 7.795 3.315 ;
      RECT 7.625 3.66 7.795 3.83 ;
      RECT 7.51 2.22 7.68 2.39 ;
      RECT 7.425 1.565 7.595 1.735 ;
      RECT 7.425 4.285 7.595 4.455 ;
      RECT 7.045 3.73 7.215 3.9 ;
      RECT 6.965 1.565 7.135 1.735 ;
      RECT 6.965 4.285 7.135 4.455 ;
      RECT 6.565 2.26 6.735 2.43 ;
      RECT 6.505 1.565 6.675 1.735 ;
      RECT 6.505 4.285 6.675 4.455 ;
      RECT 6.35 2.635 6.52 2.805 ;
      RECT 6.045 1.565 6.215 1.735 ;
      RECT 6.045 4.285 6.215 4.455 ;
      RECT 5.85 3.235 6.02 3.405 ;
      RECT 5.735 2.685 5.905 2.855 ;
      RECT 5.585 1.565 5.755 1.735 ;
      RECT 5.585 4.285 5.755 4.455 ;
      RECT 5.565 2.135 5.735 2.305 ;
      RECT 5.19 3.165 5.36 3.335 ;
      RECT 5.125 1.565 5.295 1.735 ;
      RECT 5.125 4.285 5.295 4.455 ;
      RECT 4.705 2.765 4.875 2.935 ;
      RECT 4.665 1.565 4.835 1.735 ;
      RECT 4.665 4.285 4.835 4.455 ;
      RECT 4.655 3.54 4.825 3.71 ;
      RECT 4.205 1.565 4.375 1.735 ;
      RECT 4.205 4.285 4.375 4.455 ;
      RECT 4.165 3.165 4.335 3.335 ;
      RECT 4.13 2.27 4.3 2.44 ;
      RECT 3.77 2.67 3.94 2.84 ;
      RECT 3.745 1.565 3.915 1.735 ;
      RECT 3.745 4.285 3.915 4.455 ;
      RECT 3.565 3.48 3.735 3.65 ;
      RECT 3.285 1.565 3.455 1.735 ;
      RECT 3.285 4.285 3.455 4.455 ;
      RECT 3.26 2.91 3.43 3.08 ;
      RECT 2.825 1.565 2.995 1.735 ;
      RECT 2.825 4.285 2.995 4.455 ;
      RECT 2.56 2.7 2.73 2.87 ;
      RECT 2.365 1.565 2.535 1.735 ;
      RECT 2.365 4.285 2.535 4.455 ;
      RECT 2.24 3.145 2.41 3.315 ;
      RECT 1.905 1.565 2.075 1.735 ;
      RECT 1.905 4.285 2.075 4.455 ;
      RECT 1.825 3.18 1.995 3.35 ;
      RECT 1.655 2.165 1.825 2.335 ;
      RECT 1.48 2.62 1.65 2.79 ;
      RECT 1.445 1.565 1.615 1.735 ;
      RECT 1.445 4.285 1.615 4.455 ;
      RECT 0.985 1.565 1.155 1.735 ;
      RECT 0.985 4.285 1.155 4.455 ;
      RECT 0.56 2.27 0.73 2.44 ;
      RECT 0.555 3.585 0.725 3.755 ;
      RECT 0.525 1.565 0.695 1.735 ;
      RECT 0.525 4.285 0.695 4.455 ;
    LAYER li ;
      RECT 83.105 0 83.275 2.235 ;
      RECT 82.145 0 82.315 2.235 ;
      RECT 81.185 0 81.355 2.235 ;
      RECT 80.665 0 80.835 2.235 ;
      RECT 79.705 0 79.875 2.235 ;
      RECT 78.705 0 78.875 2.235 ;
      RECT 77.745 0 77.915 2.235 ;
      RECT 76.265 0 76.435 2.235 ;
      RECT 74.345 0 74.515 2.235 ;
      RECT 72.865 0 73.035 2.235 ;
      RECT 65.185 0 65.355 2.235 ;
      RECT 64.225 0 64.395 2.235 ;
      RECT 63.265 0 63.435 2.235 ;
      RECT 62.745 0 62.915 2.235 ;
      RECT 61.785 0 61.955 2.235 ;
      RECT 60.785 0 60.955 2.235 ;
      RECT 59.825 0 59.995 2.235 ;
      RECT 58.345 0 58.515 2.235 ;
      RECT 56.425 0 56.595 2.235 ;
      RECT 54.945 0 55.115 2.235 ;
      RECT 47.265 0 47.435 2.235 ;
      RECT 46.305 0 46.475 2.235 ;
      RECT 45.345 0 45.515 2.235 ;
      RECT 44.825 0 44.995 2.235 ;
      RECT 43.865 0 44.035 2.235 ;
      RECT 42.865 0 43.035 2.235 ;
      RECT 41.905 0 42.075 2.235 ;
      RECT 40.425 0 40.595 2.235 ;
      RECT 38.505 0 38.675 2.235 ;
      RECT 37.025 0 37.195 2.235 ;
      RECT 29.35 0 29.52 2.235 ;
      RECT 28.39 0 28.56 2.235 ;
      RECT 27.43 0 27.6 2.235 ;
      RECT 26.91 0 27.08 2.235 ;
      RECT 25.95 0 26.12 2.235 ;
      RECT 24.95 0 25.12 2.235 ;
      RECT 23.99 0 24.16 2.235 ;
      RECT 22.51 0 22.68 2.235 ;
      RECT 20.59 0 20.76 2.235 ;
      RECT 19.11 0 19.28 2.235 ;
      RECT 11.43 0 11.6 2.235 ;
      RECT 10.47 0 10.64 2.235 ;
      RECT 9.51 0 9.68 2.235 ;
      RECT 8.99 0 9.16 2.235 ;
      RECT 8.03 0 8.2 2.235 ;
      RECT 7.03 0 7.2 2.235 ;
      RECT 6.07 0 6.24 2.235 ;
      RECT 4.59 0 4.76 2.235 ;
      RECT 2.67 0 2.84 2.235 ;
      RECT 1.19 0 1.36 2.235 ;
      RECT 72.055 0 84.015 1.735 ;
      RECT 54.135 0 66.095 1.735 ;
      RECT 36.215 0 48.175 1.735 ;
      RECT 18.3 0 30.26 1.735 ;
      RECT 0.38 0 12.34 1.735 ;
      RECT 72.05 0 84.015 1.68 ;
      RECT 54.13 0 66.095 1.68 ;
      RECT 36.21 0 48.175 1.68 ;
      RECT 18.295 0 30.26 1.68 ;
      RECT 0.375 0 12.34 1.68 ;
      RECT 88.635 0 88.805 0.935 ;
      RECT 87.645 0 87.815 0.935 ;
      RECT 84.9 0 85.07 0.935 ;
      RECT 70.715 0 70.885 0.935 ;
      RECT 69.725 0 69.895 0.935 ;
      RECT 66.98 0 67.15 0.935 ;
      RECT 52.795 0 52.965 0.935 ;
      RECT 51.805 0 51.975 0.935 ;
      RECT 49.06 0 49.23 0.935 ;
      RECT 34.88 0 35.05 0.935 ;
      RECT 33.89 0 34.06 0.935 ;
      RECT 31.145 0 31.315 0.935 ;
      RECT 16.96 0 17.13 0.935 ;
      RECT 15.97 0 16.14 0.935 ;
      RECT 13.225 0 13.395 0.935 ;
      RECT 0.005 0 89.605 0.305 ;
      RECT 88.635 3.405 88.805 5.475 ;
      RECT 87.645 3.405 87.815 5.475 ;
      RECT 84.9 3.405 85.07 5.475 ;
      RECT 70.715 3.405 70.885 5.475 ;
      RECT 69.725 3.405 69.895 5.475 ;
      RECT 66.98 3.405 67.15 5.475 ;
      RECT 52.795 3.405 52.965 5.475 ;
      RECT 51.805 3.405 51.975 5.475 ;
      RECT 49.06 3.405 49.23 5.475 ;
      RECT 34.88 3.405 35.05 5.475 ;
      RECT 33.89 3.405 34.06 5.475 ;
      RECT 31.145 3.405 31.315 5.475 ;
      RECT 16.96 3.405 17.13 5.475 ;
      RECT 15.97 3.405 16.14 5.475 ;
      RECT 13.225 3.405 13.395 5.475 ;
      RECT 0.005 4.285 89.605 4.745 ;
      RECT 83.645 4.135 89.605 4.745 ;
      RECT 82.145 3.785 82.315 4.745 ;
      RECT 79.705 3.785 79.875 4.745 ;
      RECT 77.745 3.785 77.915 4.745 ;
      RECT 76.785 3.785 76.955 4.745 ;
      RECT 74.825 3.785 74.995 4.745 ;
      RECT 73.825 3.785 73.995 4.745 ;
      RECT 72.865 3.785 73.035 4.745 ;
      RECT 65.725 4.135 71.685 4.745 ;
      RECT 64.225 3.785 64.395 4.745 ;
      RECT 61.785 3.785 61.955 4.745 ;
      RECT 59.825 3.785 59.995 4.745 ;
      RECT 58.865 3.785 59.035 4.745 ;
      RECT 56.905 3.785 57.075 4.745 ;
      RECT 55.905 3.785 56.075 4.745 ;
      RECT 54.945 3.785 55.115 4.745 ;
      RECT 47.805 4.135 53.765 4.745 ;
      RECT 46.305 3.785 46.475 4.745 ;
      RECT 43.865 3.785 44.035 4.745 ;
      RECT 41.905 3.785 42.075 4.745 ;
      RECT 40.945 3.785 41.115 4.745 ;
      RECT 38.985 3.785 39.155 4.745 ;
      RECT 37.985 3.785 38.155 4.745 ;
      RECT 37.025 3.785 37.195 4.745 ;
      RECT 29.89 4.135 35.85 4.745 ;
      RECT 28.39 3.785 28.56 4.745 ;
      RECT 25.95 3.785 26.12 4.745 ;
      RECT 23.99 3.785 24.16 4.745 ;
      RECT 23.03 3.785 23.2 4.745 ;
      RECT 21.07 3.785 21.24 4.745 ;
      RECT 20.07 3.785 20.24 4.745 ;
      RECT 19.11 3.785 19.28 4.745 ;
      RECT 11.97 4.135 17.93 4.745 ;
      RECT 10.47 3.785 10.64 4.745 ;
      RECT 8.03 3.785 8.2 4.745 ;
      RECT 6.07 3.785 6.24 4.745 ;
      RECT 5.11 3.785 5.28 4.745 ;
      RECT 3.15 3.785 3.32 4.745 ;
      RECT 2.15 3.785 2.32 4.745 ;
      RECT 1.19 3.785 1.36 4.745 ;
      RECT 0.01 8.575 89.605 8.88 ;
      RECT 88.635 7.945 88.805 8.88 ;
      RECT 87.645 7.945 87.815 8.88 ;
      RECT 84.9 7.945 85.07 8.88 ;
      RECT 70.715 7.945 70.885 8.88 ;
      RECT 69.725 7.945 69.895 8.88 ;
      RECT 66.98 7.945 67.15 8.88 ;
      RECT 52.795 7.945 52.965 8.88 ;
      RECT 51.805 7.945 51.975 8.88 ;
      RECT 49.06 7.945 49.23 8.88 ;
      RECT 34.88 7.945 35.05 8.88 ;
      RECT 33.89 7.945 34.06 8.88 ;
      RECT 31.145 7.945 31.315 8.88 ;
      RECT 16.96 7.945 17.13 8.88 ;
      RECT 15.97 7.945 16.14 8.88 ;
      RECT 13.225 7.945 13.395 8.88 ;
      RECT 88.695 1.74 88.865 2.935 ;
      RECT 88.695 1.74 89.16 1.91 ;
      RECT 88.695 6.97 89.16 7.14 ;
      RECT 88.695 5.945 88.865 7.14 ;
      RECT 87.705 1.74 87.875 2.935 ;
      RECT 87.705 1.74 88.17 1.91 ;
      RECT 87.705 6.97 88.17 7.14 ;
      RECT 87.705 5.945 87.875 7.14 ;
      RECT 85.85 2.635 86.02 3.865 ;
      RECT 85.905 0.855 86.075 2.805 ;
      RECT 85.85 0.575 86.02 1.025 ;
      RECT 85.85 7.855 86.02 8.305 ;
      RECT 85.905 6.075 86.075 8.025 ;
      RECT 85.85 5.015 86.02 6.245 ;
      RECT 85.33 0.575 85.5 3.865 ;
      RECT 85.33 2.075 85.735 2.405 ;
      RECT 85.33 1.235 85.735 1.565 ;
      RECT 85.33 5.015 85.5 8.305 ;
      RECT 85.33 7.315 85.735 7.645 ;
      RECT 85.33 6.475 85.735 6.805 ;
      RECT 83.43 3.392 83.445 3.443 ;
      RECT 83.425 3.372 83.43 3.49 ;
      RECT 83.41 3.362 83.425 3.558 ;
      RECT 83.385 3.342 83.41 3.613 ;
      RECT 83.345 3.327 83.385 3.633 ;
      RECT 83.3 3.321 83.345 3.661 ;
      RECT 83.23 3.311 83.3 3.678 ;
      RECT 83.21 3.303 83.23 3.678 ;
      RECT 83.15 3.297 83.21 3.67 ;
      RECT 83.091 3.288 83.15 3.658 ;
      RECT 83.005 3.277 83.091 3.641 ;
      RECT 82.983 3.268 83.005 3.629 ;
      RECT 82.897 3.261 82.983 3.616 ;
      RECT 82.811 3.248 82.897 3.597 ;
      RECT 82.725 3.236 82.811 3.577 ;
      RECT 82.695 3.225 82.725 3.564 ;
      RECT 82.645 3.211 82.695 3.556 ;
      RECT 82.625 3.2 82.645 3.548 ;
      RECT 82.576 3.189 82.625 3.54 ;
      RECT 82.49 3.168 82.576 3.525 ;
      RECT 82.445 3.155 82.49 3.51 ;
      RECT 82.4 3.155 82.445 3.49 ;
      RECT 82.345 3.155 82.4 3.425 ;
      RECT 82.32 3.155 82.345 3.348 ;
      RECT 82.845 2.892 83.015 3.075 ;
      RECT 82.845 2.892 83.03 3.033 ;
      RECT 82.845 2.892 83.035 2.975 ;
      RECT 82.905 2.66 83.04 2.951 ;
      RECT 82.905 2.664 83.045 2.934 ;
      RECT 82.85 2.827 83.045 2.934 ;
      RECT 82.875 2.672 83.015 3.075 ;
      RECT 82.875 2.676 83.055 2.875 ;
      RECT 82.86 2.762 83.055 2.875 ;
      RECT 82.87 2.692 83.015 3.075 ;
      RECT 82.87 2.695 83.065 2.788 ;
      RECT 82.865 2.712 83.065 2.788 ;
      RECT 82.635 1.932 82.805 2.415 ;
      RECT 82.63 1.927 82.78 2.405 ;
      RECT 82.63 1.934 82.81 2.399 ;
      RECT 82.62 1.928 82.78 2.378 ;
      RECT 82.62 1.944 82.825 2.337 ;
      RECT 82.59 1.929 82.78 2.3 ;
      RECT 82.59 1.959 82.835 2.24 ;
      RECT 82.585 1.931 82.78 2.238 ;
      RECT 82.565 1.94 82.81 2.195 ;
      RECT 82.54 1.956 82.825 2.107 ;
      RECT 82.54 1.975 82.85 2.098 ;
      RECT 82.535 2.012 82.85 2.05 ;
      RECT 82.54 1.992 82.855 2.018 ;
      RECT 82.635 1.926 82.745 2.415 ;
      RECT 82.721 1.925 82.745 2.415 ;
      RECT 81.955 2.71 81.96 2.921 ;
      RECT 82.555 2.71 82.56 2.895 ;
      RECT 82.62 2.75 82.625 2.863 ;
      RECT 82.615 2.742 82.62 2.869 ;
      RECT 82.61 2.732 82.615 2.877 ;
      RECT 82.605 2.722 82.61 2.886 ;
      RECT 82.6 2.712 82.605 2.89 ;
      RECT 82.56 2.71 82.6 2.893 ;
      RECT 82.532 2.709 82.555 2.897 ;
      RECT 82.446 2.706 82.532 2.904 ;
      RECT 82.36 2.702 82.446 2.915 ;
      RECT 82.34 2.7 82.36 2.921 ;
      RECT 82.322 2.699 82.34 2.924 ;
      RECT 82.236 2.697 82.322 2.931 ;
      RECT 82.15 2.692 82.236 2.944 ;
      RECT 82.131 2.689 82.15 2.949 ;
      RECT 82.045 2.687 82.131 2.94 ;
      RECT 82.035 2.687 82.045 2.933 ;
      RECT 81.96 2.7 82.035 2.927 ;
      RECT 81.945 2.711 81.955 2.921 ;
      RECT 81.935 2.713 81.945 2.92 ;
      RECT 81.925 2.717 81.935 2.916 ;
      RECT 81.92 2.72 81.925 2.91 ;
      RECT 81.91 2.722 81.92 2.904 ;
      RECT 81.905 2.725 81.91 2.898 ;
      RECT 81.885 3.311 81.89 3.515 ;
      RECT 81.87 3.298 81.885 3.608 ;
      RECT 81.855 3.279 81.87 3.885 ;
      RECT 81.82 3.245 81.855 3.885 ;
      RECT 81.816 3.215 81.82 3.885 ;
      RECT 81.73 3.097 81.816 3.885 ;
      RECT 81.72 2.972 81.73 3.885 ;
      RECT 81.705 2.94 81.72 3.885 ;
      RECT 81.7 2.915 81.705 3.885 ;
      RECT 81.695 2.905 81.7 3.841 ;
      RECT 81.68 2.877 81.695 3.746 ;
      RECT 81.665 2.843 81.68 3.645 ;
      RECT 81.66 2.821 81.665 3.598 ;
      RECT 81.655 2.81 81.66 3.568 ;
      RECT 81.65 2.8 81.655 3.534 ;
      RECT 81.64 2.787 81.65 3.502 ;
      RECT 81.615 2.763 81.64 3.428 ;
      RECT 81.61 2.743 81.615 3.353 ;
      RECT 81.605 2.737 81.61 3.328 ;
      RECT 81.6 2.732 81.605 3.293 ;
      RECT 81.595 2.727 81.6 3.268 ;
      RECT 81.59 2.725 81.595 3.248 ;
      RECT 81.585 2.725 81.59 3.233 ;
      RECT 81.58 2.725 81.585 3.193 ;
      RECT 81.57 2.725 81.58 3.165 ;
      RECT 81.56 2.725 81.57 3.11 ;
      RECT 81.545 2.725 81.56 3.048 ;
      RECT 81.54 2.724 81.545 2.993 ;
      RECT 81.525 2.723 81.54 2.973 ;
      RECT 81.465 2.721 81.525 2.947 ;
      RECT 81.43 2.722 81.465 2.927 ;
      RECT 81.425 2.724 81.43 2.917 ;
      RECT 81.415 2.743 81.425 2.907 ;
      RECT 81.41 2.77 81.415 2.838 ;
      RECT 81.525 2.195 81.695 2.44 ;
      RECT 81.56 1.966 81.695 2.44 ;
      RECT 81.56 1.968 81.705 2.435 ;
      RECT 81.56 1.97 81.73 2.423 ;
      RECT 81.56 1.973 81.755 2.405 ;
      RECT 81.56 1.978 81.805 2.378 ;
      RECT 81.56 1.983 81.825 2.343 ;
      RECT 81.54 1.985 81.835 2.318 ;
      RECT 81.53 2.08 81.835 2.318 ;
      RECT 81.56 1.965 81.67 2.44 ;
      RECT 81.57 1.962 81.665 2.44 ;
      RECT 81.09 3.227 81.28 3.585 ;
      RECT 81.09 3.239 81.315 3.584 ;
      RECT 81.09 3.267 81.335 3.582 ;
      RECT 81.09 3.292 81.34 3.581 ;
      RECT 81.09 3.35 81.355 3.58 ;
      RECT 81.075 3.223 81.235 3.565 ;
      RECT 81.055 3.232 81.28 3.518 ;
      RECT 81.03 3.243 81.315 3.455 ;
      RECT 81.03 3.327 81.35 3.455 ;
      RECT 81.03 3.302 81.345 3.455 ;
      RECT 81.09 3.218 81.235 3.585 ;
      RECT 81.176 3.217 81.235 3.585 ;
      RECT 81.176 3.216 81.22 3.585 ;
      RECT 80.875 2.732 80.88 3.11 ;
      RECT 80.87 2.7 80.875 3.11 ;
      RECT 80.865 2.672 80.87 3.11 ;
      RECT 80.86 2.652 80.865 3.11 ;
      RECT 80.805 2.635 80.86 3.11 ;
      RECT 80.765 2.62 80.805 3.11 ;
      RECT 80.71 2.607 80.765 3.11 ;
      RECT 80.675 2.598 80.71 3.11 ;
      RECT 80.671 2.596 80.675 3.109 ;
      RECT 80.585 2.592 80.671 3.092 ;
      RECT 80.5 2.584 80.585 3.055 ;
      RECT 80.49 2.58 80.5 3.028 ;
      RECT 80.48 2.58 80.49 3.01 ;
      RECT 80.47 2.582 80.48 2.993 ;
      RECT 80.465 2.587 80.47 2.979 ;
      RECT 80.46 2.591 80.465 2.966 ;
      RECT 80.45 2.596 80.46 2.95 ;
      RECT 80.435 2.61 80.45 2.925 ;
      RECT 80.43 2.616 80.435 2.905 ;
      RECT 80.425 2.618 80.43 2.898 ;
      RECT 80.42 2.622 80.425 2.773 ;
      RECT 80.6 3.422 80.845 3.885 ;
      RECT 80.52 3.395 80.84 3.881 ;
      RECT 80.45 3.43 80.845 3.874 ;
      RECT 80.24 3.685 80.845 3.87 ;
      RECT 80.42 3.453 80.845 3.87 ;
      RECT 80.26 3.645 80.845 3.87 ;
      RECT 80.41 3.465 80.845 3.87 ;
      RECT 80.295 3.582 80.845 3.87 ;
      RECT 80.35 3.507 80.845 3.87 ;
      RECT 80.6 3.372 80.84 3.885 ;
      RECT 80.63 3.365 80.84 3.885 ;
      RECT 80.62 3.367 80.84 3.885 ;
      RECT 80.63 3.362 80.76 3.885 ;
      RECT 80.185 1.925 80.271 2.364 ;
      RECT 80.18 1.925 80.271 2.362 ;
      RECT 80.18 1.925 80.34 2.361 ;
      RECT 80.18 1.925 80.37 2.358 ;
      RECT 80.165 1.932 80.37 2.349 ;
      RECT 80.165 1.932 80.375 2.345 ;
      RECT 80.16 1.942 80.375 2.338 ;
      RECT 80.155 1.947 80.375 2.313 ;
      RECT 80.155 1.947 80.39 2.295 ;
      RECT 80.18 1.925 80.41 2.21 ;
      RECT 80.15 1.952 80.41 2.208 ;
      RECT 80.16 1.945 80.415 2.146 ;
      RECT 80.15 2.067 80.42 2.129 ;
      RECT 80.135 1.962 80.415 2.08 ;
      RECT 80.13 1.972 80.415 1.98 ;
      RECT 80.21 2.743 80.215 2.82 ;
      RECT 80.2 2.737 80.21 3.01 ;
      RECT 80.19 2.729 80.2 3.031 ;
      RECT 80.18 2.72 80.19 3.053 ;
      RECT 80.175 2.715 80.18 3.07 ;
      RECT 80.135 2.715 80.175 3.11 ;
      RECT 80.115 2.715 80.135 3.165 ;
      RECT 80.11 2.715 80.115 3.193 ;
      RECT 80.1 2.715 80.11 3.208 ;
      RECT 80.065 2.715 80.1 3.25 ;
      RECT 80.06 2.715 80.065 3.293 ;
      RECT 80.05 2.715 80.06 3.308 ;
      RECT 80.035 2.715 80.05 3.328 ;
      RECT 80.02 2.715 80.035 3.355 ;
      RECT 80.015 2.716 80.02 3.373 ;
      RECT 79.995 2.717 80.015 3.38 ;
      RECT 79.94 2.718 79.995 3.4 ;
      RECT 79.93 2.719 79.94 3.414 ;
      RECT 79.925 2.722 79.93 3.413 ;
      RECT 79.885 2.795 79.925 3.411 ;
      RECT 79.87 2.875 79.885 3.409 ;
      RECT 79.845 2.93 79.87 3.407 ;
      RECT 79.83 2.995 79.845 3.406 ;
      RECT 79.785 3.027 79.83 3.403 ;
      RECT 79.7 3.05 79.785 3.398 ;
      RECT 79.675 3.07 79.7 3.393 ;
      RECT 79.605 3.075 79.675 3.389 ;
      RECT 79.585 3.077 79.605 3.386 ;
      RECT 79.5 3.088 79.585 3.38 ;
      RECT 79.495 3.099 79.5 3.375 ;
      RECT 79.485 3.101 79.495 3.375 ;
      RECT 79.45 3.105 79.485 3.373 ;
      RECT 79.4 3.115 79.45 3.36 ;
      RECT 79.38 3.123 79.4 3.345 ;
      RECT 79.3 3.135 79.38 3.328 ;
      RECT 79.465 2.685 79.635 2.895 ;
      RECT 79.581 2.681 79.635 2.895 ;
      RECT 79.386 2.685 79.635 2.886 ;
      RECT 79.386 2.685 79.64 2.875 ;
      RECT 79.3 2.685 79.64 2.866 ;
      RECT 79.3 2.693 79.65 2.81 ;
      RECT 79.3 2.705 79.655 2.723 ;
      RECT 79.3 2.712 79.66 2.715 ;
      RECT 79.495 2.683 79.635 2.895 ;
      RECT 79.25 3.628 79.495 3.96 ;
      RECT 79.245 3.62 79.25 3.957 ;
      RECT 79.215 3.64 79.495 3.938 ;
      RECT 79.195 3.672 79.495 3.911 ;
      RECT 79.245 3.625 79.422 3.957 ;
      RECT 79.245 3.622 79.336 3.957 ;
      RECT 79.185 1.97 79.355 2.39 ;
      RECT 79.18 1.97 79.355 2.388 ;
      RECT 79.18 1.97 79.38 2.378 ;
      RECT 79.18 1.97 79.4 2.353 ;
      RECT 79.175 1.97 79.4 2.348 ;
      RECT 79.175 1.97 79.41 2.338 ;
      RECT 79.175 1.97 79.415 2.333 ;
      RECT 79.175 1.975 79.42 2.328 ;
      RECT 79.175 2.007 79.435 2.318 ;
      RECT 79.175 2.077 79.46 2.301 ;
      RECT 79.155 2.077 79.46 2.293 ;
      RECT 79.155 2.137 79.47 2.27 ;
      RECT 79.155 2.177 79.48 2.215 ;
      RECT 79.14 1.97 79.415 2.195 ;
      RECT 79.13 1.985 79.42 2.093 ;
      RECT 78.72 3.375 78.89 3.9 ;
      RECT 78.715 3.375 78.89 3.893 ;
      RECT 78.705 3.375 78.895 3.858 ;
      RECT 78.7 3.385 78.895 3.83 ;
      RECT 78.695 3.405 78.895 3.813 ;
      RECT 78.705 3.38 78.9 3.803 ;
      RECT 78.69 3.425 78.9 3.795 ;
      RECT 78.685 3.445 78.9 3.78 ;
      RECT 78.68 3.475 78.9 3.77 ;
      RECT 78.67 3.52 78.9 3.745 ;
      RECT 78.7 3.39 78.905 3.728 ;
      RECT 78.665 3.572 78.905 3.723 ;
      RECT 78.7 3.4 78.91 3.693 ;
      RECT 78.66 3.605 78.91 3.69 ;
      RECT 78.655 3.63 78.91 3.67 ;
      RECT 78.695 3.417 78.92 3.61 ;
      RECT 78.69 3.439 78.93 3.503 ;
      RECT 78.64 2.686 78.655 2.955 ;
      RECT 78.595 2.67 78.64 3 ;
      RECT 78.59 2.658 78.595 3.05 ;
      RECT 78.58 2.654 78.59 3.083 ;
      RECT 78.575 2.651 78.58 3.111 ;
      RECT 78.56 2.653 78.575 3.153 ;
      RECT 78.555 2.657 78.56 3.193 ;
      RECT 78.535 2.662 78.555 3.245 ;
      RECT 78.531 2.667 78.535 3.302 ;
      RECT 78.445 2.686 78.531 3.339 ;
      RECT 78.435 2.707 78.445 3.375 ;
      RECT 78.43 2.715 78.435 3.376 ;
      RECT 78.425 2.757 78.43 3.377 ;
      RECT 78.41 2.845 78.425 3.378 ;
      RECT 78.4 2.995 78.41 3.38 ;
      RECT 78.395 3.04 78.4 3.382 ;
      RECT 78.36 3.082 78.395 3.385 ;
      RECT 78.355 3.1 78.36 3.388 ;
      RECT 78.278 3.106 78.355 3.394 ;
      RECT 78.192 3.12 78.278 3.407 ;
      RECT 78.106 3.134 78.192 3.421 ;
      RECT 78.02 3.148 78.106 3.434 ;
      RECT 77.96 3.16 78.02 3.446 ;
      RECT 77.935 3.167 77.96 3.453 ;
      RECT 77.921 3.17 77.935 3.458 ;
      RECT 77.835 3.178 77.921 3.474 ;
      RECT 77.83 3.185 77.835 3.489 ;
      RECT 77.806 3.185 77.83 3.496 ;
      RECT 77.72 3.188 77.806 3.524 ;
      RECT 77.635 3.192 77.72 3.568 ;
      RECT 77.57 3.196 77.635 3.605 ;
      RECT 77.545 3.199 77.57 3.621 ;
      RECT 77.47 3.212 77.545 3.625 ;
      RECT 77.445 3.23 77.47 3.629 ;
      RECT 77.435 3.237 77.445 3.631 ;
      RECT 77.42 3.24 77.435 3.632 ;
      RECT 77.36 3.252 77.42 3.636 ;
      RECT 77.35 3.266 77.36 3.64 ;
      RECT 77.295 3.276 77.35 3.628 ;
      RECT 77.27 3.297 77.295 3.611 ;
      RECT 77.25 3.317 77.27 3.602 ;
      RECT 77.245 3.33 77.25 3.597 ;
      RECT 77.23 3.342 77.245 3.593 ;
      RECT 78.465 1.997 78.47 2.02 ;
      RECT 78.46 1.988 78.465 2.06 ;
      RECT 78.455 1.986 78.46 2.103 ;
      RECT 78.45 1.977 78.455 2.138 ;
      RECT 78.445 1.967 78.45 2.21 ;
      RECT 78.44 1.957 78.445 2.275 ;
      RECT 78.435 1.954 78.44 2.315 ;
      RECT 78.41 1.948 78.435 2.405 ;
      RECT 78.375 1.936 78.41 2.43 ;
      RECT 78.365 1.927 78.375 2.43 ;
      RECT 78.23 1.925 78.24 2.413 ;
      RECT 78.22 1.925 78.23 2.38 ;
      RECT 78.215 1.925 78.22 2.355 ;
      RECT 78.21 1.925 78.215 2.343 ;
      RECT 78.205 1.925 78.21 2.325 ;
      RECT 78.195 1.925 78.205 2.29 ;
      RECT 78.19 1.927 78.195 2.268 ;
      RECT 78.185 1.933 78.19 2.253 ;
      RECT 78.18 1.939 78.185 2.238 ;
      RECT 78.165 1.951 78.18 2.211 ;
      RECT 78.16 1.962 78.165 2.179 ;
      RECT 78.155 1.972 78.16 2.163 ;
      RECT 78.145 1.98 78.155 2.132 ;
      RECT 78.14 1.99 78.145 2.106 ;
      RECT 78.135 2.047 78.14 2.089 ;
      RECT 78.24 1.925 78.365 2.43 ;
      RECT 77.955 2.612 78.215 2.91 ;
      RECT 77.95 2.619 78.215 2.908 ;
      RECT 77.955 2.614 78.23 2.903 ;
      RECT 77.945 2.627 78.23 2.9 ;
      RECT 77.945 2.632 78.235 2.893 ;
      RECT 77.94 2.64 78.235 2.89 ;
      RECT 77.94 2.657 78.24 2.688 ;
      RECT 77.955 2.609 78.186 2.91 ;
      RECT 78.01 2.608 78.186 2.91 ;
      RECT 78.01 2.605 78.1 2.91 ;
      RECT 78.01 2.602 78.096 2.91 ;
      RECT 77.7 2.875 77.705 2.888 ;
      RECT 77.695 2.842 77.7 2.893 ;
      RECT 77.69 2.797 77.695 2.9 ;
      RECT 77.685 2.752 77.69 2.908 ;
      RECT 77.68 2.72 77.685 2.916 ;
      RECT 77.675 2.68 77.68 2.917 ;
      RECT 77.66 2.66 77.675 2.919 ;
      RECT 77.585 2.642 77.66 2.931 ;
      RECT 77.575 2.635 77.585 2.942 ;
      RECT 77.57 2.635 77.575 2.944 ;
      RECT 77.54 2.641 77.57 2.948 ;
      RECT 77.5 2.654 77.54 2.948 ;
      RECT 77.475 2.665 77.5 2.934 ;
      RECT 77.46 2.671 77.475 2.917 ;
      RECT 77.45 2.673 77.46 2.908 ;
      RECT 77.445 2.674 77.45 2.903 ;
      RECT 77.44 2.675 77.445 2.898 ;
      RECT 77.435 2.676 77.44 2.895 ;
      RECT 77.41 2.681 77.435 2.885 ;
      RECT 77.4 2.697 77.41 2.872 ;
      RECT 77.395 2.717 77.4 2.867 ;
      RECT 77.405 2.11 77.41 2.306 ;
      RECT 77.39 2.074 77.405 2.308 ;
      RECT 77.38 2.056 77.39 2.313 ;
      RECT 77.37 2.042 77.38 2.317 ;
      RECT 77.325 2.026 77.37 2.327 ;
      RECT 77.32 2.016 77.325 2.336 ;
      RECT 77.275 2.005 77.32 2.342 ;
      RECT 77.27 1.993 77.275 2.349 ;
      RECT 77.255 1.988 77.27 2.353 ;
      RECT 77.24 1.98 77.255 2.358 ;
      RECT 77.23 1.973 77.24 2.363 ;
      RECT 77.22 1.97 77.23 2.368 ;
      RECT 77.21 1.97 77.22 2.369 ;
      RECT 77.205 1.967 77.21 2.368 ;
      RECT 77.17 1.962 77.195 2.367 ;
      RECT 77.146 1.958 77.17 2.366 ;
      RECT 77.06 1.949 77.146 2.363 ;
      RECT 77.045 1.941 77.06 2.36 ;
      RECT 77.023 1.94 77.045 2.359 ;
      RECT 76.937 1.94 77.023 2.357 ;
      RECT 76.851 1.94 76.937 2.355 ;
      RECT 76.765 1.94 76.851 2.352 ;
      RECT 76.755 1.94 76.765 2.343 ;
      RECT 76.725 1.94 76.755 2.303 ;
      RECT 76.715 1.95 76.725 2.258 ;
      RECT 76.71 1.99 76.715 2.243 ;
      RECT 76.705 2.005 76.71 2.23 ;
      RECT 76.675 2.085 76.705 2.192 ;
      RECT 77.195 1.965 77.205 2.368 ;
      RECT 77.02 2.73 77.035 3.335 ;
      RECT 77.025 2.725 77.035 3.335 ;
      RECT 77.19 2.725 77.195 2.908 ;
      RECT 77.18 2.725 77.19 2.938 ;
      RECT 77.165 2.725 77.18 2.998 ;
      RECT 77.16 2.725 77.165 3.043 ;
      RECT 77.155 2.725 77.16 3.073 ;
      RECT 77.15 2.725 77.155 3.093 ;
      RECT 77.14 2.725 77.15 3.128 ;
      RECT 77.125 2.725 77.14 3.16 ;
      RECT 77.08 2.725 77.125 3.188 ;
      RECT 77.075 2.725 77.08 3.218 ;
      RECT 77.07 2.725 77.075 3.23 ;
      RECT 77.065 2.725 77.07 3.238 ;
      RECT 77.055 2.725 77.065 3.253 ;
      RECT 77.05 2.725 77.055 3.275 ;
      RECT 77.04 2.725 77.05 3.298 ;
      RECT 77.035 2.725 77.04 3.318 ;
      RECT 77 2.74 77.02 3.335 ;
      RECT 76.975 2.757 77 3.335 ;
      RECT 76.97 2.767 76.975 3.335 ;
      RECT 76.94 2.782 76.97 3.335 ;
      RECT 76.865 2.824 76.94 3.335 ;
      RECT 76.86 2.855 76.865 3.318 ;
      RECT 76.855 2.859 76.86 3.3 ;
      RECT 76.85 2.863 76.855 3.263 ;
      RECT 76.845 3.047 76.85 3.23 ;
      RECT 76.33 3.236 76.416 3.801 ;
      RECT 76.285 3.238 76.45 3.795 ;
      RECT 76.416 3.235 76.45 3.795 ;
      RECT 76.33 3.237 76.535 3.789 ;
      RECT 76.285 3.247 76.545 3.785 ;
      RECT 76.26 3.239 76.535 3.781 ;
      RECT 76.255 3.242 76.535 3.776 ;
      RECT 76.23 3.257 76.545 3.77 ;
      RECT 76.23 3.282 76.585 3.765 ;
      RECT 76.19 3.29 76.585 3.74 ;
      RECT 76.19 3.317 76.6 3.738 ;
      RECT 76.19 3.347 76.61 3.725 ;
      RECT 76.185 3.492 76.61 3.713 ;
      RECT 76.19 3.421 76.63 3.71 ;
      RECT 76.19 3.478 76.635 3.518 ;
      RECT 76.38 2.757 76.55 2.935 ;
      RECT 76.33 2.696 76.38 2.92 ;
      RECT 76.065 2.676 76.33 2.905 ;
      RECT 76.025 2.74 76.5 2.905 ;
      RECT 76.025 2.73 76.455 2.905 ;
      RECT 76.025 2.727 76.445 2.905 ;
      RECT 76.025 2.715 76.435 2.905 ;
      RECT 76.025 2.7 76.38 2.905 ;
      RECT 76.065 2.672 76.266 2.905 ;
      RECT 76.075 2.65 76.266 2.905 ;
      RECT 76.1 2.635 76.18 2.905 ;
      RECT 75.855 3.165 75.975 3.61 ;
      RECT 75.84 3.165 75.975 3.609 ;
      RECT 75.795 3.187 75.975 3.604 ;
      RECT 75.755 3.236 75.975 3.598 ;
      RECT 75.755 3.236 75.98 3.573 ;
      RECT 75.755 3.236 76 3.463 ;
      RECT 75.75 3.266 76 3.46 ;
      RECT 75.84 3.165 76.01 3.355 ;
      RECT 75.5 1.95 75.505 2.395 ;
      RECT 75.31 1.95 75.33 2.36 ;
      RECT 75.28 1.95 75.285 2.335 ;
      RECT 75.96 2.257 75.975 2.445 ;
      RECT 75.955 2.242 75.96 2.451 ;
      RECT 75.935 2.215 75.955 2.454 ;
      RECT 75.885 2.182 75.935 2.463 ;
      RECT 75.855 2.162 75.885 2.467 ;
      RECT 75.836 2.15 75.855 2.463 ;
      RECT 75.75 2.122 75.836 2.453 ;
      RECT 75.74 2.097 75.75 2.443 ;
      RECT 75.67 2.065 75.74 2.435 ;
      RECT 75.645 2.025 75.67 2.427 ;
      RECT 75.625 2.007 75.645 2.421 ;
      RECT 75.615 1.997 75.625 2.418 ;
      RECT 75.605 1.99 75.615 2.416 ;
      RECT 75.585 1.977 75.605 2.413 ;
      RECT 75.575 1.967 75.585 2.41 ;
      RECT 75.565 1.96 75.575 2.408 ;
      RECT 75.515 1.952 75.565 2.402 ;
      RECT 75.505 1.95 75.515 2.396 ;
      RECT 75.475 1.95 75.5 2.393 ;
      RECT 75.446 1.95 75.475 2.388 ;
      RECT 75.36 1.95 75.446 2.378 ;
      RECT 75.33 1.95 75.36 2.365 ;
      RECT 75.285 1.95 75.31 2.348 ;
      RECT 75.27 1.95 75.28 2.33 ;
      RECT 75.25 1.957 75.27 2.315 ;
      RECT 75.245 1.972 75.25 2.303 ;
      RECT 75.24 1.977 75.245 2.243 ;
      RECT 75.235 1.982 75.24 2.085 ;
      RECT 75.23 1.985 75.235 2.003 ;
      RECT 75.495 2.67 75.581 2.991 ;
      RECT 75.495 2.67 75.615 2.984 ;
      RECT 75.445 2.67 75.615 2.98 ;
      RECT 75.445 2.672 75.701 2.978 ;
      RECT 75.445 2.674 75.725 2.972 ;
      RECT 75.445 2.681 75.735 2.971 ;
      RECT 75.445 2.69 75.74 2.968 ;
      RECT 75.445 2.696 75.745 2.963 ;
      RECT 75.445 2.74 75.75 2.96 ;
      RECT 75.445 2.832 75.755 2.957 ;
      RECT 74.97 3.275 75.005 3.595 ;
      RECT 75.555 3.46 75.56 3.642 ;
      RECT 75.51 3.342 75.555 3.661 ;
      RECT 75.495 3.319 75.51 3.684 ;
      RECT 75.485 3.309 75.495 3.694 ;
      RECT 75.465 3.304 75.485 3.707 ;
      RECT 75.44 3.302 75.465 3.728 ;
      RECT 75.421 3.301 75.44 3.74 ;
      RECT 75.335 3.298 75.421 3.74 ;
      RECT 75.265 3.293 75.335 3.728 ;
      RECT 75.19 3.289 75.265 3.703 ;
      RECT 75.125 3.285 75.19 3.67 ;
      RECT 75.055 3.282 75.125 3.63 ;
      RECT 75.025 3.278 75.055 3.605 ;
      RECT 75.005 3.276 75.025 3.598 ;
      RECT 74.921 3.274 74.97 3.596 ;
      RECT 74.835 3.271 74.921 3.597 ;
      RECT 74.76 3.27 74.835 3.599 ;
      RECT 74.675 3.27 74.76 3.625 ;
      RECT 74.598 3.271 74.675 3.65 ;
      RECT 74.512 3.272 74.598 3.65 ;
      RECT 74.426 3.272 74.512 3.65 ;
      RECT 74.34 3.273 74.426 3.65 ;
      RECT 74.32 3.274 74.34 3.642 ;
      RECT 74.305 3.28 74.32 3.627 ;
      RECT 74.27 3.3 74.305 3.607 ;
      RECT 74.26 3.32 74.27 3.589 ;
      RECT 75.23 2.625 75.235 2.895 ;
      RECT 75.225 2.616 75.23 2.9 ;
      RECT 75.215 2.606 75.225 2.912 ;
      RECT 75.21 2.595 75.215 2.923 ;
      RECT 75.19 2.589 75.21 2.941 ;
      RECT 75.145 2.586 75.19 2.99 ;
      RECT 75.13 2.585 75.145 3.035 ;
      RECT 75.125 2.585 75.13 3.048 ;
      RECT 75.115 2.585 75.125 3.06 ;
      RECT 75.11 2.586 75.115 3.075 ;
      RECT 75.09 2.594 75.11 3.08 ;
      RECT 75.06 2.61 75.09 3.08 ;
      RECT 75.05 2.622 75.055 3.08 ;
      RECT 75.015 2.637 75.05 3.08 ;
      RECT 74.985 2.657 75.015 3.08 ;
      RECT 74.975 2.682 74.985 3.08 ;
      RECT 74.97 2.71 74.975 3.08 ;
      RECT 74.965 2.74 74.97 3.08 ;
      RECT 74.96 2.757 74.965 3.08 ;
      RECT 74.95 2.785 74.96 3.08 ;
      RECT 74.94 2.82 74.95 3.08 ;
      RECT 74.935 2.855 74.94 3.08 ;
      RECT 75.055 2.62 75.06 3.08 ;
      RECT 74.57 2.722 74.755 2.895 ;
      RECT 74.53 2.64 74.715 2.893 ;
      RECT 74.491 2.645 74.715 2.889 ;
      RECT 74.405 2.654 74.715 2.884 ;
      RECT 74.321 2.67 74.72 2.879 ;
      RECT 74.235 2.69 74.745 2.873 ;
      RECT 74.235 2.71 74.75 2.873 ;
      RECT 74.321 2.68 74.745 2.879 ;
      RECT 74.405 2.655 74.72 2.884 ;
      RECT 74.57 2.637 74.715 2.895 ;
      RECT 74.57 2.632 74.67 2.895 ;
      RECT 74.656 2.626 74.67 2.895 ;
      RECT 74.045 1.95 74.05 2.349 ;
      RECT 73.79 1.95 73.825 2.347 ;
      RECT 73.385 1.985 73.39 2.341 ;
      RECT 74.13 1.988 74.135 2.243 ;
      RECT 74.125 1.986 74.13 2.249 ;
      RECT 74.12 1.985 74.125 2.256 ;
      RECT 74.095 1.978 74.12 2.28 ;
      RECT 74.09 1.971 74.095 2.304 ;
      RECT 74.085 1.967 74.09 2.313 ;
      RECT 74.075 1.962 74.085 2.326 ;
      RECT 74.07 1.959 74.075 2.335 ;
      RECT 74.065 1.957 74.07 2.34 ;
      RECT 74.05 1.953 74.065 2.35 ;
      RECT 74.035 1.947 74.045 2.349 ;
      RECT 73.997 1.945 74.035 2.349 ;
      RECT 73.911 1.947 73.997 2.349 ;
      RECT 73.825 1.949 73.911 2.348 ;
      RECT 73.754 1.95 73.79 2.347 ;
      RECT 73.668 1.952 73.754 2.347 ;
      RECT 73.582 1.954 73.668 2.346 ;
      RECT 73.496 1.956 73.582 2.346 ;
      RECT 73.41 1.959 73.496 2.345 ;
      RECT 73.4 1.965 73.41 2.344 ;
      RECT 73.39 1.977 73.4 2.342 ;
      RECT 73.33 2.012 73.385 2.338 ;
      RECT 73.325 2.042 73.33 2.1 ;
      RECT 74.07 3.122 74.085 3.315 ;
      RECT 74.065 3.09 74.07 3.315 ;
      RECT 74.055 3.065 74.065 3.315 ;
      RECT 74.05 3.037 74.055 3.315 ;
      RECT 74.02 2.96 74.05 3.315 ;
      RECT 73.995 2.842 74.02 3.315 ;
      RECT 73.99 2.78 73.995 3.315 ;
      RECT 73.98 2.767 73.99 3.315 ;
      RECT 73.96 2.757 73.98 3.315 ;
      RECT 73.945 2.74 73.96 3.315 ;
      RECT 73.915 2.728 73.945 3.315 ;
      RECT 73.91 2.727 73.915 3.26 ;
      RECT 73.905 2.727 73.91 3.218 ;
      RECT 73.89 2.726 73.905 3.17 ;
      RECT 73.875 2.726 73.89 3.108 ;
      RECT 73.855 2.726 73.875 3.068 ;
      RECT 73.85 2.726 73.855 3.053 ;
      RECT 73.825 2.725 73.85 3.048 ;
      RECT 73.755 2.724 73.825 3.035 ;
      RECT 73.74 2.723 73.755 3.02 ;
      RECT 73.71 2.722 73.74 3.003 ;
      RECT 73.705 2.722 73.71 2.988 ;
      RECT 73.655 2.721 73.705 2.968 ;
      RECT 73.59 2.72 73.655 2.923 ;
      RECT 73.585 2.72 73.59 2.895 ;
      RECT 73.67 3.257 73.675 3.514 ;
      RECT 73.65 3.176 73.67 3.531 ;
      RECT 73.63 3.17 73.65 3.56 ;
      RECT 73.57 3.157 73.63 3.58 ;
      RECT 73.525 3.141 73.57 3.581 ;
      RECT 73.441 3.129 73.525 3.569 ;
      RECT 73.355 3.116 73.441 3.553 ;
      RECT 73.345 3.109 73.355 3.545 ;
      RECT 73.3 3.106 73.345 3.485 ;
      RECT 73.28 3.102 73.3 3.4 ;
      RECT 73.265 3.1 73.28 3.353 ;
      RECT 73.235 3.097 73.265 3.323 ;
      RECT 73.2 3.093 73.235 3.3 ;
      RECT 73.157 3.088 73.2 3.288 ;
      RECT 73.071 3.079 73.157 3.297 ;
      RECT 72.985 3.068 73.071 3.309 ;
      RECT 72.92 3.059 72.985 3.318 ;
      RECT 72.9 3.05 72.92 3.323 ;
      RECT 72.895 3.043 72.9 3.325 ;
      RECT 72.855 3.028 72.895 3.322 ;
      RECT 72.835 3.007 72.855 3.317 ;
      RECT 72.82 2.995 72.835 3.31 ;
      RECT 72.815 2.987 72.82 3.303 ;
      RECT 72.8 2.967 72.815 3.296 ;
      RECT 72.795 2.83 72.8 3.29 ;
      RECT 72.715 2.719 72.795 3.262 ;
      RECT 72.706 2.712 72.715 3.228 ;
      RECT 72.62 2.706 72.706 3.153 ;
      RECT 72.595 2.697 72.62 3.065 ;
      RECT 72.565 2.692 72.595 3.04 ;
      RECT 72.5 2.701 72.565 3.025 ;
      RECT 72.48 2.717 72.5 3 ;
      RECT 72.47 2.723 72.48 2.948 ;
      RECT 72.45 2.745 72.47 2.83 ;
      RECT 73.105 2.71 73.275 2.895 ;
      RECT 73.105 2.71 73.31 2.893 ;
      RECT 73.155 2.62 73.325 2.884 ;
      RECT 73.105 2.777 73.33 2.877 ;
      RECT 73.12 2.655 73.325 2.884 ;
      RECT 72.32 3.388 72.385 3.831 ;
      RECT 72.26 3.413 72.385 3.829 ;
      RECT 72.26 3.413 72.44 3.823 ;
      RECT 72.245 3.438 72.44 3.822 ;
      RECT 72.385 3.375 72.46 3.819 ;
      RECT 72.32 3.4 72.54 3.813 ;
      RECT 72.245 3.439 72.585 3.807 ;
      RECT 72.23 3.466 72.585 3.798 ;
      RECT 72.245 3.459 72.605 3.79 ;
      RECT 72.23 3.468 72.61 3.773 ;
      RECT 72.225 3.485 72.61 3.6 ;
      RECT 72.23 2.207 72.265 2.445 ;
      RECT 72.23 2.207 72.295 2.444 ;
      RECT 72.23 2.207 72.41 2.44 ;
      RECT 72.23 2.207 72.465 2.418 ;
      RECT 72.24 2.15 72.52 2.318 ;
      RECT 72.345 1.99 72.375 2.441 ;
      RECT 72.375 1.985 72.555 2.198 ;
      RECT 72.245 2.126 72.555 2.198 ;
      RECT 72.295 2.022 72.345 2.442 ;
      RECT 72.265 2.078 72.555 2.198 ;
      RECT 70.775 1.74 70.945 2.935 ;
      RECT 70.775 1.74 71.24 1.91 ;
      RECT 70.775 6.97 71.24 7.14 ;
      RECT 70.775 5.945 70.945 7.14 ;
      RECT 69.785 1.74 69.955 2.935 ;
      RECT 69.785 1.74 70.25 1.91 ;
      RECT 69.785 6.97 70.25 7.14 ;
      RECT 69.785 5.945 69.955 7.14 ;
      RECT 67.93 2.635 68.1 3.865 ;
      RECT 67.985 0.855 68.155 2.805 ;
      RECT 67.93 0.575 68.1 1.025 ;
      RECT 67.93 7.855 68.1 8.305 ;
      RECT 67.985 6.075 68.155 8.025 ;
      RECT 67.93 5.015 68.1 6.245 ;
      RECT 67.41 0.575 67.58 3.865 ;
      RECT 67.41 2.075 67.815 2.405 ;
      RECT 67.41 1.235 67.815 1.565 ;
      RECT 67.41 5.015 67.58 8.305 ;
      RECT 67.41 7.315 67.815 7.645 ;
      RECT 67.41 6.475 67.815 6.805 ;
      RECT 65.51 3.392 65.525 3.443 ;
      RECT 65.505 3.372 65.51 3.49 ;
      RECT 65.49 3.362 65.505 3.558 ;
      RECT 65.465 3.342 65.49 3.613 ;
      RECT 65.425 3.327 65.465 3.633 ;
      RECT 65.38 3.321 65.425 3.661 ;
      RECT 65.31 3.311 65.38 3.678 ;
      RECT 65.29 3.303 65.31 3.678 ;
      RECT 65.23 3.297 65.29 3.67 ;
      RECT 65.171 3.288 65.23 3.658 ;
      RECT 65.085 3.277 65.171 3.641 ;
      RECT 65.063 3.268 65.085 3.629 ;
      RECT 64.977 3.261 65.063 3.616 ;
      RECT 64.891 3.248 64.977 3.597 ;
      RECT 64.805 3.236 64.891 3.577 ;
      RECT 64.775 3.225 64.805 3.564 ;
      RECT 64.725 3.211 64.775 3.556 ;
      RECT 64.705 3.2 64.725 3.548 ;
      RECT 64.656 3.189 64.705 3.54 ;
      RECT 64.57 3.168 64.656 3.525 ;
      RECT 64.525 3.155 64.57 3.51 ;
      RECT 64.48 3.155 64.525 3.49 ;
      RECT 64.425 3.155 64.48 3.425 ;
      RECT 64.4 3.155 64.425 3.348 ;
      RECT 64.925 2.892 65.095 3.075 ;
      RECT 64.925 2.892 65.11 3.033 ;
      RECT 64.925 2.892 65.115 2.975 ;
      RECT 64.985 2.66 65.12 2.951 ;
      RECT 64.985 2.664 65.125 2.934 ;
      RECT 64.93 2.827 65.125 2.934 ;
      RECT 64.955 2.672 65.095 3.075 ;
      RECT 64.955 2.676 65.135 2.875 ;
      RECT 64.94 2.762 65.135 2.875 ;
      RECT 64.95 2.692 65.095 3.075 ;
      RECT 64.95 2.695 65.145 2.788 ;
      RECT 64.945 2.712 65.145 2.788 ;
      RECT 64.715 1.932 64.885 2.415 ;
      RECT 64.71 1.927 64.86 2.405 ;
      RECT 64.71 1.934 64.89 2.399 ;
      RECT 64.7 1.928 64.86 2.378 ;
      RECT 64.7 1.944 64.905 2.337 ;
      RECT 64.67 1.929 64.86 2.3 ;
      RECT 64.67 1.959 64.915 2.24 ;
      RECT 64.665 1.931 64.86 2.238 ;
      RECT 64.645 1.94 64.89 2.195 ;
      RECT 64.62 1.956 64.905 2.107 ;
      RECT 64.62 1.975 64.93 2.098 ;
      RECT 64.615 2.012 64.93 2.05 ;
      RECT 64.62 1.992 64.935 2.018 ;
      RECT 64.715 1.926 64.825 2.415 ;
      RECT 64.801 1.925 64.825 2.415 ;
      RECT 64.035 2.71 64.04 2.921 ;
      RECT 64.635 2.71 64.64 2.895 ;
      RECT 64.7 2.75 64.705 2.863 ;
      RECT 64.695 2.742 64.7 2.869 ;
      RECT 64.69 2.732 64.695 2.877 ;
      RECT 64.685 2.722 64.69 2.886 ;
      RECT 64.68 2.712 64.685 2.89 ;
      RECT 64.64 2.71 64.68 2.893 ;
      RECT 64.612 2.709 64.635 2.897 ;
      RECT 64.526 2.706 64.612 2.904 ;
      RECT 64.44 2.702 64.526 2.915 ;
      RECT 64.42 2.7 64.44 2.921 ;
      RECT 64.402 2.699 64.42 2.924 ;
      RECT 64.316 2.697 64.402 2.931 ;
      RECT 64.23 2.692 64.316 2.944 ;
      RECT 64.211 2.689 64.23 2.949 ;
      RECT 64.125 2.687 64.211 2.94 ;
      RECT 64.115 2.687 64.125 2.933 ;
      RECT 64.04 2.7 64.115 2.927 ;
      RECT 64.025 2.711 64.035 2.921 ;
      RECT 64.015 2.713 64.025 2.92 ;
      RECT 64.005 2.717 64.015 2.916 ;
      RECT 64 2.72 64.005 2.91 ;
      RECT 63.99 2.722 64 2.904 ;
      RECT 63.985 2.725 63.99 2.898 ;
      RECT 63.965 3.311 63.97 3.515 ;
      RECT 63.95 3.298 63.965 3.608 ;
      RECT 63.935 3.279 63.95 3.885 ;
      RECT 63.9 3.245 63.935 3.885 ;
      RECT 63.896 3.215 63.9 3.885 ;
      RECT 63.81 3.097 63.896 3.885 ;
      RECT 63.8 2.972 63.81 3.885 ;
      RECT 63.785 2.94 63.8 3.885 ;
      RECT 63.78 2.915 63.785 3.885 ;
      RECT 63.775 2.905 63.78 3.841 ;
      RECT 63.76 2.877 63.775 3.746 ;
      RECT 63.745 2.843 63.76 3.645 ;
      RECT 63.74 2.821 63.745 3.598 ;
      RECT 63.735 2.81 63.74 3.568 ;
      RECT 63.73 2.8 63.735 3.534 ;
      RECT 63.72 2.787 63.73 3.502 ;
      RECT 63.695 2.763 63.72 3.428 ;
      RECT 63.69 2.743 63.695 3.353 ;
      RECT 63.685 2.737 63.69 3.328 ;
      RECT 63.68 2.732 63.685 3.293 ;
      RECT 63.675 2.727 63.68 3.268 ;
      RECT 63.67 2.725 63.675 3.248 ;
      RECT 63.665 2.725 63.67 3.233 ;
      RECT 63.66 2.725 63.665 3.193 ;
      RECT 63.65 2.725 63.66 3.165 ;
      RECT 63.64 2.725 63.65 3.11 ;
      RECT 63.625 2.725 63.64 3.048 ;
      RECT 63.62 2.724 63.625 2.993 ;
      RECT 63.605 2.723 63.62 2.973 ;
      RECT 63.545 2.721 63.605 2.947 ;
      RECT 63.51 2.722 63.545 2.927 ;
      RECT 63.505 2.724 63.51 2.917 ;
      RECT 63.495 2.743 63.505 2.907 ;
      RECT 63.49 2.77 63.495 2.838 ;
      RECT 63.605 2.195 63.775 2.44 ;
      RECT 63.64 1.966 63.775 2.44 ;
      RECT 63.64 1.968 63.785 2.435 ;
      RECT 63.64 1.97 63.81 2.423 ;
      RECT 63.64 1.973 63.835 2.405 ;
      RECT 63.64 1.978 63.885 2.378 ;
      RECT 63.64 1.983 63.905 2.343 ;
      RECT 63.62 1.985 63.915 2.318 ;
      RECT 63.61 2.08 63.915 2.318 ;
      RECT 63.64 1.965 63.75 2.44 ;
      RECT 63.65 1.962 63.745 2.44 ;
      RECT 63.17 3.227 63.36 3.585 ;
      RECT 63.17 3.239 63.395 3.584 ;
      RECT 63.17 3.267 63.415 3.582 ;
      RECT 63.17 3.292 63.42 3.581 ;
      RECT 63.17 3.35 63.435 3.58 ;
      RECT 63.155 3.223 63.315 3.565 ;
      RECT 63.135 3.232 63.36 3.518 ;
      RECT 63.11 3.243 63.395 3.455 ;
      RECT 63.11 3.327 63.43 3.455 ;
      RECT 63.11 3.302 63.425 3.455 ;
      RECT 63.17 3.218 63.315 3.585 ;
      RECT 63.256 3.217 63.315 3.585 ;
      RECT 63.256 3.216 63.3 3.585 ;
      RECT 62.955 2.732 62.96 3.11 ;
      RECT 62.95 2.7 62.955 3.11 ;
      RECT 62.945 2.672 62.95 3.11 ;
      RECT 62.94 2.652 62.945 3.11 ;
      RECT 62.885 2.635 62.94 3.11 ;
      RECT 62.845 2.62 62.885 3.11 ;
      RECT 62.79 2.607 62.845 3.11 ;
      RECT 62.755 2.598 62.79 3.11 ;
      RECT 62.751 2.596 62.755 3.109 ;
      RECT 62.665 2.592 62.751 3.092 ;
      RECT 62.58 2.584 62.665 3.055 ;
      RECT 62.57 2.58 62.58 3.028 ;
      RECT 62.56 2.58 62.57 3.01 ;
      RECT 62.55 2.582 62.56 2.993 ;
      RECT 62.545 2.587 62.55 2.979 ;
      RECT 62.54 2.591 62.545 2.966 ;
      RECT 62.53 2.596 62.54 2.95 ;
      RECT 62.515 2.61 62.53 2.925 ;
      RECT 62.51 2.616 62.515 2.905 ;
      RECT 62.505 2.618 62.51 2.898 ;
      RECT 62.5 2.622 62.505 2.773 ;
      RECT 62.68 3.422 62.925 3.885 ;
      RECT 62.6 3.395 62.92 3.881 ;
      RECT 62.53 3.43 62.925 3.874 ;
      RECT 62.32 3.685 62.925 3.87 ;
      RECT 62.5 3.453 62.925 3.87 ;
      RECT 62.34 3.645 62.925 3.87 ;
      RECT 62.49 3.465 62.925 3.87 ;
      RECT 62.375 3.582 62.925 3.87 ;
      RECT 62.43 3.507 62.925 3.87 ;
      RECT 62.68 3.372 62.92 3.885 ;
      RECT 62.71 3.365 62.92 3.885 ;
      RECT 62.7 3.367 62.92 3.885 ;
      RECT 62.71 3.362 62.84 3.885 ;
      RECT 62.265 1.925 62.351 2.364 ;
      RECT 62.26 1.925 62.351 2.362 ;
      RECT 62.26 1.925 62.42 2.361 ;
      RECT 62.26 1.925 62.45 2.358 ;
      RECT 62.245 1.932 62.45 2.349 ;
      RECT 62.245 1.932 62.455 2.345 ;
      RECT 62.24 1.942 62.455 2.338 ;
      RECT 62.235 1.947 62.455 2.313 ;
      RECT 62.235 1.947 62.47 2.295 ;
      RECT 62.26 1.925 62.49 2.21 ;
      RECT 62.23 1.952 62.49 2.208 ;
      RECT 62.24 1.945 62.495 2.146 ;
      RECT 62.23 2.067 62.5 2.129 ;
      RECT 62.215 1.962 62.495 2.08 ;
      RECT 62.21 1.972 62.495 1.98 ;
      RECT 62.29 2.743 62.295 2.82 ;
      RECT 62.28 2.737 62.29 3.01 ;
      RECT 62.27 2.729 62.28 3.031 ;
      RECT 62.26 2.72 62.27 3.053 ;
      RECT 62.255 2.715 62.26 3.07 ;
      RECT 62.215 2.715 62.255 3.11 ;
      RECT 62.195 2.715 62.215 3.165 ;
      RECT 62.19 2.715 62.195 3.193 ;
      RECT 62.18 2.715 62.19 3.208 ;
      RECT 62.145 2.715 62.18 3.25 ;
      RECT 62.14 2.715 62.145 3.293 ;
      RECT 62.13 2.715 62.14 3.308 ;
      RECT 62.115 2.715 62.13 3.328 ;
      RECT 62.1 2.715 62.115 3.355 ;
      RECT 62.095 2.716 62.1 3.373 ;
      RECT 62.075 2.717 62.095 3.38 ;
      RECT 62.02 2.718 62.075 3.4 ;
      RECT 62.01 2.719 62.02 3.414 ;
      RECT 62.005 2.722 62.01 3.413 ;
      RECT 61.965 2.795 62.005 3.411 ;
      RECT 61.95 2.875 61.965 3.409 ;
      RECT 61.925 2.93 61.95 3.407 ;
      RECT 61.91 2.995 61.925 3.406 ;
      RECT 61.865 3.027 61.91 3.403 ;
      RECT 61.78 3.05 61.865 3.398 ;
      RECT 61.755 3.07 61.78 3.393 ;
      RECT 61.685 3.075 61.755 3.389 ;
      RECT 61.665 3.077 61.685 3.386 ;
      RECT 61.58 3.088 61.665 3.38 ;
      RECT 61.575 3.099 61.58 3.375 ;
      RECT 61.565 3.101 61.575 3.375 ;
      RECT 61.53 3.105 61.565 3.373 ;
      RECT 61.48 3.115 61.53 3.36 ;
      RECT 61.46 3.123 61.48 3.345 ;
      RECT 61.38 3.135 61.46 3.328 ;
      RECT 61.545 2.685 61.715 2.895 ;
      RECT 61.661 2.681 61.715 2.895 ;
      RECT 61.466 2.685 61.715 2.886 ;
      RECT 61.466 2.685 61.72 2.875 ;
      RECT 61.38 2.685 61.72 2.866 ;
      RECT 61.38 2.693 61.73 2.81 ;
      RECT 61.38 2.705 61.735 2.723 ;
      RECT 61.38 2.712 61.74 2.715 ;
      RECT 61.575 2.683 61.715 2.895 ;
      RECT 61.33 3.628 61.575 3.96 ;
      RECT 61.325 3.62 61.33 3.957 ;
      RECT 61.295 3.64 61.575 3.938 ;
      RECT 61.275 3.672 61.575 3.911 ;
      RECT 61.325 3.625 61.502 3.957 ;
      RECT 61.325 3.622 61.416 3.957 ;
      RECT 61.265 1.97 61.435 2.39 ;
      RECT 61.26 1.97 61.435 2.388 ;
      RECT 61.26 1.97 61.46 2.378 ;
      RECT 61.26 1.97 61.48 2.353 ;
      RECT 61.255 1.97 61.48 2.348 ;
      RECT 61.255 1.97 61.49 2.338 ;
      RECT 61.255 1.97 61.495 2.333 ;
      RECT 61.255 1.975 61.5 2.328 ;
      RECT 61.255 2.007 61.515 2.318 ;
      RECT 61.255 2.077 61.54 2.301 ;
      RECT 61.235 2.077 61.54 2.293 ;
      RECT 61.235 2.137 61.55 2.27 ;
      RECT 61.235 2.177 61.56 2.215 ;
      RECT 61.22 1.97 61.495 2.195 ;
      RECT 61.21 1.985 61.5 2.093 ;
      RECT 60.8 3.375 60.97 3.9 ;
      RECT 60.795 3.375 60.97 3.893 ;
      RECT 60.785 3.375 60.975 3.858 ;
      RECT 60.78 3.385 60.975 3.83 ;
      RECT 60.775 3.405 60.975 3.813 ;
      RECT 60.785 3.38 60.98 3.803 ;
      RECT 60.77 3.425 60.98 3.795 ;
      RECT 60.765 3.445 60.98 3.78 ;
      RECT 60.76 3.475 60.98 3.77 ;
      RECT 60.75 3.52 60.98 3.745 ;
      RECT 60.78 3.39 60.985 3.728 ;
      RECT 60.745 3.572 60.985 3.723 ;
      RECT 60.78 3.4 60.99 3.693 ;
      RECT 60.74 3.605 60.99 3.69 ;
      RECT 60.735 3.63 60.99 3.67 ;
      RECT 60.775 3.417 61 3.61 ;
      RECT 60.77 3.439 61.01 3.503 ;
      RECT 60.72 2.686 60.735 2.955 ;
      RECT 60.675 2.67 60.72 3 ;
      RECT 60.67 2.658 60.675 3.05 ;
      RECT 60.66 2.654 60.67 3.083 ;
      RECT 60.655 2.651 60.66 3.111 ;
      RECT 60.64 2.653 60.655 3.153 ;
      RECT 60.635 2.657 60.64 3.193 ;
      RECT 60.615 2.662 60.635 3.245 ;
      RECT 60.611 2.667 60.615 3.302 ;
      RECT 60.525 2.686 60.611 3.339 ;
      RECT 60.515 2.707 60.525 3.375 ;
      RECT 60.51 2.715 60.515 3.376 ;
      RECT 60.505 2.757 60.51 3.377 ;
      RECT 60.49 2.845 60.505 3.378 ;
      RECT 60.48 2.995 60.49 3.38 ;
      RECT 60.475 3.04 60.48 3.382 ;
      RECT 60.44 3.082 60.475 3.385 ;
      RECT 60.435 3.1 60.44 3.388 ;
      RECT 60.358 3.106 60.435 3.394 ;
      RECT 60.272 3.12 60.358 3.407 ;
      RECT 60.186 3.134 60.272 3.421 ;
      RECT 60.1 3.148 60.186 3.434 ;
      RECT 60.04 3.16 60.1 3.446 ;
      RECT 60.015 3.167 60.04 3.453 ;
      RECT 60.001 3.17 60.015 3.458 ;
      RECT 59.915 3.178 60.001 3.474 ;
      RECT 59.91 3.185 59.915 3.489 ;
      RECT 59.886 3.185 59.91 3.496 ;
      RECT 59.8 3.188 59.886 3.524 ;
      RECT 59.715 3.192 59.8 3.568 ;
      RECT 59.65 3.196 59.715 3.605 ;
      RECT 59.625 3.199 59.65 3.621 ;
      RECT 59.55 3.212 59.625 3.625 ;
      RECT 59.525 3.23 59.55 3.629 ;
      RECT 59.515 3.237 59.525 3.631 ;
      RECT 59.5 3.24 59.515 3.632 ;
      RECT 59.44 3.252 59.5 3.636 ;
      RECT 59.43 3.266 59.44 3.64 ;
      RECT 59.375 3.276 59.43 3.628 ;
      RECT 59.35 3.297 59.375 3.611 ;
      RECT 59.33 3.317 59.35 3.602 ;
      RECT 59.325 3.33 59.33 3.597 ;
      RECT 59.31 3.342 59.325 3.593 ;
      RECT 60.545 1.997 60.55 2.02 ;
      RECT 60.54 1.988 60.545 2.06 ;
      RECT 60.535 1.986 60.54 2.103 ;
      RECT 60.53 1.977 60.535 2.138 ;
      RECT 60.525 1.967 60.53 2.21 ;
      RECT 60.52 1.957 60.525 2.275 ;
      RECT 60.515 1.954 60.52 2.315 ;
      RECT 60.49 1.948 60.515 2.405 ;
      RECT 60.455 1.936 60.49 2.43 ;
      RECT 60.445 1.927 60.455 2.43 ;
      RECT 60.31 1.925 60.32 2.413 ;
      RECT 60.3 1.925 60.31 2.38 ;
      RECT 60.295 1.925 60.3 2.355 ;
      RECT 60.29 1.925 60.295 2.343 ;
      RECT 60.285 1.925 60.29 2.325 ;
      RECT 60.275 1.925 60.285 2.29 ;
      RECT 60.27 1.927 60.275 2.268 ;
      RECT 60.265 1.933 60.27 2.253 ;
      RECT 60.26 1.939 60.265 2.238 ;
      RECT 60.245 1.951 60.26 2.211 ;
      RECT 60.24 1.962 60.245 2.179 ;
      RECT 60.235 1.972 60.24 2.163 ;
      RECT 60.225 1.98 60.235 2.132 ;
      RECT 60.22 1.99 60.225 2.106 ;
      RECT 60.215 2.047 60.22 2.089 ;
      RECT 60.32 1.925 60.445 2.43 ;
      RECT 60.035 2.612 60.295 2.91 ;
      RECT 60.03 2.619 60.295 2.908 ;
      RECT 60.035 2.614 60.31 2.903 ;
      RECT 60.025 2.627 60.31 2.9 ;
      RECT 60.025 2.632 60.315 2.893 ;
      RECT 60.02 2.64 60.315 2.89 ;
      RECT 60.02 2.657 60.32 2.688 ;
      RECT 60.035 2.609 60.266 2.91 ;
      RECT 60.09 2.608 60.266 2.91 ;
      RECT 60.09 2.605 60.18 2.91 ;
      RECT 60.09 2.602 60.176 2.91 ;
      RECT 59.78 2.875 59.785 2.888 ;
      RECT 59.775 2.842 59.78 2.893 ;
      RECT 59.77 2.797 59.775 2.9 ;
      RECT 59.765 2.752 59.77 2.908 ;
      RECT 59.76 2.72 59.765 2.916 ;
      RECT 59.755 2.68 59.76 2.917 ;
      RECT 59.74 2.66 59.755 2.919 ;
      RECT 59.665 2.642 59.74 2.931 ;
      RECT 59.655 2.635 59.665 2.942 ;
      RECT 59.65 2.635 59.655 2.944 ;
      RECT 59.62 2.641 59.65 2.948 ;
      RECT 59.58 2.654 59.62 2.948 ;
      RECT 59.555 2.665 59.58 2.934 ;
      RECT 59.54 2.671 59.555 2.917 ;
      RECT 59.53 2.673 59.54 2.908 ;
      RECT 59.525 2.674 59.53 2.903 ;
      RECT 59.52 2.675 59.525 2.898 ;
      RECT 59.515 2.676 59.52 2.895 ;
      RECT 59.49 2.681 59.515 2.885 ;
      RECT 59.48 2.697 59.49 2.872 ;
      RECT 59.475 2.717 59.48 2.867 ;
      RECT 59.485 2.11 59.49 2.306 ;
      RECT 59.47 2.074 59.485 2.308 ;
      RECT 59.46 2.056 59.47 2.313 ;
      RECT 59.45 2.042 59.46 2.317 ;
      RECT 59.405 2.026 59.45 2.327 ;
      RECT 59.4 2.016 59.405 2.336 ;
      RECT 59.355 2.005 59.4 2.342 ;
      RECT 59.35 1.993 59.355 2.349 ;
      RECT 59.335 1.988 59.35 2.353 ;
      RECT 59.32 1.98 59.335 2.358 ;
      RECT 59.31 1.973 59.32 2.363 ;
      RECT 59.3 1.97 59.31 2.368 ;
      RECT 59.29 1.97 59.3 2.369 ;
      RECT 59.285 1.967 59.29 2.368 ;
      RECT 59.25 1.962 59.275 2.367 ;
      RECT 59.226 1.958 59.25 2.366 ;
      RECT 59.14 1.949 59.226 2.363 ;
      RECT 59.125 1.941 59.14 2.36 ;
      RECT 59.103 1.94 59.125 2.359 ;
      RECT 59.017 1.94 59.103 2.357 ;
      RECT 58.931 1.94 59.017 2.355 ;
      RECT 58.845 1.94 58.931 2.352 ;
      RECT 58.835 1.94 58.845 2.343 ;
      RECT 58.805 1.94 58.835 2.303 ;
      RECT 58.795 1.95 58.805 2.258 ;
      RECT 58.79 1.99 58.795 2.243 ;
      RECT 58.785 2.005 58.79 2.23 ;
      RECT 58.755 2.085 58.785 2.192 ;
      RECT 59.275 1.965 59.285 2.368 ;
      RECT 59.1 2.73 59.115 3.335 ;
      RECT 59.105 2.725 59.115 3.335 ;
      RECT 59.27 2.725 59.275 2.908 ;
      RECT 59.26 2.725 59.27 2.938 ;
      RECT 59.245 2.725 59.26 2.998 ;
      RECT 59.24 2.725 59.245 3.043 ;
      RECT 59.235 2.725 59.24 3.073 ;
      RECT 59.23 2.725 59.235 3.093 ;
      RECT 59.22 2.725 59.23 3.128 ;
      RECT 59.205 2.725 59.22 3.16 ;
      RECT 59.16 2.725 59.205 3.188 ;
      RECT 59.155 2.725 59.16 3.218 ;
      RECT 59.15 2.725 59.155 3.23 ;
      RECT 59.145 2.725 59.15 3.238 ;
      RECT 59.135 2.725 59.145 3.253 ;
      RECT 59.13 2.725 59.135 3.275 ;
      RECT 59.12 2.725 59.13 3.298 ;
      RECT 59.115 2.725 59.12 3.318 ;
      RECT 59.08 2.74 59.1 3.335 ;
      RECT 59.055 2.757 59.08 3.335 ;
      RECT 59.05 2.767 59.055 3.335 ;
      RECT 59.02 2.782 59.05 3.335 ;
      RECT 58.945 2.824 59.02 3.335 ;
      RECT 58.94 2.855 58.945 3.318 ;
      RECT 58.935 2.859 58.94 3.3 ;
      RECT 58.93 2.863 58.935 3.263 ;
      RECT 58.925 3.047 58.93 3.23 ;
      RECT 58.41 3.236 58.496 3.801 ;
      RECT 58.365 3.238 58.53 3.795 ;
      RECT 58.496 3.235 58.53 3.795 ;
      RECT 58.41 3.237 58.615 3.789 ;
      RECT 58.365 3.247 58.625 3.785 ;
      RECT 58.34 3.239 58.615 3.781 ;
      RECT 58.335 3.242 58.615 3.776 ;
      RECT 58.31 3.257 58.625 3.77 ;
      RECT 58.31 3.282 58.665 3.765 ;
      RECT 58.27 3.29 58.665 3.74 ;
      RECT 58.27 3.317 58.68 3.738 ;
      RECT 58.27 3.347 58.69 3.725 ;
      RECT 58.265 3.492 58.69 3.713 ;
      RECT 58.27 3.421 58.71 3.71 ;
      RECT 58.27 3.478 58.715 3.518 ;
      RECT 58.46 2.757 58.63 2.935 ;
      RECT 58.41 2.696 58.46 2.92 ;
      RECT 58.145 2.676 58.41 2.905 ;
      RECT 58.105 2.74 58.58 2.905 ;
      RECT 58.105 2.73 58.535 2.905 ;
      RECT 58.105 2.727 58.525 2.905 ;
      RECT 58.105 2.715 58.515 2.905 ;
      RECT 58.105 2.7 58.46 2.905 ;
      RECT 58.145 2.672 58.346 2.905 ;
      RECT 58.155 2.65 58.346 2.905 ;
      RECT 58.18 2.635 58.26 2.905 ;
      RECT 57.935 3.165 58.055 3.61 ;
      RECT 57.92 3.165 58.055 3.609 ;
      RECT 57.875 3.187 58.055 3.604 ;
      RECT 57.835 3.236 58.055 3.598 ;
      RECT 57.835 3.236 58.06 3.573 ;
      RECT 57.835 3.236 58.08 3.463 ;
      RECT 57.83 3.266 58.08 3.46 ;
      RECT 57.92 3.165 58.09 3.355 ;
      RECT 57.58 1.95 57.585 2.395 ;
      RECT 57.39 1.95 57.41 2.36 ;
      RECT 57.36 1.95 57.365 2.335 ;
      RECT 58.04 2.257 58.055 2.445 ;
      RECT 58.035 2.242 58.04 2.451 ;
      RECT 58.015 2.215 58.035 2.454 ;
      RECT 57.965 2.182 58.015 2.463 ;
      RECT 57.935 2.162 57.965 2.467 ;
      RECT 57.916 2.15 57.935 2.463 ;
      RECT 57.83 2.122 57.916 2.453 ;
      RECT 57.82 2.097 57.83 2.443 ;
      RECT 57.75 2.065 57.82 2.435 ;
      RECT 57.725 2.025 57.75 2.427 ;
      RECT 57.705 2.007 57.725 2.421 ;
      RECT 57.695 1.997 57.705 2.418 ;
      RECT 57.685 1.99 57.695 2.416 ;
      RECT 57.665 1.977 57.685 2.413 ;
      RECT 57.655 1.967 57.665 2.41 ;
      RECT 57.645 1.96 57.655 2.408 ;
      RECT 57.595 1.952 57.645 2.402 ;
      RECT 57.585 1.95 57.595 2.396 ;
      RECT 57.555 1.95 57.58 2.393 ;
      RECT 57.526 1.95 57.555 2.388 ;
      RECT 57.44 1.95 57.526 2.378 ;
      RECT 57.41 1.95 57.44 2.365 ;
      RECT 57.365 1.95 57.39 2.348 ;
      RECT 57.35 1.95 57.36 2.33 ;
      RECT 57.33 1.957 57.35 2.315 ;
      RECT 57.325 1.972 57.33 2.303 ;
      RECT 57.32 1.977 57.325 2.243 ;
      RECT 57.315 1.982 57.32 2.085 ;
      RECT 57.31 1.985 57.315 2.003 ;
      RECT 57.575 2.67 57.661 2.991 ;
      RECT 57.575 2.67 57.695 2.984 ;
      RECT 57.525 2.67 57.695 2.98 ;
      RECT 57.525 2.672 57.781 2.978 ;
      RECT 57.525 2.674 57.805 2.972 ;
      RECT 57.525 2.681 57.815 2.971 ;
      RECT 57.525 2.69 57.82 2.968 ;
      RECT 57.525 2.696 57.825 2.963 ;
      RECT 57.525 2.74 57.83 2.96 ;
      RECT 57.525 2.832 57.835 2.957 ;
      RECT 57.05 3.275 57.085 3.595 ;
      RECT 57.635 3.46 57.64 3.642 ;
      RECT 57.59 3.342 57.635 3.661 ;
      RECT 57.575 3.319 57.59 3.684 ;
      RECT 57.565 3.309 57.575 3.694 ;
      RECT 57.545 3.304 57.565 3.707 ;
      RECT 57.52 3.302 57.545 3.728 ;
      RECT 57.501 3.301 57.52 3.74 ;
      RECT 57.415 3.298 57.501 3.74 ;
      RECT 57.345 3.293 57.415 3.728 ;
      RECT 57.27 3.289 57.345 3.703 ;
      RECT 57.205 3.285 57.27 3.67 ;
      RECT 57.135 3.282 57.205 3.63 ;
      RECT 57.105 3.278 57.135 3.605 ;
      RECT 57.085 3.276 57.105 3.598 ;
      RECT 57.001 3.274 57.05 3.596 ;
      RECT 56.915 3.271 57.001 3.597 ;
      RECT 56.84 3.27 56.915 3.599 ;
      RECT 56.755 3.27 56.84 3.625 ;
      RECT 56.678 3.271 56.755 3.65 ;
      RECT 56.592 3.272 56.678 3.65 ;
      RECT 56.506 3.272 56.592 3.65 ;
      RECT 56.42 3.273 56.506 3.65 ;
      RECT 56.4 3.274 56.42 3.642 ;
      RECT 56.385 3.28 56.4 3.627 ;
      RECT 56.35 3.3 56.385 3.607 ;
      RECT 56.34 3.32 56.35 3.589 ;
      RECT 57.31 2.625 57.315 2.895 ;
      RECT 57.305 2.616 57.31 2.9 ;
      RECT 57.295 2.606 57.305 2.912 ;
      RECT 57.29 2.595 57.295 2.923 ;
      RECT 57.27 2.589 57.29 2.941 ;
      RECT 57.225 2.586 57.27 2.99 ;
      RECT 57.21 2.585 57.225 3.035 ;
      RECT 57.205 2.585 57.21 3.048 ;
      RECT 57.195 2.585 57.205 3.06 ;
      RECT 57.19 2.586 57.195 3.075 ;
      RECT 57.17 2.594 57.19 3.08 ;
      RECT 57.14 2.61 57.17 3.08 ;
      RECT 57.13 2.622 57.135 3.08 ;
      RECT 57.095 2.637 57.13 3.08 ;
      RECT 57.065 2.657 57.095 3.08 ;
      RECT 57.055 2.682 57.065 3.08 ;
      RECT 57.05 2.71 57.055 3.08 ;
      RECT 57.045 2.74 57.05 3.08 ;
      RECT 57.04 2.757 57.045 3.08 ;
      RECT 57.03 2.785 57.04 3.08 ;
      RECT 57.02 2.82 57.03 3.08 ;
      RECT 57.015 2.855 57.02 3.08 ;
      RECT 57.135 2.62 57.14 3.08 ;
      RECT 56.65 2.722 56.835 2.895 ;
      RECT 56.61 2.64 56.795 2.893 ;
      RECT 56.571 2.645 56.795 2.889 ;
      RECT 56.485 2.654 56.795 2.884 ;
      RECT 56.401 2.67 56.8 2.879 ;
      RECT 56.315 2.69 56.825 2.873 ;
      RECT 56.315 2.71 56.83 2.873 ;
      RECT 56.401 2.68 56.825 2.879 ;
      RECT 56.485 2.655 56.8 2.884 ;
      RECT 56.65 2.637 56.795 2.895 ;
      RECT 56.65 2.632 56.75 2.895 ;
      RECT 56.736 2.626 56.75 2.895 ;
      RECT 56.125 1.95 56.13 2.349 ;
      RECT 55.87 1.95 55.905 2.347 ;
      RECT 55.465 1.985 55.47 2.341 ;
      RECT 56.21 1.988 56.215 2.243 ;
      RECT 56.205 1.986 56.21 2.249 ;
      RECT 56.2 1.985 56.205 2.256 ;
      RECT 56.175 1.978 56.2 2.28 ;
      RECT 56.17 1.971 56.175 2.304 ;
      RECT 56.165 1.967 56.17 2.313 ;
      RECT 56.155 1.962 56.165 2.326 ;
      RECT 56.15 1.959 56.155 2.335 ;
      RECT 56.145 1.957 56.15 2.34 ;
      RECT 56.13 1.953 56.145 2.35 ;
      RECT 56.115 1.947 56.125 2.349 ;
      RECT 56.077 1.945 56.115 2.349 ;
      RECT 55.991 1.947 56.077 2.349 ;
      RECT 55.905 1.949 55.991 2.348 ;
      RECT 55.834 1.95 55.87 2.347 ;
      RECT 55.748 1.952 55.834 2.347 ;
      RECT 55.662 1.954 55.748 2.346 ;
      RECT 55.576 1.956 55.662 2.346 ;
      RECT 55.49 1.959 55.576 2.345 ;
      RECT 55.48 1.965 55.49 2.344 ;
      RECT 55.47 1.977 55.48 2.342 ;
      RECT 55.41 2.012 55.465 2.338 ;
      RECT 55.405 2.042 55.41 2.1 ;
      RECT 56.15 3.122 56.165 3.315 ;
      RECT 56.145 3.09 56.15 3.315 ;
      RECT 56.135 3.065 56.145 3.315 ;
      RECT 56.13 3.037 56.135 3.315 ;
      RECT 56.1 2.96 56.13 3.315 ;
      RECT 56.075 2.842 56.1 3.315 ;
      RECT 56.07 2.78 56.075 3.315 ;
      RECT 56.06 2.767 56.07 3.315 ;
      RECT 56.04 2.757 56.06 3.315 ;
      RECT 56.025 2.74 56.04 3.315 ;
      RECT 55.995 2.728 56.025 3.315 ;
      RECT 55.99 2.727 55.995 3.26 ;
      RECT 55.985 2.727 55.99 3.218 ;
      RECT 55.97 2.726 55.985 3.17 ;
      RECT 55.955 2.726 55.97 3.108 ;
      RECT 55.935 2.726 55.955 3.068 ;
      RECT 55.93 2.726 55.935 3.053 ;
      RECT 55.905 2.725 55.93 3.048 ;
      RECT 55.835 2.724 55.905 3.035 ;
      RECT 55.82 2.723 55.835 3.02 ;
      RECT 55.79 2.722 55.82 3.003 ;
      RECT 55.785 2.722 55.79 2.988 ;
      RECT 55.735 2.721 55.785 2.968 ;
      RECT 55.67 2.72 55.735 2.923 ;
      RECT 55.665 2.72 55.67 2.895 ;
      RECT 55.75 3.257 55.755 3.514 ;
      RECT 55.73 3.176 55.75 3.531 ;
      RECT 55.71 3.17 55.73 3.56 ;
      RECT 55.65 3.157 55.71 3.58 ;
      RECT 55.605 3.141 55.65 3.581 ;
      RECT 55.521 3.129 55.605 3.569 ;
      RECT 55.435 3.116 55.521 3.553 ;
      RECT 55.425 3.109 55.435 3.545 ;
      RECT 55.38 3.106 55.425 3.485 ;
      RECT 55.36 3.102 55.38 3.4 ;
      RECT 55.345 3.1 55.36 3.353 ;
      RECT 55.315 3.097 55.345 3.323 ;
      RECT 55.28 3.093 55.315 3.3 ;
      RECT 55.237 3.088 55.28 3.288 ;
      RECT 55.151 3.079 55.237 3.297 ;
      RECT 55.065 3.068 55.151 3.309 ;
      RECT 55 3.059 55.065 3.318 ;
      RECT 54.98 3.05 55 3.323 ;
      RECT 54.975 3.043 54.98 3.325 ;
      RECT 54.935 3.028 54.975 3.322 ;
      RECT 54.915 3.007 54.935 3.317 ;
      RECT 54.9 2.995 54.915 3.31 ;
      RECT 54.895 2.987 54.9 3.303 ;
      RECT 54.88 2.967 54.895 3.296 ;
      RECT 54.875 2.83 54.88 3.29 ;
      RECT 54.795 2.719 54.875 3.262 ;
      RECT 54.786 2.712 54.795 3.228 ;
      RECT 54.7 2.706 54.786 3.153 ;
      RECT 54.675 2.697 54.7 3.065 ;
      RECT 54.645 2.692 54.675 3.04 ;
      RECT 54.58 2.701 54.645 3.025 ;
      RECT 54.56 2.717 54.58 3 ;
      RECT 54.55 2.723 54.56 2.948 ;
      RECT 54.53 2.745 54.55 2.83 ;
      RECT 55.185 2.71 55.355 2.895 ;
      RECT 55.185 2.71 55.39 2.893 ;
      RECT 55.235 2.62 55.405 2.884 ;
      RECT 55.185 2.777 55.41 2.877 ;
      RECT 55.2 2.655 55.405 2.884 ;
      RECT 54.4 3.388 54.465 3.831 ;
      RECT 54.34 3.413 54.465 3.829 ;
      RECT 54.34 3.413 54.52 3.823 ;
      RECT 54.325 3.438 54.52 3.822 ;
      RECT 54.465 3.375 54.54 3.819 ;
      RECT 54.4 3.4 54.62 3.813 ;
      RECT 54.325 3.439 54.665 3.807 ;
      RECT 54.31 3.466 54.665 3.798 ;
      RECT 54.325 3.459 54.685 3.79 ;
      RECT 54.31 3.468 54.69 3.773 ;
      RECT 54.305 3.485 54.69 3.6 ;
      RECT 54.31 2.207 54.345 2.445 ;
      RECT 54.31 2.207 54.375 2.444 ;
      RECT 54.31 2.207 54.49 2.44 ;
      RECT 54.31 2.207 54.545 2.418 ;
      RECT 54.32 2.15 54.6 2.318 ;
      RECT 54.425 1.99 54.455 2.441 ;
      RECT 54.455 1.985 54.635 2.198 ;
      RECT 54.325 2.126 54.635 2.198 ;
      RECT 54.375 2.022 54.425 2.442 ;
      RECT 54.345 2.078 54.635 2.198 ;
      RECT 52.855 1.74 53.025 2.935 ;
      RECT 52.855 1.74 53.32 1.91 ;
      RECT 52.855 6.97 53.32 7.14 ;
      RECT 52.855 5.945 53.025 7.14 ;
      RECT 51.865 1.74 52.035 2.935 ;
      RECT 51.865 1.74 52.33 1.91 ;
      RECT 51.865 6.97 52.33 7.14 ;
      RECT 51.865 5.945 52.035 7.14 ;
      RECT 50.01 2.635 50.18 3.865 ;
      RECT 50.065 0.855 50.235 2.805 ;
      RECT 50.01 0.575 50.18 1.025 ;
      RECT 50.01 7.855 50.18 8.305 ;
      RECT 50.065 6.075 50.235 8.025 ;
      RECT 50.01 5.015 50.18 6.245 ;
      RECT 49.49 0.575 49.66 3.865 ;
      RECT 49.49 2.075 49.895 2.405 ;
      RECT 49.49 1.235 49.895 1.565 ;
      RECT 49.49 5.015 49.66 8.305 ;
      RECT 49.49 7.315 49.895 7.645 ;
      RECT 49.49 6.475 49.895 6.805 ;
      RECT 47.59 3.392 47.605 3.443 ;
      RECT 47.585 3.372 47.59 3.49 ;
      RECT 47.57 3.362 47.585 3.558 ;
      RECT 47.545 3.342 47.57 3.613 ;
      RECT 47.505 3.327 47.545 3.633 ;
      RECT 47.46 3.321 47.505 3.661 ;
      RECT 47.39 3.311 47.46 3.678 ;
      RECT 47.37 3.303 47.39 3.678 ;
      RECT 47.31 3.297 47.37 3.67 ;
      RECT 47.251 3.288 47.31 3.658 ;
      RECT 47.165 3.277 47.251 3.641 ;
      RECT 47.143 3.268 47.165 3.629 ;
      RECT 47.057 3.261 47.143 3.616 ;
      RECT 46.971 3.248 47.057 3.597 ;
      RECT 46.885 3.236 46.971 3.577 ;
      RECT 46.855 3.225 46.885 3.564 ;
      RECT 46.805 3.211 46.855 3.556 ;
      RECT 46.785 3.2 46.805 3.548 ;
      RECT 46.736 3.189 46.785 3.54 ;
      RECT 46.65 3.168 46.736 3.525 ;
      RECT 46.605 3.155 46.65 3.51 ;
      RECT 46.56 3.155 46.605 3.49 ;
      RECT 46.505 3.155 46.56 3.425 ;
      RECT 46.48 3.155 46.505 3.348 ;
      RECT 47.005 2.892 47.175 3.075 ;
      RECT 47.005 2.892 47.19 3.033 ;
      RECT 47.005 2.892 47.195 2.975 ;
      RECT 47.065 2.66 47.2 2.951 ;
      RECT 47.065 2.664 47.205 2.934 ;
      RECT 47.01 2.827 47.205 2.934 ;
      RECT 47.035 2.672 47.175 3.075 ;
      RECT 47.035 2.676 47.215 2.875 ;
      RECT 47.02 2.762 47.215 2.875 ;
      RECT 47.03 2.692 47.175 3.075 ;
      RECT 47.03 2.695 47.225 2.788 ;
      RECT 47.025 2.712 47.225 2.788 ;
      RECT 46.795 1.932 46.965 2.415 ;
      RECT 46.79 1.927 46.94 2.405 ;
      RECT 46.79 1.934 46.97 2.399 ;
      RECT 46.78 1.928 46.94 2.378 ;
      RECT 46.78 1.944 46.985 2.337 ;
      RECT 46.75 1.929 46.94 2.3 ;
      RECT 46.75 1.959 46.995 2.24 ;
      RECT 46.745 1.931 46.94 2.238 ;
      RECT 46.725 1.94 46.97 2.195 ;
      RECT 46.7 1.956 46.985 2.107 ;
      RECT 46.7 1.975 47.01 2.098 ;
      RECT 46.695 2.012 47.01 2.05 ;
      RECT 46.7 1.992 47.015 2.018 ;
      RECT 46.795 1.926 46.905 2.415 ;
      RECT 46.881 1.925 46.905 2.415 ;
      RECT 46.115 2.71 46.12 2.921 ;
      RECT 46.715 2.71 46.72 2.895 ;
      RECT 46.78 2.75 46.785 2.863 ;
      RECT 46.775 2.742 46.78 2.869 ;
      RECT 46.77 2.732 46.775 2.877 ;
      RECT 46.765 2.722 46.77 2.886 ;
      RECT 46.76 2.712 46.765 2.89 ;
      RECT 46.72 2.71 46.76 2.893 ;
      RECT 46.692 2.709 46.715 2.897 ;
      RECT 46.606 2.706 46.692 2.904 ;
      RECT 46.52 2.702 46.606 2.915 ;
      RECT 46.5 2.7 46.52 2.921 ;
      RECT 46.482 2.699 46.5 2.924 ;
      RECT 46.396 2.697 46.482 2.931 ;
      RECT 46.31 2.692 46.396 2.944 ;
      RECT 46.291 2.689 46.31 2.949 ;
      RECT 46.205 2.687 46.291 2.94 ;
      RECT 46.195 2.687 46.205 2.933 ;
      RECT 46.12 2.7 46.195 2.927 ;
      RECT 46.105 2.711 46.115 2.921 ;
      RECT 46.095 2.713 46.105 2.92 ;
      RECT 46.085 2.717 46.095 2.916 ;
      RECT 46.08 2.72 46.085 2.91 ;
      RECT 46.07 2.722 46.08 2.904 ;
      RECT 46.065 2.725 46.07 2.898 ;
      RECT 46.045 3.311 46.05 3.515 ;
      RECT 46.03 3.298 46.045 3.608 ;
      RECT 46.015 3.279 46.03 3.885 ;
      RECT 45.98 3.245 46.015 3.885 ;
      RECT 45.976 3.215 45.98 3.885 ;
      RECT 45.89 3.097 45.976 3.885 ;
      RECT 45.88 2.972 45.89 3.885 ;
      RECT 45.865 2.94 45.88 3.885 ;
      RECT 45.86 2.915 45.865 3.885 ;
      RECT 45.855 2.905 45.86 3.841 ;
      RECT 45.84 2.877 45.855 3.746 ;
      RECT 45.825 2.843 45.84 3.645 ;
      RECT 45.82 2.821 45.825 3.598 ;
      RECT 45.815 2.81 45.82 3.568 ;
      RECT 45.81 2.8 45.815 3.534 ;
      RECT 45.8 2.787 45.81 3.502 ;
      RECT 45.775 2.763 45.8 3.428 ;
      RECT 45.77 2.743 45.775 3.353 ;
      RECT 45.765 2.737 45.77 3.328 ;
      RECT 45.76 2.732 45.765 3.293 ;
      RECT 45.755 2.727 45.76 3.268 ;
      RECT 45.75 2.725 45.755 3.248 ;
      RECT 45.745 2.725 45.75 3.233 ;
      RECT 45.74 2.725 45.745 3.193 ;
      RECT 45.73 2.725 45.74 3.165 ;
      RECT 45.72 2.725 45.73 3.11 ;
      RECT 45.705 2.725 45.72 3.048 ;
      RECT 45.7 2.724 45.705 2.993 ;
      RECT 45.685 2.723 45.7 2.973 ;
      RECT 45.625 2.721 45.685 2.947 ;
      RECT 45.59 2.722 45.625 2.927 ;
      RECT 45.585 2.724 45.59 2.917 ;
      RECT 45.575 2.743 45.585 2.907 ;
      RECT 45.57 2.77 45.575 2.838 ;
      RECT 45.685 2.195 45.855 2.44 ;
      RECT 45.72 1.966 45.855 2.44 ;
      RECT 45.72 1.968 45.865 2.435 ;
      RECT 45.72 1.97 45.89 2.423 ;
      RECT 45.72 1.973 45.915 2.405 ;
      RECT 45.72 1.978 45.965 2.378 ;
      RECT 45.72 1.983 45.985 2.343 ;
      RECT 45.7 1.985 45.995 2.318 ;
      RECT 45.69 2.08 45.995 2.318 ;
      RECT 45.72 1.965 45.83 2.44 ;
      RECT 45.73 1.962 45.825 2.44 ;
      RECT 45.25 3.227 45.44 3.585 ;
      RECT 45.25 3.239 45.475 3.584 ;
      RECT 45.25 3.267 45.495 3.582 ;
      RECT 45.25 3.292 45.5 3.581 ;
      RECT 45.25 3.35 45.515 3.58 ;
      RECT 45.235 3.223 45.395 3.565 ;
      RECT 45.215 3.232 45.44 3.518 ;
      RECT 45.19 3.243 45.475 3.455 ;
      RECT 45.19 3.327 45.51 3.455 ;
      RECT 45.19 3.302 45.505 3.455 ;
      RECT 45.25 3.218 45.395 3.585 ;
      RECT 45.336 3.217 45.395 3.585 ;
      RECT 45.336 3.216 45.38 3.585 ;
      RECT 45.035 2.732 45.04 3.11 ;
      RECT 45.03 2.7 45.035 3.11 ;
      RECT 45.025 2.672 45.03 3.11 ;
      RECT 45.02 2.652 45.025 3.11 ;
      RECT 44.965 2.635 45.02 3.11 ;
      RECT 44.925 2.62 44.965 3.11 ;
      RECT 44.87 2.607 44.925 3.11 ;
      RECT 44.835 2.598 44.87 3.11 ;
      RECT 44.831 2.596 44.835 3.109 ;
      RECT 44.745 2.592 44.831 3.092 ;
      RECT 44.66 2.584 44.745 3.055 ;
      RECT 44.65 2.58 44.66 3.028 ;
      RECT 44.64 2.58 44.65 3.01 ;
      RECT 44.63 2.582 44.64 2.993 ;
      RECT 44.625 2.587 44.63 2.979 ;
      RECT 44.62 2.591 44.625 2.966 ;
      RECT 44.61 2.596 44.62 2.95 ;
      RECT 44.595 2.61 44.61 2.925 ;
      RECT 44.59 2.616 44.595 2.905 ;
      RECT 44.585 2.618 44.59 2.898 ;
      RECT 44.58 2.622 44.585 2.773 ;
      RECT 44.76 3.422 45.005 3.885 ;
      RECT 44.68 3.395 45 3.881 ;
      RECT 44.61 3.43 45.005 3.874 ;
      RECT 44.4 3.685 45.005 3.87 ;
      RECT 44.58 3.453 45.005 3.87 ;
      RECT 44.42 3.645 45.005 3.87 ;
      RECT 44.57 3.465 45.005 3.87 ;
      RECT 44.455 3.582 45.005 3.87 ;
      RECT 44.51 3.507 45.005 3.87 ;
      RECT 44.76 3.372 45 3.885 ;
      RECT 44.79 3.365 45 3.885 ;
      RECT 44.78 3.367 45 3.885 ;
      RECT 44.79 3.362 44.92 3.885 ;
      RECT 44.345 1.925 44.431 2.364 ;
      RECT 44.34 1.925 44.431 2.362 ;
      RECT 44.34 1.925 44.5 2.361 ;
      RECT 44.34 1.925 44.53 2.358 ;
      RECT 44.325 1.932 44.53 2.349 ;
      RECT 44.325 1.932 44.535 2.345 ;
      RECT 44.32 1.942 44.535 2.338 ;
      RECT 44.315 1.947 44.535 2.313 ;
      RECT 44.315 1.947 44.55 2.295 ;
      RECT 44.34 1.925 44.57 2.21 ;
      RECT 44.31 1.952 44.57 2.208 ;
      RECT 44.32 1.945 44.575 2.146 ;
      RECT 44.31 2.067 44.58 2.129 ;
      RECT 44.295 1.962 44.575 2.08 ;
      RECT 44.29 1.972 44.575 1.98 ;
      RECT 44.37 2.743 44.375 2.82 ;
      RECT 44.36 2.737 44.37 3.01 ;
      RECT 44.35 2.729 44.36 3.031 ;
      RECT 44.34 2.72 44.35 3.053 ;
      RECT 44.335 2.715 44.34 3.07 ;
      RECT 44.295 2.715 44.335 3.11 ;
      RECT 44.275 2.715 44.295 3.165 ;
      RECT 44.27 2.715 44.275 3.193 ;
      RECT 44.26 2.715 44.27 3.208 ;
      RECT 44.225 2.715 44.26 3.25 ;
      RECT 44.22 2.715 44.225 3.293 ;
      RECT 44.21 2.715 44.22 3.308 ;
      RECT 44.195 2.715 44.21 3.328 ;
      RECT 44.18 2.715 44.195 3.355 ;
      RECT 44.175 2.716 44.18 3.373 ;
      RECT 44.155 2.717 44.175 3.38 ;
      RECT 44.1 2.718 44.155 3.4 ;
      RECT 44.09 2.719 44.1 3.414 ;
      RECT 44.085 2.722 44.09 3.413 ;
      RECT 44.045 2.795 44.085 3.411 ;
      RECT 44.03 2.875 44.045 3.409 ;
      RECT 44.005 2.93 44.03 3.407 ;
      RECT 43.99 2.995 44.005 3.406 ;
      RECT 43.945 3.027 43.99 3.403 ;
      RECT 43.86 3.05 43.945 3.398 ;
      RECT 43.835 3.07 43.86 3.393 ;
      RECT 43.765 3.075 43.835 3.389 ;
      RECT 43.745 3.077 43.765 3.386 ;
      RECT 43.66 3.088 43.745 3.38 ;
      RECT 43.655 3.099 43.66 3.375 ;
      RECT 43.645 3.101 43.655 3.375 ;
      RECT 43.61 3.105 43.645 3.373 ;
      RECT 43.56 3.115 43.61 3.36 ;
      RECT 43.54 3.123 43.56 3.345 ;
      RECT 43.46 3.135 43.54 3.328 ;
      RECT 43.625 2.685 43.795 2.895 ;
      RECT 43.741 2.681 43.795 2.895 ;
      RECT 43.546 2.685 43.795 2.886 ;
      RECT 43.546 2.685 43.8 2.875 ;
      RECT 43.46 2.685 43.8 2.866 ;
      RECT 43.46 2.693 43.81 2.81 ;
      RECT 43.46 2.705 43.815 2.723 ;
      RECT 43.46 2.712 43.82 2.715 ;
      RECT 43.655 2.683 43.795 2.895 ;
      RECT 43.41 3.628 43.655 3.96 ;
      RECT 43.405 3.62 43.41 3.957 ;
      RECT 43.375 3.64 43.655 3.938 ;
      RECT 43.355 3.672 43.655 3.911 ;
      RECT 43.405 3.625 43.582 3.957 ;
      RECT 43.405 3.622 43.496 3.957 ;
      RECT 43.345 1.97 43.515 2.39 ;
      RECT 43.34 1.97 43.515 2.388 ;
      RECT 43.34 1.97 43.54 2.378 ;
      RECT 43.34 1.97 43.56 2.353 ;
      RECT 43.335 1.97 43.56 2.348 ;
      RECT 43.335 1.97 43.57 2.338 ;
      RECT 43.335 1.97 43.575 2.333 ;
      RECT 43.335 1.975 43.58 2.328 ;
      RECT 43.335 2.007 43.595 2.318 ;
      RECT 43.335 2.077 43.62 2.301 ;
      RECT 43.315 2.077 43.62 2.293 ;
      RECT 43.315 2.137 43.63 2.27 ;
      RECT 43.315 2.177 43.64 2.215 ;
      RECT 43.3 1.97 43.575 2.195 ;
      RECT 43.29 1.985 43.58 2.093 ;
      RECT 42.88 3.375 43.05 3.9 ;
      RECT 42.875 3.375 43.05 3.893 ;
      RECT 42.865 3.375 43.055 3.858 ;
      RECT 42.86 3.385 43.055 3.83 ;
      RECT 42.855 3.405 43.055 3.813 ;
      RECT 42.865 3.38 43.06 3.803 ;
      RECT 42.85 3.425 43.06 3.795 ;
      RECT 42.845 3.445 43.06 3.78 ;
      RECT 42.84 3.475 43.06 3.77 ;
      RECT 42.83 3.52 43.06 3.745 ;
      RECT 42.86 3.39 43.065 3.728 ;
      RECT 42.825 3.572 43.065 3.723 ;
      RECT 42.86 3.4 43.07 3.693 ;
      RECT 42.82 3.605 43.07 3.69 ;
      RECT 42.815 3.63 43.07 3.67 ;
      RECT 42.855 3.417 43.08 3.61 ;
      RECT 42.85 3.439 43.09 3.503 ;
      RECT 42.8 2.686 42.815 2.955 ;
      RECT 42.755 2.67 42.8 3 ;
      RECT 42.75 2.658 42.755 3.05 ;
      RECT 42.74 2.654 42.75 3.083 ;
      RECT 42.735 2.651 42.74 3.111 ;
      RECT 42.72 2.653 42.735 3.153 ;
      RECT 42.715 2.657 42.72 3.193 ;
      RECT 42.695 2.662 42.715 3.245 ;
      RECT 42.691 2.667 42.695 3.302 ;
      RECT 42.605 2.686 42.691 3.339 ;
      RECT 42.595 2.707 42.605 3.375 ;
      RECT 42.59 2.715 42.595 3.376 ;
      RECT 42.585 2.757 42.59 3.377 ;
      RECT 42.57 2.845 42.585 3.378 ;
      RECT 42.56 2.995 42.57 3.38 ;
      RECT 42.555 3.04 42.56 3.382 ;
      RECT 42.52 3.082 42.555 3.385 ;
      RECT 42.515 3.1 42.52 3.388 ;
      RECT 42.438 3.106 42.515 3.394 ;
      RECT 42.352 3.12 42.438 3.407 ;
      RECT 42.266 3.134 42.352 3.421 ;
      RECT 42.18 3.148 42.266 3.434 ;
      RECT 42.12 3.16 42.18 3.446 ;
      RECT 42.095 3.167 42.12 3.453 ;
      RECT 42.081 3.17 42.095 3.458 ;
      RECT 41.995 3.178 42.081 3.474 ;
      RECT 41.99 3.185 41.995 3.489 ;
      RECT 41.966 3.185 41.99 3.496 ;
      RECT 41.88 3.188 41.966 3.524 ;
      RECT 41.795 3.192 41.88 3.568 ;
      RECT 41.73 3.196 41.795 3.605 ;
      RECT 41.705 3.199 41.73 3.621 ;
      RECT 41.63 3.212 41.705 3.625 ;
      RECT 41.605 3.23 41.63 3.629 ;
      RECT 41.595 3.237 41.605 3.631 ;
      RECT 41.58 3.24 41.595 3.632 ;
      RECT 41.52 3.252 41.58 3.636 ;
      RECT 41.51 3.266 41.52 3.64 ;
      RECT 41.455 3.276 41.51 3.628 ;
      RECT 41.43 3.297 41.455 3.611 ;
      RECT 41.41 3.317 41.43 3.602 ;
      RECT 41.405 3.33 41.41 3.597 ;
      RECT 41.39 3.342 41.405 3.593 ;
      RECT 42.625 1.997 42.63 2.02 ;
      RECT 42.62 1.988 42.625 2.06 ;
      RECT 42.615 1.986 42.62 2.103 ;
      RECT 42.61 1.977 42.615 2.138 ;
      RECT 42.605 1.967 42.61 2.21 ;
      RECT 42.6 1.957 42.605 2.275 ;
      RECT 42.595 1.954 42.6 2.315 ;
      RECT 42.57 1.948 42.595 2.405 ;
      RECT 42.535 1.936 42.57 2.43 ;
      RECT 42.525 1.927 42.535 2.43 ;
      RECT 42.39 1.925 42.4 2.413 ;
      RECT 42.38 1.925 42.39 2.38 ;
      RECT 42.375 1.925 42.38 2.355 ;
      RECT 42.37 1.925 42.375 2.343 ;
      RECT 42.365 1.925 42.37 2.325 ;
      RECT 42.355 1.925 42.365 2.29 ;
      RECT 42.35 1.927 42.355 2.268 ;
      RECT 42.345 1.933 42.35 2.253 ;
      RECT 42.34 1.939 42.345 2.238 ;
      RECT 42.325 1.951 42.34 2.211 ;
      RECT 42.32 1.962 42.325 2.179 ;
      RECT 42.315 1.972 42.32 2.163 ;
      RECT 42.305 1.98 42.315 2.132 ;
      RECT 42.3 1.99 42.305 2.106 ;
      RECT 42.295 2.047 42.3 2.089 ;
      RECT 42.4 1.925 42.525 2.43 ;
      RECT 42.115 2.612 42.375 2.91 ;
      RECT 42.11 2.619 42.375 2.908 ;
      RECT 42.115 2.614 42.39 2.903 ;
      RECT 42.105 2.627 42.39 2.9 ;
      RECT 42.105 2.632 42.395 2.893 ;
      RECT 42.1 2.64 42.395 2.89 ;
      RECT 42.1 2.657 42.4 2.688 ;
      RECT 42.115 2.609 42.346 2.91 ;
      RECT 42.17 2.608 42.346 2.91 ;
      RECT 42.17 2.605 42.26 2.91 ;
      RECT 42.17 2.602 42.256 2.91 ;
      RECT 41.86 2.875 41.865 2.888 ;
      RECT 41.855 2.842 41.86 2.893 ;
      RECT 41.85 2.797 41.855 2.9 ;
      RECT 41.845 2.752 41.85 2.908 ;
      RECT 41.84 2.72 41.845 2.916 ;
      RECT 41.835 2.68 41.84 2.917 ;
      RECT 41.82 2.66 41.835 2.919 ;
      RECT 41.745 2.642 41.82 2.931 ;
      RECT 41.735 2.635 41.745 2.942 ;
      RECT 41.73 2.635 41.735 2.944 ;
      RECT 41.7 2.641 41.73 2.948 ;
      RECT 41.66 2.654 41.7 2.948 ;
      RECT 41.635 2.665 41.66 2.934 ;
      RECT 41.62 2.671 41.635 2.917 ;
      RECT 41.61 2.673 41.62 2.908 ;
      RECT 41.605 2.674 41.61 2.903 ;
      RECT 41.6 2.675 41.605 2.898 ;
      RECT 41.595 2.676 41.6 2.895 ;
      RECT 41.57 2.681 41.595 2.885 ;
      RECT 41.56 2.697 41.57 2.872 ;
      RECT 41.555 2.717 41.56 2.867 ;
      RECT 41.565 2.11 41.57 2.306 ;
      RECT 41.55 2.074 41.565 2.308 ;
      RECT 41.54 2.056 41.55 2.313 ;
      RECT 41.53 2.042 41.54 2.317 ;
      RECT 41.485 2.026 41.53 2.327 ;
      RECT 41.48 2.016 41.485 2.336 ;
      RECT 41.435 2.005 41.48 2.342 ;
      RECT 41.43 1.993 41.435 2.349 ;
      RECT 41.415 1.988 41.43 2.353 ;
      RECT 41.4 1.98 41.415 2.358 ;
      RECT 41.39 1.973 41.4 2.363 ;
      RECT 41.38 1.97 41.39 2.368 ;
      RECT 41.37 1.97 41.38 2.369 ;
      RECT 41.365 1.967 41.37 2.368 ;
      RECT 41.33 1.962 41.355 2.367 ;
      RECT 41.306 1.958 41.33 2.366 ;
      RECT 41.22 1.949 41.306 2.363 ;
      RECT 41.205 1.941 41.22 2.36 ;
      RECT 41.183 1.94 41.205 2.359 ;
      RECT 41.097 1.94 41.183 2.357 ;
      RECT 41.011 1.94 41.097 2.355 ;
      RECT 40.925 1.94 41.011 2.352 ;
      RECT 40.915 1.94 40.925 2.343 ;
      RECT 40.885 1.94 40.915 2.303 ;
      RECT 40.875 1.95 40.885 2.258 ;
      RECT 40.87 1.99 40.875 2.243 ;
      RECT 40.865 2.005 40.87 2.23 ;
      RECT 40.835 2.085 40.865 2.192 ;
      RECT 41.355 1.965 41.365 2.368 ;
      RECT 41.18 2.73 41.195 3.335 ;
      RECT 41.185 2.725 41.195 3.335 ;
      RECT 41.35 2.725 41.355 2.908 ;
      RECT 41.34 2.725 41.35 2.938 ;
      RECT 41.325 2.725 41.34 2.998 ;
      RECT 41.32 2.725 41.325 3.043 ;
      RECT 41.315 2.725 41.32 3.073 ;
      RECT 41.31 2.725 41.315 3.093 ;
      RECT 41.3 2.725 41.31 3.128 ;
      RECT 41.285 2.725 41.3 3.16 ;
      RECT 41.24 2.725 41.285 3.188 ;
      RECT 41.235 2.725 41.24 3.218 ;
      RECT 41.23 2.725 41.235 3.23 ;
      RECT 41.225 2.725 41.23 3.238 ;
      RECT 41.215 2.725 41.225 3.253 ;
      RECT 41.21 2.725 41.215 3.275 ;
      RECT 41.2 2.725 41.21 3.298 ;
      RECT 41.195 2.725 41.2 3.318 ;
      RECT 41.16 2.74 41.18 3.335 ;
      RECT 41.135 2.757 41.16 3.335 ;
      RECT 41.13 2.767 41.135 3.335 ;
      RECT 41.1 2.782 41.13 3.335 ;
      RECT 41.025 2.824 41.1 3.335 ;
      RECT 41.02 2.855 41.025 3.318 ;
      RECT 41.015 2.859 41.02 3.3 ;
      RECT 41.01 2.863 41.015 3.263 ;
      RECT 41.005 3.047 41.01 3.23 ;
      RECT 40.49 3.236 40.576 3.801 ;
      RECT 40.445 3.238 40.61 3.795 ;
      RECT 40.576 3.235 40.61 3.795 ;
      RECT 40.49 3.237 40.695 3.789 ;
      RECT 40.445 3.247 40.705 3.785 ;
      RECT 40.42 3.239 40.695 3.781 ;
      RECT 40.415 3.242 40.695 3.776 ;
      RECT 40.39 3.257 40.705 3.77 ;
      RECT 40.39 3.282 40.745 3.765 ;
      RECT 40.35 3.29 40.745 3.74 ;
      RECT 40.35 3.317 40.76 3.738 ;
      RECT 40.35 3.347 40.77 3.725 ;
      RECT 40.345 3.492 40.77 3.713 ;
      RECT 40.35 3.421 40.79 3.71 ;
      RECT 40.35 3.478 40.795 3.518 ;
      RECT 40.54 2.757 40.71 2.935 ;
      RECT 40.49 2.696 40.54 2.92 ;
      RECT 40.225 2.676 40.49 2.905 ;
      RECT 40.185 2.74 40.66 2.905 ;
      RECT 40.185 2.73 40.615 2.905 ;
      RECT 40.185 2.727 40.605 2.905 ;
      RECT 40.185 2.715 40.595 2.905 ;
      RECT 40.185 2.7 40.54 2.905 ;
      RECT 40.225 2.672 40.426 2.905 ;
      RECT 40.235 2.65 40.426 2.905 ;
      RECT 40.26 2.635 40.34 2.905 ;
      RECT 40.015 3.165 40.135 3.61 ;
      RECT 40 3.165 40.135 3.609 ;
      RECT 39.955 3.187 40.135 3.604 ;
      RECT 39.915 3.236 40.135 3.598 ;
      RECT 39.915 3.236 40.14 3.573 ;
      RECT 39.915 3.236 40.16 3.463 ;
      RECT 39.91 3.266 40.16 3.46 ;
      RECT 40 3.165 40.17 3.355 ;
      RECT 39.66 1.95 39.665 2.395 ;
      RECT 39.47 1.95 39.49 2.36 ;
      RECT 39.44 1.95 39.445 2.335 ;
      RECT 40.12 2.257 40.135 2.445 ;
      RECT 40.115 2.242 40.12 2.451 ;
      RECT 40.095 2.215 40.115 2.454 ;
      RECT 40.045 2.182 40.095 2.463 ;
      RECT 40.015 2.162 40.045 2.467 ;
      RECT 39.996 2.15 40.015 2.463 ;
      RECT 39.91 2.122 39.996 2.453 ;
      RECT 39.9 2.097 39.91 2.443 ;
      RECT 39.83 2.065 39.9 2.435 ;
      RECT 39.805 2.025 39.83 2.427 ;
      RECT 39.785 2.007 39.805 2.421 ;
      RECT 39.775 1.997 39.785 2.418 ;
      RECT 39.765 1.99 39.775 2.416 ;
      RECT 39.745 1.977 39.765 2.413 ;
      RECT 39.735 1.967 39.745 2.41 ;
      RECT 39.725 1.96 39.735 2.408 ;
      RECT 39.675 1.952 39.725 2.402 ;
      RECT 39.665 1.95 39.675 2.396 ;
      RECT 39.635 1.95 39.66 2.393 ;
      RECT 39.606 1.95 39.635 2.388 ;
      RECT 39.52 1.95 39.606 2.378 ;
      RECT 39.49 1.95 39.52 2.365 ;
      RECT 39.445 1.95 39.47 2.348 ;
      RECT 39.43 1.95 39.44 2.33 ;
      RECT 39.41 1.957 39.43 2.315 ;
      RECT 39.405 1.972 39.41 2.303 ;
      RECT 39.4 1.977 39.405 2.243 ;
      RECT 39.395 1.982 39.4 2.085 ;
      RECT 39.39 1.985 39.395 2.003 ;
      RECT 39.655 2.67 39.741 2.991 ;
      RECT 39.655 2.67 39.775 2.984 ;
      RECT 39.605 2.67 39.775 2.98 ;
      RECT 39.605 2.672 39.861 2.978 ;
      RECT 39.605 2.674 39.885 2.972 ;
      RECT 39.605 2.681 39.895 2.971 ;
      RECT 39.605 2.69 39.9 2.968 ;
      RECT 39.605 2.696 39.905 2.963 ;
      RECT 39.605 2.74 39.91 2.96 ;
      RECT 39.605 2.832 39.915 2.957 ;
      RECT 39.13 3.275 39.165 3.595 ;
      RECT 39.715 3.46 39.72 3.642 ;
      RECT 39.67 3.342 39.715 3.661 ;
      RECT 39.655 3.319 39.67 3.684 ;
      RECT 39.645 3.309 39.655 3.694 ;
      RECT 39.625 3.304 39.645 3.707 ;
      RECT 39.6 3.302 39.625 3.728 ;
      RECT 39.581 3.301 39.6 3.74 ;
      RECT 39.495 3.298 39.581 3.74 ;
      RECT 39.425 3.293 39.495 3.728 ;
      RECT 39.35 3.289 39.425 3.703 ;
      RECT 39.285 3.285 39.35 3.67 ;
      RECT 39.215 3.282 39.285 3.63 ;
      RECT 39.185 3.278 39.215 3.605 ;
      RECT 39.165 3.276 39.185 3.598 ;
      RECT 39.081 3.274 39.13 3.596 ;
      RECT 38.995 3.271 39.081 3.597 ;
      RECT 38.92 3.27 38.995 3.599 ;
      RECT 38.835 3.27 38.92 3.625 ;
      RECT 38.758 3.271 38.835 3.65 ;
      RECT 38.672 3.272 38.758 3.65 ;
      RECT 38.586 3.272 38.672 3.65 ;
      RECT 38.5 3.273 38.586 3.65 ;
      RECT 38.48 3.274 38.5 3.642 ;
      RECT 38.465 3.28 38.48 3.627 ;
      RECT 38.43 3.3 38.465 3.607 ;
      RECT 38.42 3.32 38.43 3.589 ;
      RECT 39.39 2.625 39.395 2.895 ;
      RECT 39.385 2.616 39.39 2.9 ;
      RECT 39.375 2.606 39.385 2.912 ;
      RECT 39.37 2.595 39.375 2.923 ;
      RECT 39.35 2.589 39.37 2.941 ;
      RECT 39.305 2.586 39.35 2.99 ;
      RECT 39.29 2.585 39.305 3.035 ;
      RECT 39.285 2.585 39.29 3.048 ;
      RECT 39.275 2.585 39.285 3.06 ;
      RECT 39.27 2.586 39.275 3.075 ;
      RECT 39.25 2.594 39.27 3.08 ;
      RECT 39.22 2.61 39.25 3.08 ;
      RECT 39.21 2.622 39.215 3.08 ;
      RECT 39.175 2.637 39.21 3.08 ;
      RECT 39.145 2.657 39.175 3.08 ;
      RECT 39.135 2.682 39.145 3.08 ;
      RECT 39.13 2.71 39.135 3.08 ;
      RECT 39.125 2.74 39.13 3.08 ;
      RECT 39.12 2.757 39.125 3.08 ;
      RECT 39.11 2.785 39.12 3.08 ;
      RECT 39.1 2.82 39.11 3.08 ;
      RECT 39.095 2.855 39.1 3.08 ;
      RECT 39.215 2.62 39.22 3.08 ;
      RECT 38.73 2.722 38.915 2.895 ;
      RECT 38.69 2.64 38.875 2.893 ;
      RECT 38.651 2.645 38.875 2.889 ;
      RECT 38.565 2.654 38.875 2.884 ;
      RECT 38.481 2.67 38.88 2.879 ;
      RECT 38.395 2.69 38.905 2.873 ;
      RECT 38.395 2.71 38.91 2.873 ;
      RECT 38.481 2.68 38.905 2.879 ;
      RECT 38.565 2.655 38.88 2.884 ;
      RECT 38.73 2.637 38.875 2.895 ;
      RECT 38.73 2.632 38.83 2.895 ;
      RECT 38.816 2.626 38.83 2.895 ;
      RECT 38.205 1.95 38.21 2.349 ;
      RECT 37.95 1.95 37.985 2.347 ;
      RECT 37.545 1.985 37.55 2.341 ;
      RECT 38.29 1.988 38.295 2.243 ;
      RECT 38.285 1.986 38.29 2.249 ;
      RECT 38.28 1.985 38.285 2.256 ;
      RECT 38.255 1.978 38.28 2.28 ;
      RECT 38.25 1.971 38.255 2.304 ;
      RECT 38.245 1.967 38.25 2.313 ;
      RECT 38.235 1.962 38.245 2.326 ;
      RECT 38.23 1.959 38.235 2.335 ;
      RECT 38.225 1.957 38.23 2.34 ;
      RECT 38.21 1.953 38.225 2.35 ;
      RECT 38.195 1.947 38.205 2.349 ;
      RECT 38.157 1.945 38.195 2.349 ;
      RECT 38.071 1.947 38.157 2.349 ;
      RECT 37.985 1.949 38.071 2.348 ;
      RECT 37.914 1.95 37.95 2.347 ;
      RECT 37.828 1.952 37.914 2.347 ;
      RECT 37.742 1.954 37.828 2.346 ;
      RECT 37.656 1.956 37.742 2.346 ;
      RECT 37.57 1.959 37.656 2.345 ;
      RECT 37.56 1.965 37.57 2.344 ;
      RECT 37.55 1.977 37.56 2.342 ;
      RECT 37.49 2.012 37.545 2.338 ;
      RECT 37.485 2.042 37.49 2.1 ;
      RECT 38.23 3.122 38.245 3.315 ;
      RECT 38.225 3.09 38.23 3.315 ;
      RECT 38.215 3.065 38.225 3.315 ;
      RECT 38.21 3.037 38.215 3.315 ;
      RECT 38.18 2.96 38.21 3.315 ;
      RECT 38.155 2.842 38.18 3.315 ;
      RECT 38.15 2.78 38.155 3.315 ;
      RECT 38.14 2.767 38.15 3.315 ;
      RECT 38.12 2.757 38.14 3.315 ;
      RECT 38.105 2.74 38.12 3.315 ;
      RECT 38.075 2.728 38.105 3.315 ;
      RECT 38.07 2.727 38.075 3.26 ;
      RECT 38.065 2.727 38.07 3.218 ;
      RECT 38.05 2.726 38.065 3.17 ;
      RECT 38.035 2.726 38.05 3.108 ;
      RECT 38.015 2.726 38.035 3.068 ;
      RECT 38.01 2.726 38.015 3.053 ;
      RECT 37.985 2.725 38.01 3.048 ;
      RECT 37.915 2.724 37.985 3.035 ;
      RECT 37.9 2.723 37.915 3.02 ;
      RECT 37.87 2.722 37.9 3.003 ;
      RECT 37.865 2.722 37.87 2.988 ;
      RECT 37.815 2.721 37.865 2.968 ;
      RECT 37.75 2.72 37.815 2.923 ;
      RECT 37.745 2.72 37.75 2.895 ;
      RECT 37.83 3.257 37.835 3.514 ;
      RECT 37.81 3.176 37.83 3.531 ;
      RECT 37.79 3.17 37.81 3.56 ;
      RECT 37.73 3.157 37.79 3.58 ;
      RECT 37.685 3.141 37.73 3.581 ;
      RECT 37.601 3.129 37.685 3.569 ;
      RECT 37.515 3.116 37.601 3.553 ;
      RECT 37.505 3.109 37.515 3.545 ;
      RECT 37.46 3.106 37.505 3.485 ;
      RECT 37.44 3.102 37.46 3.4 ;
      RECT 37.425 3.1 37.44 3.353 ;
      RECT 37.395 3.097 37.425 3.323 ;
      RECT 37.36 3.093 37.395 3.3 ;
      RECT 37.317 3.088 37.36 3.288 ;
      RECT 37.231 3.079 37.317 3.297 ;
      RECT 37.145 3.068 37.231 3.309 ;
      RECT 37.08 3.059 37.145 3.318 ;
      RECT 37.06 3.05 37.08 3.323 ;
      RECT 37.055 3.043 37.06 3.325 ;
      RECT 37.015 3.028 37.055 3.322 ;
      RECT 36.995 3.007 37.015 3.317 ;
      RECT 36.98 2.995 36.995 3.31 ;
      RECT 36.975 2.987 36.98 3.303 ;
      RECT 36.96 2.967 36.975 3.296 ;
      RECT 36.955 2.83 36.96 3.29 ;
      RECT 36.875 2.719 36.955 3.262 ;
      RECT 36.866 2.712 36.875 3.228 ;
      RECT 36.78 2.706 36.866 3.153 ;
      RECT 36.755 2.697 36.78 3.065 ;
      RECT 36.725 2.692 36.755 3.04 ;
      RECT 36.66 2.701 36.725 3.025 ;
      RECT 36.64 2.717 36.66 3 ;
      RECT 36.63 2.723 36.64 2.948 ;
      RECT 36.61 2.745 36.63 2.83 ;
      RECT 37.265 2.71 37.435 2.895 ;
      RECT 37.265 2.71 37.47 2.893 ;
      RECT 37.315 2.62 37.485 2.884 ;
      RECT 37.265 2.777 37.49 2.877 ;
      RECT 37.28 2.655 37.485 2.884 ;
      RECT 36.48 3.388 36.545 3.831 ;
      RECT 36.42 3.413 36.545 3.829 ;
      RECT 36.42 3.413 36.6 3.823 ;
      RECT 36.405 3.438 36.6 3.822 ;
      RECT 36.545 3.375 36.62 3.819 ;
      RECT 36.48 3.4 36.7 3.813 ;
      RECT 36.405 3.439 36.745 3.807 ;
      RECT 36.39 3.466 36.745 3.798 ;
      RECT 36.405 3.459 36.765 3.79 ;
      RECT 36.39 3.468 36.77 3.773 ;
      RECT 36.385 3.485 36.77 3.6 ;
      RECT 36.39 2.207 36.425 2.445 ;
      RECT 36.39 2.207 36.455 2.444 ;
      RECT 36.39 2.207 36.57 2.44 ;
      RECT 36.39 2.207 36.625 2.418 ;
      RECT 36.4 2.15 36.68 2.318 ;
      RECT 36.505 1.99 36.535 2.441 ;
      RECT 36.535 1.985 36.715 2.198 ;
      RECT 36.405 2.126 36.715 2.198 ;
      RECT 36.455 2.022 36.505 2.442 ;
      RECT 36.425 2.078 36.715 2.198 ;
      RECT 34.94 1.74 35.11 2.935 ;
      RECT 34.94 1.74 35.405 1.91 ;
      RECT 34.94 6.97 35.405 7.14 ;
      RECT 34.94 5.945 35.11 7.14 ;
      RECT 33.95 1.74 34.12 2.935 ;
      RECT 33.95 1.74 34.415 1.91 ;
      RECT 33.95 6.97 34.415 7.14 ;
      RECT 33.95 5.945 34.12 7.14 ;
      RECT 32.095 2.635 32.265 3.865 ;
      RECT 32.15 0.855 32.32 2.805 ;
      RECT 32.095 0.575 32.265 1.025 ;
      RECT 32.095 7.855 32.265 8.305 ;
      RECT 32.15 6.075 32.32 8.025 ;
      RECT 32.095 5.015 32.265 6.245 ;
      RECT 31.575 0.575 31.745 3.865 ;
      RECT 31.575 2.075 31.98 2.405 ;
      RECT 31.575 1.235 31.98 1.565 ;
      RECT 31.575 5.015 31.745 8.305 ;
      RECT 31.575 7.315 31.98 7.645 ;
      RECT 31.575 6.475 31.98 6.805 ;
      RECT 29.675 3.392 29.69 3.443 ;
      RECT 29.67 3.372 29.675 3.49 ;
      RECT 29.655 3.362 29.67 3.558 ;
      RECT 29.63 3.342 29.655 3.613 ;
      RECT 29.59 3.327 29.63 3.633 ;
      RECT 29.545 3.321 29.59 3.661 ;
      RECT 29.475 3.311 29.545 3.678 ;
      RECT 29.455 3.303 29.475 3.678 ;
      RECT 29.395 3.297 29.455 3.67 ;
      RECT 29.336 3.288 29.395 3.658 ;
      RECT 29.25 3.277 29.336 3.641 ;
      RECT 29.228 3.268 29.25 3.629 ;
      RECT 29.142 3.261 29.228 3.616 ;
      RECT 29.056 3.248 29.142 3.597 ;
      RECT 28.97 3.236 29.056 3.577 ;
      RECT 28.94 3.225 28.97 3.564 ;
      RECT 28.89 3.211 28.94 3.556 ;
      RECT 28.87 3.2 28.89 3.548 ;
      RECT 28.821 3.189 28.87 3.54 ;
      RECT 28.735 3.168 28.821 3.525 ;
      RECT 28.69 3.155 28.735 3.51 ;
      RECT 28.645 3.155 28.69 3.49 ;
      RECT 28.59 3.155 28.645 3.425 ;
      RECT 28.565 3.155 28.59 3.348 ;
      RECT 29.09 2.892 29.26 3.075 ;
      RECT 29.09 2.892 29.275 3.033 ;
      RECT 29.09 2.892 29.28 2.975 ;
      RECT 29.15 2.66 29.285 2.951 ;
      RECT 29.15 2.664 29.29 2.934 ;
      RECT 29.095 2.827 29.29 2.934 ;
      RECT 29.12 2.672 29.26 3.075 ;
      RECT 29.12 2.676 29.3 2.875 ;
      RECT 29.105 2.762 29.3 2.875 ;
      RECT 29.115 2.692 29.26 3.075 ;
      RECT 29.115 2.695 29.31 2.788 ;
      RECT 29.11 2.712 29.31 2.788 ;
      RECT 28.88 1.932 29.05 2.415 ;
      RECT 28.875 1.927 29.025 2.405 ;
      RECT 28.875 1.934 29.055 2.399 ;
      RECT 28.865 1.928 29.025 2.378 ;
      RECT 28.865 1.944 29.07 2.337 ;
      RECT 28.835 1.929 29.025 2.3 ;
      RECT 28.835 1.959 29.08 2.24 ;
      RECT 28.83 1.931 29.025 2.238 ;
      RECT 28.81 1.94 29.055 2.195 ;
      RECT 28.785 1.956 29.07 2.107 ;
      RECT 28.785 1.975 29.095 2.098 ;
      RECT 28.78 2.012 29.095 2.05 ;
      RECT 28.785 1.992 29.1 2.018 ;
      RECT 28.88 1.926 28.99 2.415 ;
      RECT 28.966 1.925 28.99 2.415 ;
      RECT 28.2 2.71 28.205 2.921 ;
      RECT 28.8 2.71 28.805 2.895 ;
      RECT 28.865 2.75 28.87 2.863 ;
      RECT 28.86 2.742 28.865 2.869 ;
      RECT 28.855 2.732 28.86 2.877 ;
      RECT 28.85 2.722 28.855 2.886 ;
      RECT 28.845 2.712 28.85 2.89 ;
      RECT 28.805 2.71 28.845 2.893 ;
      RECT 28.777 2.709 28.8 2.897 ;
      RECT 28.691 2.706 28.777 2.904 ;
      RECT 28.605 2.702 28.691 2.915 ;
      RECT 28.585 2.7 28.605 2.921 ;
      RECT 28.567 2.699 28.585 2.924 ;
      RECT 28.481 2.697 28.567 2.931 ;
      RECT 28.395 2.692 28.481 2.944 ;
      RECT 28.376 2.689 28.395 2.949 ;
      RECT 28.29 2.687 28.376 2.94 ;
      RECT 28.28 2.687 28.29 2.933 ;
      RECT 28.205 2.7 28.28 2.927 ;
      RECT 28.19 2.711 28.2 2.921 ;
      RECT 28.18 2.713 28.19 2.92 ;
      RECT 28.17 2.717 28.18 2.916 ;
      RECT 28.165 2.72 28.17 2.91 ;
      RECT 28.155 2.722 28.165 2.904 ;
      RECT 28.15 2.725 28.155 2.898 ;
      RECT 28.13 3.311 28.135 3.515 ;
      RECT 28.115 3.298 28.13 3.608 ;
      RECT 28.1 3.279 28.115 3.885 ;
      RECT 28.065 3.245 28.1 3.885 ;
      RECT 28.061 3.215 28.065 3.885 ;
      RECT 27.975 3.097 28.061 3.885 ;
      RECT 27.965 2.972 27.975 3.885 ;
      RECT 27.95 2.94 27.965 3.885 ;
      RECT 27.945 2.915 27.95 3.885 ;
      RECT 27.94 2.905 27.945 3.841 ;
      RECT 27.925 2.877 27.94 3.746 ;
      RECT 27.91 2.843 27.925 3.645 ;
      RECT 27.905 2.821 27.91 3.598 ;
      RECT 27.9 2.81 27.905 3.568 ;
      RECT 27.895 2.8 27.9 3.534 ;
      RECT 27.885 2.787 27.895 3.502 ;
      RECT 27.86 2.763 27.885 3.428 ;
      RECT 27.855 2.743 27.86 3.353 ;
      RECT 27.85 2.737 27.855 3.328 ;
      RECT 27.845 2.732 27.85 3.293 ;
      RECT 27.84 2.727 27.845 3.268 ;
      RECT 27.835 2.725 27.84 3.248 ;
      RECT 27.83 2.725 27.835 3.233 ;
      RECT 27.825 2.725 27.83 3.193 ;
      RECT 27.815 2.725 27.825 3.165 ;
      RECT 27.805 2.725 27.815 3.11 ;
      RECT 27.79 2.725 27.805 3.048 ;
      RECT 27.785 2.724 27.79 2.993 ;
      RECT 27.77 2.723 27.785 2.973 ;
      RECT 27.71 2.721 27.77 2.947 ;
      RECT 27.675 2.722 27.71 2.927 ;
      RECT 27.67 2.724 27.675 2.917 ;
      RECT 27.66 2.743 27.67 2.907 ;
      RECT 27.655 2.77 27.66 2.838 ;
      RECT 27.77 2.195 27.94 2.44 ;
      RECT 27.805 1.966 27.94 2.44 ;
      RECT 27.805 1.968 27.95 2.435 ;
      RECT 27.805 1.97 27.975 2.423 ;
      RECT 27.805 1.973 28 2.405 ;
      RECT 27.805 1.978 28.05 2.378 ;
      RECT 27.805 1.983 28.07 2.343 ;
      RECT 27.785 1.985 28.08 2.318 ;
      RECT 27.775 2.08 28.08 2.318 ;
      RECT 27.805 1.965 27.915 2.44 ;
      RECT 27.815 1.962 27.91 2.44 ;
      RECT 27.335 3.227 27.525 3.585 ;
      RECT 27.335 3.239 27.56 3.584 ;
      RECT 27.335 3.267 27.58 3.582 ;
      RECT 27.335 3.292 27.585 3.581 ;
      RECT 27.335 3.35 27.6 3.58 ;
      RECT 27.32 3.223 27.48 3.565 ;
      RECT 27.3 3.232 27.525 3.518 ;
      RECT 27.275 3.243 27.56 3.455 ;
      RECT 27.275 3.327 27.595 3.455 ;
      RECT 27.275 3.302 27.59 3.455 ;
      RECT 27.335 3.218 27.48 3.585 ;
      RECT 27.421 3.217 27.48 3.585 ;
      RECT 27.421 3.216 27.465 3.585 ;
      RECT 27.12 2.732 27.125 3.11 ;
      RECT 27.115 2.7 27.12 3.11 ;
      RECT 27.11 2.672 27.115 3.11 ;
      RECT 27.105 2.652 27.11 3.11 ;
      RECT 27.05 2.635 27.105 3.11 ;
      RECT 27.01 2.62 27.05 3.11 ;
      RECT 26.955 2.607 27.01 3.11 ;
      RECT 26.92 2.598 26.955 3.11 ;
      RECT 26.916 2.596 26.92 3.109 ;
      RECT 26.83 2.592 26.916 3.092 ;
      RECT 26.745 2.584 26.83 3.055 ;
      RECT 26.735 2.58 26.745 3.028 ;
      RECT 26.725 2.58 26.735 3.01 ;
      RECT 26.715 2.582 26.725 2.993 ;
      RECT 26.71 2.587 26.715 2.979 ;
      RECT 26.705 2.591 26.71 2.966 ;
      RECT 26.695 2.596 26.705 2.95 ;
      RECT 26.68 2.61 26.695 2.925 ;
      RECT 26.675 2.616 26.68 2.905 ;
      RECT 26.67 2.618 26.675 2.898 ;
      RECT 26.665 2.622 26.67 2.773 ;
      RECT 26.845 3.422 27.09 3.885 ;
      RECT 26.765 3.395 27.085 3.881 ;
      RECT 26.695 3.43 27.09 3.874 ;
      RECT 26.485 3.685 27.09 3.87 ;
      RECT 26.665 3.453 27.09 3.87 ;
      RECT 26.505 3.645 27.09 3.87 ;
      RECT 26.655 3.465 27.09 3.87 ;
      RECT 26.54 3.582 27.09 3.87 ;
      RECT 26.595 3.507 27.09 3.87 ;
      RECT 26.845 3.372 27.085 3.885 ;
      RECT 26.875 3.365 27.085 3.885 ;
      RECT 26.865 3.367 27.085 3.885 ;
      RECT 26.875 3.362 27.005 3.885 ;
      RECT 26.43 1.925 26.516 2.364 ;
      RECT 26.425 1.925 26.516 2.362 ;
      RECT 26.425 1.925 26.585 2.361 ;
      RECT 26.425 1.925 26.615 2.358 ;
      RECT 26.41 1.932 26.615 2.349 ;
      RECT 26.41 1.932 26.62 2.345 ;
      RECT 26.405 1.942 26.62 2.338 ;
      RECT 26.4 1.947 26.62 2.313 ;
      RECT 26.4 1.947 26.635 2.295 ;
      RECT 26.425 1.925 26.655 2.21 ;
      RECT 26.395 1.952 26.655 2.208 ;
      RECT 26.405 1.945 26.66 2.146 ;
      RECT 26.395 2.067 26.665 2.129 ;
      RECT 26.38 1.962 26.66 2.08 ;
      RECT 26.375 1.972 26.66 1.98 ;
      RECT 26.455 2.743 26.46 2.82 ;
      RECT 26.445 2.737 26.455 3.01 ;
      RECT 26.435 2.729 26.445 3.031 ;
      RECT 26.425 2.72 26.435 3.053 ;
      RECT 26.42 2.715 26.425 3.07 ;
      RECT 26.38 2.715 26.42 3.11 ;
      RECT 26.36 2.715 26.38 3.165 ;
      RECT 26.355 2.715 26.36 3.193 ;
      RECT 26.345 2.715 26.355 3.208 ;
      RECT 26.31 2.715 26.345 3.25 ;
      RECT 26.305 2.715 26.31 3.293 ;
      RECT 26.295 2.715 26.305 3.308 ;
      RECT 26.28 2.715 26.295 3.328 ;
      RECT 26.265 2.715 26.28 3.355 ;
      RECT 26.26 2.716 26.265 3.373 ;
      RECT 26.24 2.717 26.26 3.38 ;
      RECT 26.185 2.718 26.24 3.4 ;
      RECT 26.175 2.719 26.185 3.414 ;
      RECT 26.17 2.722 26.175 3.413 ;
      RECT 26.13 2.795 26.17 3.411 ;
      RECT 26.115 2.875 26.13 3.409 ;
      RECT 26.09 2.93 26.115 3.407 ;
      RECT 26.075 2.995 26.09 3.406 ;
      RECT 26.03 3.027 26.075 3.403 ;
      RECT 25.945 3.05 26.03 3.398 ;
      RECT 25.92 3.07 25.945 3.393 ;
      RECT 25.85 3.075 25.92 3.389 ;
      RECT 25.83 3.077 25.85 3.386 ;
      RECT 25.745 3.088 25.83 3.38 ;
      RECT 25.74 3.099 25.745 3.375 ;
      RECT 25.73 3.101 25.74 3.375 ;
      RECT 25.695 3.105 25.73 3.373 ;
      RECT 25.645 3.115 25.695 3.36 ;
      RECT 25.625 3.123 25.645 3.345 ;
      RECT 25.545 3.135 25.625 3.328 ;
      RECT 25.71 2.685 25.88 2.895 ;
      RECT 25.826 2.681 25.88 2.895 ;
      RECT 25.631 2.685 25.88 2.886 ;
      RECT 25.631 2.685 25.885 2.875 ;
      RECT 25.545 2.685 25.885 2.866 ;
      RECT 25.545 2.693 25.895 2.81 ;
      RECT 25.545 2.705 25.9 2.723 ;
      RECT 25.545 2.712 25.905 2.715 ;
      RECT 25.74 2.683 25.88 2.895 ;
      RECT 25.495 3.628 25.74 3.96 ;
      RECT 25.49 3.62 25.495 3.957 ;
      RECT 25.46 3.64 25.74 3.938 ;
      RECT 25.44 3.672 25.74 3.911 ;
      RECT 25.49 3.625 25.667 3.957 ;
      RECT 25.49 3.622 25.581 3.957 ;
      RECT 25.43 1.97 25.6 2.39 ;
      RECT 25.425 1.97 25.6 2.388 ;
      RECT 25.425 1.97 25.625 2.378 ;
      RECT 25.425 1.97 25.645 2.353 ;
      RECT 25.42 1.97 25.645 2.348 ;
      RECT 25.42 1.97 25.655 2.338 ;
      RECT 25.42 1.97 25.66 2.333 ;
      RECT 25.42 1.975 25.665 2.328 ;
      RECT 25.42 2.007 25.68 2.318 ;
      RECT 25.42 2.077 25.705 2.301 ;
      RECT 25.4 2.077 25.705 2.293 ;
      RECT 25.4 2.137 25.715 2.27 ;
      RECT 25.4 2.177 25.725 2.215 ;
      RECT 25.385 1.97 25.66 2.195 ;
      RECT 25.375 1.985 25.665 2.093 ;
      RECT 24.965 3.375 25.135 3.9 ;
      RECT 24.96 3.375 25.135 3.893 ;
      RECT 24.95 3.375 25.14 3.858 ;
      RECT 24.945 3.385 25.14 3.83 ;
      RECT 24.94 3.405 25.14 3.813 ;
      RECT 24.95 3.38 25.145 3.803 ;
      RECT 24.935 3.425 25.145 3.795 ;
      RECT 24.93 3.445 25.145 3.78 ;
      RECT 24.925 3.475 25.145 3.77 ;
      RECT 24.915 3.52 25.145 3.745 ;
      RECT 24.945 3.39 25.15 3.728 ;
      RECT 24.91 3.572 25.15 3.723 ;
      RECT 24.945 3.4 25.155 3.693 ;
      RECT 24.905 3.605 25.155 3.69 ;
      RECT 24.9 3.63 25.155 3.67 ;
      RECT 24.94 3.417 25.165 3.61 ;
      RECT 24.935 3.439 25.175 3.503 ;
      RECT 24.885 2.686 24.9 2.955 ;
      RECT 24.84 2.67 24.885 3 ;
      RECT 24.835 2.658 24.84 3.05 ;
      RECT 24.825 2.654 24.835 3.083 ;
      RECT 24.82 2.651 24.825 3.111 ;
      RECT 24.805 2.653 24.82 3.153 ;
      RECT 24.8 2.657 24.805 3.193 ;
      RECT 24.78 2.662 24.8 3.245 ;
      RECT 24.776 2.667 24.78 3.302 ;
      RECT 24.69 2.686 24.776 3.339 ;
      RECT 24.68 2.707 24.69 3.375 ;
      RECT 24.675 2.715 24.68 3.376 ;
      RECT 24.67 2.757 24.675 3.377 ;
      RECT 24.655 2.845 24.67 3.378 ;
      RECT 24.645 2.995 24.655 3.38 ;
      RECT 24.64 3.04 24.645 3.382 ;
      RECT 24.605 3.082 24.64 3.385 ;
      RECT 24.6 3.1 24.605 3.388 ;
      RECT 24.523 3.106 24.6 3.394 ;
      RECT 24.437 3.12 24.523 3.407 ;
      RECT 24.351 3.134 24.437 3.421 ;
      RECT 24.265 3.148 24.351 3.434 ;
      RECT 24.205 3.16 24.265 3.446 ;
      RECT 24.18 3.167 24.205 3.453 ;
      RECT 24.166 3.17 24.18 3.458 ;
      RECT 24.08 3.178 24.166 3.474 ;
      RECT 24.075 3.185 24.08 3.489 ;
      RECT 24.051 3.185 24.075 3.496 ;
      RECT 23.965 3.188 24.051 3.524 ;
      RECT 23.88 3.192 23.965 3.568 ;
      RECT 23.815 3.196 23.88 3.605 ;
      RECT 23.79 3.199 23.815 3.621 ;
      RECT 23.715 3.212 23.79 3.625 ;
      RECT 23.69 3.23 23.715 3.629 ;
      RECT 23.68 3.237 23.69 3.631 ;
      RECT 23.665 3.24 23.68 3.632 ;
      RECT 23.605 3.252 23.665 3.636 ;
      RECT 23.595 3.266 23.605 3.64 ;
      RECT 23.54 3.276 23.595 3.628 ;
      RECT 23.515 3.297 23.54 3.611 ;
      RECT 23.495 3.317 23.515 3.602 ;
      RECT 23.49 3.33 23.495 3.597 ;
      RECT 23.475 3.342 23.49 3.593 ;
      RECT 24.71 1.997 24.715 2.02 ;
      RECT 24.705 1.988 24.71 2.06 ;
      RECT 24.7 1.986 24.705 2.103 ;
      RECT 24.695 1.977 24.7 2.138 ;
      RECT 24.69 1.967 24.695 2.21 ;
      RECT 24.685 1.957 24.69 2.275 ;
      RECT 24.68 1.954 24.685 2.315 ;
      RECT 24.655 1.948 24.68 2.405 ;
      RECT 24.62 1.936 24.655 2.43 ;
      RECT 24.61 1.927 24.62 2.43 ;
      RECT 24.475 1.925 24.485 2.413 ;
      RECT 24.465 1.925 24.475 2.38 ;
      RECT 24.46 1.925 24.465 2.355 ;
      RECT 24.455 1.925 24.46 2.343 ;
      RECT 24.45 1.925 24.455 2.325 ;
      RECT 24.44 1.925 24.45 2.29 ;
      RECT 24.435 1.927 24.44 2.268 ;
      RECT 24.43 1.933 24.435 2.253 ;
      RECT 24.425 1.939 24.43 2.238 ;
      RECT 24.41 1.951 24.425 2.211 ;
      RECT 24.405 1.962 24.41 2.179 ;
      RECT 24.4 1.972 24.405 2.163 ;
      RECT 24.39 1.98 24.4 2.132 ;
      RECT 24.385 1.99 24.39 2.106 ;
      RECT 24.38 2.047 24.385 2.089 ;
      RECT 24.485 1.925 24.61 2.43 ;
      RECT 24.2 2.612 24.46 2.91 ;
      RECT 24.195 2.619 24.46 2.908 ;
      RECT 24.2 2.614 24.475 2.903 ;
      RECT 24.19 2.627 24.475 2.9 ;
      RECT 24.19 2.632 24.48 2.893 ;
      RECT 24.185 2.64 24.48 2.89 ;
      RECT 24.185 2.657 24.485 2.688 ;
      RECT 24.2 2.609 24.431 2.91 ;
      RECT 24.255 2.608 24.431 2.91 ;
      RECT 24.255 2.605 24.345 2.91 ;
      RECT 24.255 2.602 24.341 2.91 ;
      RECT 23.945 2.875 23.95 2.888 ;
      RECT 23.94 2.842 23.945 2.893 ;
      RECT 23.935 2.797 23.94 2.9 ;
      RECT 23.93 2.752 23.935 2.908 ;
      RECT 23.925 2.72 23.93 2.916 ;
      RECT 23.92 2.68 23.925 2.917 ;
      RECT 23.905 2.66 23.92 2.919 ;
      RECT 23.83 2.642 23.905 2.931 ;
      RECT 23.82 2.635 23.83 2.942 ;
      RECT 23.815 2.635 23.82 2.944 ;
      RECT 23.785 2.641 23.815 2.948 ;
      RECT 23.745 2.654 23.785 2.948 ;
      RECT 23.72 2.665 23.745 2.934 ;
      RECT 23.705 2.671 23.72 2.917 ;
      RECT 23.695 2.673 23.705 2.908 ;
      RECT 23.69 2.674 23.695 2.903 ;
      RECT 23.685 2.675 23.69 2.898 ;
      RECT 23.68 2.676 23.685 2.895 ;
      RECT 23.655 2.681 23.68 2.885 ;
      RECT 23.645 2.697 23.655 2.872 ;
      RECT 23.64 2.717 23.645 2.867 ;
      RECT 23.65 2.11 23.655 2.306 ;
      RECT 23.635 2.074 23.65 2.308 ;
      RECT 23.625 2.056 23.635 2.313 ;
      RECT 23.615 2.042 23.625 2.317 ;
      RECT 23.57 2.026 23.615 2.327 ;
      RECT 23.565 2.016 23.57 2.336 ;
      RECT 23.52 2.005 23.565 2.342 ;
      RECT 23.515 1.993 23.52 2.349 ;
      RECT 23.5 1.988 23.515 2.353 ;
      RECT 23.485 1.98 23.5 2.358 ;
      RECT 23.475 1.973 23.485 2.363 ;
      RECT 23.465 1.97 23.475 2.368 ;
      RECT 23.455 1.97 23.465 2.369 ;
      RECT 23.45 1.967 23.455 2.368 ;
      RECT 23.415 1.962 23.44 2.367 ;
      RECT 23.391 1.958 23.415 2.366 ;
      RECT 23.305 1.949 23.391 2.363 ;
      RECT 23.29 1.941 23.305 2.36 ;
      RECT 23.268 1.94 23.29 2.359 ;
      RECT 23.182 1.94 23.268 2.357 ;
      RECT 23.096 1.94 23.182 2.355 ;
      RECT 23.01 1.94 23.096 2.352 ;
      RECT 23 1.94 23.01 2.343 ;
      RECT 22.97 1.94 23 2.303 ;
      RECT 22.96 1.95 22.97 2.258 ;
      RECT 22.955 1.99 22.96 2.243 ;
      RECT 22.95 2.005 22.955 2.23 ;
      RECT 22.92 2.085 22.95 2.192 ;
      RECT 23.44 1.965 23.45 2.368 ;
      RECT 23.265 2.73 23.28 3.335 ;
      RECT 23.27 2.725 23.28 3.335 ;
      RECT 23.435 2.725 23.44 2.908 ;
      RECT 23.425 2.725 23.435 2.938 ;
      RECT 23.41 2.725 23.425 2.998 ;
      RECT 23.405 2.725 23.41 3.043 ;
      RECT 23.4 2.725 23.405 3.073 ;
      RECT 23.395 2.725 23.4 3.093 ;
      RECT 23.385 2.725 23.395 3.128 ;
      RECT 23.37 2.725 23.385 3.16 ;
      RECT 23.325 2.725 23.37 3.188 ;
      RECT 23.32 2.725 23.325 3.218 ;
      RECT 23.315 2.725 23.32 3.23 ;
      RECT 23.31 2.725 23.315 3.238 ;
      RECT 23.3 2.725 23.31 3.253 ;
      RECT 23.295 2.725 23.3 3.275 ;
      RECT 23.285 2.725 23.295 3.298 ;
      RECT 23.28 2.725 23.285 3.318 ;
      RECT 23.245 2.74 23.265 3.335 ;
      RECT 23.22 2.757 23.245 3.335 ;
      RECT 23.215 2.767 23.22 3.335 ;
      RECT 23.185 2.782 23.215 3.335 ;
      RECT 23.11 2.824 23.185 3.335 ;
      RECT 23.105 2.855 23.11 3.318 ;
      RECT 23.1 2.859 23.105 3.3 ;
      RECT 23.095 2.863 23.1 3.263 ;
      RECT 23.09 3.047 23.095 3.23 ;
      RECT 22.575 3.236 22.661 3.801 ;
      RECT 22.53 3.238 22.695 3.795 ;
      RECT 22.661 3.235 22.695 3.795 ;
      RECT 22.575 3.237 22.78 3.789 ;
      RECT 22.53 3.247 22.79 3.785 ;
      RECT 22.505 3.239 22.78 3.781 ;
      RECT 22.5 3.242 22.78 3.776 ;
      RECT 22.475 3.257 22.79 3.77 ;
      RECT 22.475 3.282 22.83 3.765 ;
      RECT 22.435 3.29 22.83 3.74 ;
      RECT 22.435 3.317 22.845 3.738 ;
      RECT 22.435 3.347 22.855 3.725 ;
      RECT 22.43 3.492 22.855 3.713 ;
      RECT 22.435 3.421 22.875 3.71 ;
      RECT 22.435 3.478 22.88 3.518 ;
      RECT 22.625 2.757 22.795 2.935 ;
      RECT 22.575 2.696 22.625 2.92 ;
      RECT 22.31 2.676 22.575 2.905 ;
      RECT 22.27 2.74 22.745 2.905 ;
      RECT 22.27 2.73 22.7 2.905 ;
      RECT 22.27 2.727 22.69 2.905 ;
      RECT 22.27 2.715 22.68 2.905 ;
      RECT 22.27 2.7 22.625 2.905 ;
      RECT 22.31 2.672 22.511 2.905 ;
      RECT 22.32 2.65 22.511 2.905 ;
      RECT 22.345 2.635 22.425 2.905 ;
      RECT 22.1 3.165 22.22 3.61 ;
      RECT 22.085 3.165 22.22 3.609 ;
      RECT 22.04 3.187 22.22 3.604 ;
      RECT 22 3.236 22.22 3.598 ;
      RECT 22 3.236 22.225 3.573 ;
      RECT 22 3.236 22.245 3.463 ;
      RECT 21.995 3.266 22.245 3.46 ;
      RECT 22.085 3.165 22.255 3.355 ;
      RECT 21.745 1.95 21.75 2.395 ;
      RECT 21.555 1.95 21.575 2.36 ;
      RECT 21.525 1.95 21.53 2.335 ;
      RECT 22.205 2.257 22.22 2.445 ;
      RECT 22.2 2.242 22.205 2.451 ;
      RECT 22.18 2.215 22.2 2.454 ;
      RECT 22.13 2.182 22.18 2.463 ;
      RECT 22.1 2.162 22.13 2.467 ;
      RECT 22.081 2.15 22.1 2.463 ;
      RECT 21.995 2.122 22.081 2.453 ;
      RECT 21.985 2.097 21.995 2.443 ;
      RECT 21.915 2.065 21.985 2.435 ;
      RECT 21.89 2.025 21.915 2.427 ;
      RECT 21.87 2.007 21.89 2.421 ;
      RECT 21.86 1.997 21.87 2.418 ;
      RECT 21.85 1.99 21.86 2.416 ;
      RECT 21.83 1.977 21.85 2.413 ;
      RECT 21.82 1.967 21.83 2.41 ;
      RECT 21.81 1.96 21.82 2.408 ;
      RECT 21.76 1.952 21.81 2.402 ;
      RECT 21.75 1.95 21.76 2.396 ;
      RECT 21.72 1.95 21.745 2.393 ;
      RECT 21.691 1.95 21.72 2.388 ;
      RECT 21.605 1.95 21.691 2.378 ;
      RECT 21.575 1.95 21.605 2.365 ;
      RECT 21.53 1.95 21.555 2.348 ;
      RECT 21.515 1.95 21.525 2.33 ;
      RECT 21.495 1.957 21.515 2.315 ;
      RECT 21.49 1.972 21.495 2.303 ;
      RECT 21.485 1.977 21.49 2.243 ;
      RECT 21.48 1.982 21.485 2.085 ;
      RECT 21.475 1.985 21.48 2.003 ;
      RECT 21.74 2.67 21.826 2.991 ;
      RECT 21.74 2.67 21.86 2.984 ;
      RECT 21.69 2.67 21.86 2.98 ;
      RECT 21.69 2.672 21.946 2.978 ;
      RECT 21.69 2.674 21.97 2.972 ;
      RECT 21.69 2.681 21.98 2.971 ;
      RECT 21.69 2.69 21.985 2.968 ;
      RECT 21.69 2.696 21.99 2.963 ;
      RECT 21.69 2.74 21.995 2.96 ;
      RECT 21.69 2.832 22 2.957 ;
      RECT 21.215 3.275 21.25 3.595 ;
      RECT 21.8 3.46 21.805 3.642 ;
      RECT 21.755 3.342 21.8 3.661 ;
      RECT 21.74 3.319 21.755 3.684 ;
      RECT 21.73 3.309 21.74 3.694 ;
      RECT 21.71 3.304 21.73 3.707 ;
      RECT 21.685 3.302 21.71 3.728 ;
      RECT 21.666 3.301 21.685 3.74 ;
      RECT 21.58 3.298 21.666 3.74 ;
      RECT 21.51 3.293 21.58 3.728 ;
      RECT 21.435 3.289 21.51 3.703 ;
      RECT 21.37 3.285 21.435 3.67 ;
      RECT 21.3 3.282 21.37 3.63 ;
      RECT 21.27 3.278 21.3 3.605 ;
      RECT 21.25 3.276 21.27 3.598 ;
      RECT 21.166 3.274 21.215 3.596 ;
      RECT 21.08 3.271 21.166 3.597 ;
      RECT 21.005 3.27 21.08 3.599 ;
      RECT 20.92 3.27 21.005 3.625 ;
      RECT 20.843 3.271 20.92 3.65 ;
      RECT 20.757 3.272 20.843 3.65 ;
      RECT 20.671 3.272 20.757 3.65 ;
      RECT 20.585 3.273 20.671 3.65 ;
      RECT 20.565 3.274 20.585 3.642 ;
      RECT 20.55 3.28 20.565 3.627 ;
      RECT 20.515 3.3 20.55 3.607 ;
      RECT 20.505 3.32 20.515 3.589 ;
      RECT 21.475 2.625 21.48 2.895 ;
      RECT 21.47 2.616 21.475 2.9 ;
      RECT 21.46 2.606 21.47 2.912 ;
      RECT 21.455 2.595 21.46 2.923 ;
      RECT 21.435 2.589 21.455 2.941 ;
      RECT 21.39 2.586 21.435 2.99 ;
      RECT 21.375 2.585 21.39 3.035 ;
      RECT 21.37 2.585 21.375 3.048 ;
      RECT 21.36 2.585 21.37 3.06 ;
      RECT 21.355 2.586 21.36 3.075 ;
      RECT 21.335 2.594 21.355 3.08 ;
      RECT 21.305 2.61 21.335 3.08 ;
      RECT 21.295 2.622 21.3 3.08 ;
      RECT 21.26 2.637 21.295 3.08 ;
      RECT 21.23 2.657 21.26 3.08 ;
      RECT 21.22 2.682 21.23 3.08 ;
      RECT 21.215 2.71 21.22 3.08 ;
      RECT 21.21 2.74 21.215 3.08 ;
      RECT 21.205 2.757 21.21 3.08 ;
      RECT 21.195 2.785 21.205 3.08 ;
      RECT 21.185 2.82 21.195 3.08 ;
      RECT 21.18 2.855 21.185 3.08 ;
      RECT 21.3 2.62 21.305 3.08 ;
      RECT 20.815 2.722 21 2.895 ;
      RECT 20.775 2.64 20.96 2.893 ;
      RECT 20.736 2.645 20.96 2.889 ;
      RECT 20.65 2.654 20.96 2.884 ;
      RECT 20.566 2.67 20.965 2.879 ;
      RECT 20.48 2.69 20.99 2.873 ;
      RECT 20.48 2.71 20.995 2.873 ;
      RECT 20.566 2.68 20.99 2.879 ;
      RECT 20.65 2.655 20.965 2.884 ;
      RECT 20.815 2.637 20.96 2.895 ;
      RECT 20.815 2.632 20.915 2.895 ;
      RECT 20.901 2.626 20.915 2.895 ;
      RECT 20.29 1.95 20.295 2.349 ;
      RECT 20.035 1.95 20.07 2.347 ;
      RECT 19.63 1.985 19.635 2.341 ;
      RECT 20.375 1.988 20.38 2.243 ;
      RECT 20.37 1.986 20.375 2.249 ;
      RECT 20.365 1.985 20.37 2.256 ;
      RECT 20.34 1.978 20.365 2.28 ;
      RECT 20.335 1.971 20.34 2.304 ;
      RECT 20.33 1.967 20.335 2.313 ;
      RECT 20.32 1.962 20.33 2.326 ;
      RECT 20.315 1.959 20.32 2.335 ;
      RECT 20.31 1.957 20.315 2.34 ;
      RECT 20.295 1.953 20.31 2.35 ;
      RECT 20.28 1.947 20.29 2.349 ;
      RECT 20.242 1.945 20.28 2.349 ;
      RECT 20.156 1.947 20.242 2.349 ;
      RECT 20.07 1.949 20.156 2.348 ;
      RECT 19.999 1.95 20.035 2.347 ;
      RECT 19.913 1.952 19.999 2.347 ;
      RECT 19.827 1.954 19.913 2.346 ;
      RECT 19.741 1.956 19.827 2.346 ;
      RECT 19.655 1.959 19.741 2.345 ;
      RECT 19.645 1.965 19.655 2.344 ;
      RECT 19.635 1.977 19.645 2.342 ;
      RECT 19.575 2.012 19.63 2.338 ;
      RECT 19.57 2.042 19.575 2.1 ;
      RECT 20.315 3.122 20.33 3.315 ;
      RECT 20.31 3.09 20.315 3.315 ;
      RECT 20.3 3.065 20.31 3.315 ;
      RECT 20.295 3.037 20.3 3.315 ;
      RECT 20.265 2.96 20.295 3.315 ;
      RECT 20.24 2.842 20.265 3.315 ;
      RECT 20.235 2.78 20.24 3.315 ;
      RECT 20.225 2.767 20.235 3.315 ;
      RECT 20.205 2.757 20.225 3.315 ;
      RECT 20.19 2.74 20.205 3.315 ;
      RECT 20.16 2.728 20.19 3.315 ;
      RECT 20.155 2.727 20.16 3.26 ;
      RECT 20.15 2.727 20.155 3.218 ;
      RECT 20.135 2.726 20.15 3.17 ;
      RECT 20.12 2.726 20.135 3.108 ;
      RECT 20.1 2.726 20.12 3.068 ;
      RECT 20.095 2.726 20.1 3.053 ;
      RECT 20.07 2.725 20.095 3.048 ;
      RECT 20 2.724 20.07 3.035 ;
      RECT 19.985 2.723 20 3.02 ;
      RECT 19.955 2.722 19.985 3.003 ;
      RECT 19.95 2.722 19.955 2.988 ;
      RECT 19.9 2.721 19.95 2.968 ;
      RECT 19.835 2.72 19.9 2.923 ;
      RECT 19.83 2.72 19.835 2.895 ;
      RECT 19.915 3.257 19.92 3.514 ;
      RECT 19.895 3.176 19.915 3.531 ;
      RECT 19.875 3.17 19.895 3.56 ;
      RECT 19.815 3.157 19.875 3.58 ;
      RECT 19.77 3.141 19.815 3.581 ;
      RECT 19.686 3.129 19.77 3.569 ;
      RECT 19.6 3.116 19.686 3.553 ;
      RECT 19.59 3.109 19.6 3.545 ;
      RECT 19.545 3.106 19.59 3.485 ;
      RECT 19.525 3.102 19.545 3.4 ;
      RECT 19.51 3.1 19.525 3.353 ;
      RECT 19.48 3.097 19.51 3.323 ;
      RECT 19.445 3.093 19.48 3.3 ;
      RECT 19.402 3.088 19.445 3.288 ;
      RECT 19.316 3.079 19.402 3.297 ;
      RECT 19.23 3.068 19.316 3.309 ;
      RECT 19.165 3.059 19.23 3.318 ;
      RECT 19.145 3.05 19.165 3.323 ;
      RECT 19.14 3.043 19.145 3.325 ;
      RECT 19.1 3.028 19.14 3.322 ;
      RECT 19.08 3.007 19.1 3.317 ;
      RECT 19.065 2.995 19.08 3.31 ;
      RECT 19.06 2.987 19.065 3.303 ;
      RECT 19.045 2.967 19.06 3.296 ;
      RECT 19.04 2.83 19.045 3.29 ;
      RECT 18.96 2.719 19.04 3.262 ;
      RECT 18.951 2.712 18.96 3.228 ;
      RECT 18.865 2.706 18.951 3.153 ;
      RECT 18.84 2.697 18.865 3.065 ;
      RECT 18.81 2.692 18.84 3.04 ;
      RECT 18.745 2.701 18.81 3.025 ;
      RECT 18.725 2.717 18.745 3 ;
      RECT 18.715 2.723 18.725 2.948 ;
      RECT 18.695 2.745 18.715 2.83 ;
      RECT 19.35 2.71 19.52 2.895 ;
      RECT 19.35 2.71 19.555 2.893 ;
      RECT 19.4 2.62 19.57 2.884 ;
      RECT 19.35 2.777 19.575 2.877 ;
      RECT 19.365 2.655 19.57 2.884 ;
      RECT 18.565 3.388 18.63 3.831 ;
      RECT 18.505 3.413 18.63 3.829 ;
      RECT 18.505 3.413 18.685 3.823 ;
      RECT 18.49 3.438 18.685 3.822 ;
      RECT 18.63 3.375 18.705 3.819 ;
      RECT 18.565 3.4 18.785 3.813 ;
      RECT 18.49 3.439 18.83 3.807 ;
      RECT 18.475 3.466 18.83 3.798 ;
      RECT 18.49 3.459 18.85 3.79 ;
      RECT 18.475 3.468 18.855 3.773 ;
      RECT 18.47 3.485 18.855 3.6 ;
      RECT 18.475 2.207 18.51 2.445 ;
      RECT 18.475 2.207 18.54 2.444 ;
      RECT 18.475 2.207 18.655 2.44 ;
      RECT 18.475 2.207 18.71 2.418 ;
      RECT 18.485 2.15 18.765 2.318 ;
      RECT 18.59 1.99 18.62 2.441 ;
      RECT 18.62 1.985 18.8 2.198 ;
      RECT 18.49 2.126 18.8 2.198 ;
      RECT 18.54 2.022 18.59 2.442 ;
      RECT 18.51 2.078 18.8 2.198 ;
      RECT 17.02 1.74 17.19 2.935 ;
      RECT 17.02 1.74 17.485 1.91 ;
      RECT 17.02 6.97 17.485 7.14 ;
      RECT 17.02 5.945 17.19 7.14 ;
      RECT 16.03 1.74 16.2 2.935 ;
      RECT 16.03 1.74 16.495 1.91 ;
      RECT 16.03 6.97 16.495 7.14 ;
      RECT 16.03 5.945 16.2 7.14 ;
      RECT 14.175 2.635 14.345 3.865 ;
      RECT 14.23 0.855 14.4 2.805 ;
      RECT 14.175 0.575 14.345 1.025 ;
      RECT 14.175 7.855 14.345 8.305 ;
      RECT 14.23 6.075 14.4 8.025 ;
      RECT 14.175 5.015 14.345 6.245 ;
      RECT 13.655 0.575 13.825 3.865 ;
      RECT 13.655 2.075 14.06 2.405 ;
      RECT 13.655 1.235 14.06 1.565 ;
      RECT 13.655 5.015 13.825 8.305 ;
      RECT 13.655 7.315 14.06 7.645 ;
      RECT 13.655 6.475 14.06 6.805 ;
      RECT 11.755 3.392 11.77 3.443 ;
      RECT 11.75 3.372 11.755 3.49 ;
      RECT 11.735 3.362 11.75 3.558 ;
      RECT 11.71 3.342 11.735 3.613 ;
      RECT 11.67 3.327 11.71 3.633 ;
      RECT 11.625 3.321 11.67 3.661 ;
      RECT 11.555 3.311 11.625 3.678 ;
      RECT 11.535 3.303 11.555 3.678 ;
      RECT 11.475 3.297 11.535 3.67 ;
      RECT 11.416 3.288 11.475 3.658 ;
      RECT 11.33 3.277 11.416 3.641 ;
      RECT 11.308 3.268 11.33 3.629 ;
      RECT 11.222 3.261 11.308 3.616 ;
      RECT 11.136 3.248 11.222 3.597 ;
      RECT 11.05 3.236 11.136 3.577 ;
      RECT 11.02 3.225 11.05 3.564 ;
      RECT 10.97 3.211 11.02 3.556 ;
      RECT 10.95 3.2 10.97 3.548 ;
      RECT 10.901 3.189 10.95 3.54 ;
      RECT 10.815 3.168 10.901 3.525 ;
      RECT 10.77 3.155 10.815 3.51 ;
      RECT 10.725 3.155 10.77 3.49 ;
      RECT 10.67 3.155 10.725 3.425 ;
      RECT 10.645 3.155 10.67 3.348 ;
      RECT 11.17 2.892 11.34 3.075 ;
      RECT 11.17 2.892 11.355 3.033 ;
      RECT 11.17 2.892 11.36 2.975 ;
      RECT 11.23 2.66 11.365 2.951 ;
      RECT 11.23 2.664 11.37 2.934 ;
      RECT 11.175 2.827 11.37 2.934 ;
      RECT 11.2 2.672 11.34 3.075 ;
      RECT 11.2 2.676 11.38 2.875 ;
      RECT 11.185 2.762 11.38 2.875 ;
      RECT 11.195 2.692 11.34 3.075 ;
      RECT 11.195 2.695 11.39 2.788 ;
      RECT 11.19 2.712 11.39 2.788 ;
      RECT 10.96 1.932 11.13 2.415 ;
      RECT 10.955 1.927 11.105 2.405 ;
      RECT 10.955 1.934 11.135 2.399 ;
      RECT 10.945 1.928 11.105 2.378 ;
      RECT 10.945 1.944 11.15 2.337 ;
      RECT 10.915 1.929 11.105 2.3 ;
      RECT 10.915 1.959 11.16 2.24 ;
      RECT 10.91 1.931 11.105 2.238 ;
      RECT 10.89 1.94 11.135 2.195 ;
      RECT 10.865 1.956 11.15 2.107 ;
      RECT 10.865 1.975 11.175 2.098 ;
      RECT 10.86 2.012 11.175 2.05 ;
      RECT 10.865 1.992 11.18 2.018 ;
      RECT 10.96 1.926 11.07 2.415 ;
      RECT 11.046 1.925 11.07 2.415 ;
      RECT 10.28 2.71 10.285 2.921 ;
      RECT 10.88 2.71 10.885 2.895 ;
      RECT 10.945 2.75 10.95 2.863 ;
      RECT 10.94 2.742 10.945 2.869 ;
      RECT 10.935 2.732 10.94 2.877 ;
      RECT 10.93 2.722 10.935 2.886 ;
      RECT 10.925 2.712 10.93 2.89 ;
      RECT 10.885 2.71 10.925 2.893 ;
      RECT 10.857 2.709 10.88 2.897 ;
      RECT 10.771 2.706 10.857 2.904 ;
      RECT 10.685 2.702 10.771 2.915 ;
      RECT 10.665 2.7 10.685 2.921 ;
      RECT 10.647 2.699 10.665 2.924 ;
      RECT 10.561 2.697 10.647 2.931 ;
      RECT 10.475 2.692 10.561 2.944 ;
      RECT 10.456 2.689 10.475 2.949 ;
      RECT 10.37 2.687 10.456 2.94 ;
      RECT 10.36 2.687 10.37 2.933 ;
      RECT 10.285 2.7 10.36 2.927 ;
      RECT 10.27 2.711 10.28 2.921 ;
      RECT 10.26 2.713 10.27 2.92 ;
      RECT 10.25 2.717 10.26 2.916 ;
      RECT 10.245 2.72 10.25 2.91 ;
      RECT 10.235 2.722 10.245 2.904 ;
      RECT 10.23 2.725 10.235 2.898 ;
      RECT 10.21 3.311 10.215 3.515 ;
      RECT 10.195 3.298 10.21 3.608 ;
      RECT 10.18 3.279 10.195 3.885 ;
      RECT 10.145 3.245 10.18 3.885 ;
      RECT 10.141 3.215 10.145 3.885 ;
      RECT 10.055 3.097 10.141 3.885 ;
      RECT 10.045 2.972 10.055 3.885 ;
      RECT 10.03 2.94 10.045 3.885 ;
      RECT 10.025 2.915 10.03 3.885 ;
      RECT 10.02 2.905 10.025 3.841 ;
      RECT 10.005 2.877 10.02 3.746 ;
      RECT 9.99 2.843 10.005 3.645 ;
      RECT 9.985 2.821 9.99 3.598 ;
      RECT 9.98 2.81 9.985 3.568 ;
      RECT 9.975 2.8 9.98 3.534 ;
      RECT 9.965 2.787 9.975 3.502 ;
      RECT 9.94 2.763 9.965 3.428 ;
      RECT 9.935 2.743 9.94 3.353 ;
      RECT 9.93 2.737 9.935 3.328 ;
      RECT 9.925 2.732 9.93 3.293 ;
      RECT 9.92 2.727 9.925 3.268 ;
      RECT 9.915 2.725 9.92 3.248 ;
      RECT 9.91 2.725 9.915 3.233 ;
      RECT 9.905 2.725 9.91 3.193 ;
      RECT 9.895 2.725 9.905 3.165 ;
      RECT 9.885 2.725 9.895 3.11 ;
      RECT 9.87 2.725 9.885 3.048 ;
      RECT 9.865 2.724 9.87 2.993 ;
      RECT 9.85 2.723 9.865 2.973 ;
      RECT 9.79 2.721 9.85 2.947 ;
      RECT 9.755 2.722 9.79 2.927 ;
      RECT 9.75 2.724 9.755 2.917 ;
      RECT 9.74 2.743 9.75 2.907 ;
      RECT 9.735 2.77 9.74 2.838 ;
      RECT 9.85 2.195 10.02 2.44 ;
      RECT 9.885 1.966 10.02 2.44 ;
      RECT 9.885 1.968 10.03 2.435 ;
      RECT 9.885 1.97 10.055 2.423 ;
      RECT 9.885 1.973 10.08 2.405 ;
      RECT 9.885 1.978 10.13 2.378 ;
      RECT 9.885 1.983 10.15 2.343 ;
      RECT 9.865 1.985 10.16 2.318 ;
      RECT 9.855 2.08 10.16 2.318 ;
      RECT 9.885 1.965 9.995 2.44 ;
      RECT 9.895 1.962 9.99 2.44 ;
      RECT 9.415 3.227 9.605 3.585 ;
      RECT 9.415 3.239 9.64 3.584 ;
      RECT 9.415 3.267 9.66 3.582 ;
      RECT 9.415 3.292 9.665 3.581 ;
      RECT 9.415 3.35 9.68 3.58 ;
      RECT 9.4 3.223 9.56 3.565 ;
      RECT 9.38 3.232 9.605 3.518 ;
      RECT 9.355 3.243 9.64 3.455 ;
      RECT 9.355 3.327 9.675 3.455 ;
      RECT 9.355 3.302 9.67 3.455 ;
      RECT 9.415 3.218 9.56 3.585 ;
      RECT 9.501 3.217 9.56 3.585 ;
      RECT 9.501 3.216 9.545 3.585 ;
      RECT 9.2 2.732 9.205 3.11 ;
      RECT 9.195 2.7 9.2 3.11 ;
      RECT 9.19 2.672 9.195 3.11 ;
      RECT 9.185 2.652 9.19 3.11 ;
      RECT 9.13 2.635 9.185 3.11 ;
      RECT 9.09 2.62 9.13 3.11 ;
      RECT 9.035 2.607 9.09 3.11 ;
      RECT 9 2.598 9.035 3.11 ;
      RECT 8.996 2.596 9 3.109 ;
      RECT 8.91 2.592 8.996 3.092 ;
      RECT 8.825 2.584 8.91 3.055 ;
      RECT 8.815 2.58 8.825 3.028 ;
      RECT 8.805 2.58 8.815 3.01 ;
      RECT 8.795 2.582 8.805 2.993 ;
      RECT 8.79 2.587 8.795 2.979 ;
      RECT 8.785 2.591 8.79 2.966 ;
      RECT 8.775 2.596 8.785 2.95 ;
      RECT 8.76 2.61 8.775 2.925 ;
      RECT 8.755 2.616 8.76 2.905 ;
      RECT 8.75 2.618 8.755 2.898 ;
      RECT 8.745 2.622 8.75 2.773 ;
      RECT 8.925 3.422 9.17 3.885 ;
      RECT 8.845 3.395 9.165 3.881 ;
      RECT 8.775 3.43 9.17 3.874 ;
      RECT 8.565 3.685 9.17 3.87 ;
      RECT 8.745 3.453 9.17 3.87 ;
      RECT 8.585 3.645 9.17 3.87 ;
      RECT 8.735 3.465 9.17 3.87 ;
      RECT 8.62 3.582 9.17 3.87 ;
      RECT 8.675 3.507 9.17 3.87 ;
      RECT 8.925 3.372 9.165 3.885 ;
      RECT 8.955 3.365 9.165 3.885 ;
      RECT 8.945 3.367 9.165 3.885 ;
      RECT 8.955 3.362 9.085 3.885 ;
      RECT 8.51 1.925 8.596 2.364 ;
      RECT 8.505 1.925 8.596 2.362 ;
      RECT 8.505 1.925 8.665 2.361 ;
      RECT 8.505 1.925 8.695 2.358 ;
      RECT 8.49 1.932 8.695 2.349 ;
      RECT 8.49 1.932 8.7 2.345 ;
      RECT 8.485 1.942 8.7 2.338 ;
      RECT 8.48 1.947 8.7 2.313 ;
      RECT 8.48 1.947 8.715 2.295 ;
      RECT 8.505 1.925 8.735 2.21 ;
      RECT 8.475 1.952 8.735 2.208 ;
      RECT 8.485 1.945 8.74 2.146 ;
      RECT 8.475 2.067 8.745 2.129 ;
      RECT 8.46 1.962 8.74 2.08 ;
      RECT 8.455 1.972 8.74 1.98 ;
      RECT 8.535 2.743 8.54 2.82 ;
      RECT 8.525 2.737 8.535 3.01 ;
      RECT 8.515 2.729 8.525 3.031 ;
      RECT 8.505 2.72 8.515 3.053 ;
      RECT 8.5 2.715 8.505 3.07 ;
      RECT 8.46 2.715 8.5 3.11 ;
      RECT 8.44 2.715 8.46 3.165 ;
      RECT 8.435 2.715 8.44 3.193 ;
      RECT 8.425 2.715 8.435 3.208 ;
      RECT 8.39 2.715 8.425 3.25 ;
      RECT 8.385 2.715 8.39 3.293 ;
      RECT 8.375 2.715 8.385 3.308 ;
      RECT 8.36 2.715 8.375 3.328 ;
      RECT 8.345 2.715 8.36 3.355 ;
      RECT 8.34 2.716 8.345 3.373 ;
      RECT 8.32 2.717 8.34 3.38 ;
      RECT 8.265 2.718 8.32 3.4 ;
      RECT 8.255 2.719 8.265 3.414 ;
      RECT 8.25 2.722 8.255 3.413 ;
      RECT 8.21 2.795 8.25 3.411 ;
      RECT 8.195 2.875 8.21 3.409 ;
      RECT 8.17 2.93 8.195 3.407 ;
      RECT 8.155 2.995 8.17 3.406 ;
      RECT 8.11 3.027 8.155 3.403 ;
      RECT 8.025 3.05 8.11 3.398 ;
      RECT 8 3.07 8.025 3.393 ;
      RECT 7.93 3.075 8 3.389 ;
      RECT 7.91 3.077 7.93 3.386 ;
      RECT 7.825 3.088 7.91 3.38 ;
      RECT 7.82 3.099 7.825 3.375 ;
      RECT 7.81 3.101 7.82 3.375 ;
      RECT 7.775 3.105 7.81 3.373 ;
      RECT 7.725 3.115 7.775 3.36 ;
      RECT 7.705 3.123 7.725 3.345 ;
      RECT 7.625 3.135 7.705 3.328 ;
      RECT 7.79 2.685 7.96 2.895 ;
      RECT 7.906 2.681 7.96 2.895 ;
      RECT 7.711 2.685 7.96 2.886 ;
      RECT 7.711 2.685 7.965 2.875 ;
      RECT 7.625 2.685 7.965 2.866 ;
      RECT 7.625 2.693 7.975 2.81 ;
      RECT 7.625 2.705 7.98 2.723 ;
      RECT 7.625 2.712 7.985 2.715 ;
      RECT 7.82 2.683 7.96 2.895 ;
      RECT 7.575 3.628 7.82 3.96 ;
      RECT 7.57 3.62 7.575 3.957 ;
      RECT 7.54 3.64 7.82 3.938 ;
      RECT 7.52 3.672 7.82 3.911 ;
      RECT 7.57 3.625 7.747 3.957 ;
      RECT 7.57 3.622 7.661 3.957 ;
      RECT 7.51 1.97 7.68 2.39 ;
      RECT 7.505 1.97 7.68 2.388 ;
      RECT 7.505 1.97 7.705 2.378 ;
      RECT 7.505 1.97 7.725 2.353 ;
      RECT 7.5 1.97 7.725 2.348 ;
      RECT 7.5 1.97 7.735 2.338 ;
      RECT 7.5 1.97 7.74 2.333 ;
      RECT 7.5 1.975 7.745 2.328 ;
      RECT 7.5 2.007 7.76 2.318 ;
      RECT 7.5 2.077 7.785 2.301 ;
      RECT 7.48 2.077 7.785 2.293 ;
      RECT 7.48 2.137 7.795 2.27 ;
      RECT 7.48 2.177 7.805 2.215 ;
      RECT 7.465 1.97 7.74 2.195 ;
      RECT 7.455 1.985 7.745 2.093 ;
      RECT 7.045 3.375 7.215 3.9 ;
      RECT 7.04 3.375 7.215 3.893 ;
      RECT 7.03 3.375 7.22 3.858 ;
      RECT 7.025 3.385 7.22 3.83 ;
      RECT 7.02 3.405 7.22 3.813 ;
      RECT 7.03 3.38 7.225 3.803 ;
      RECT 7.015 3.425 7.225 3.795 ;
      RECT 7.01 3.445 7.225 3.78 ;
      RECT 7.005 3.475 7.225 3.77 ;
      RECT 6.995 3.52 7.225 3.745 ;
      RECT 7.025 3.39 7.23 3.728 ;
      RECT 6.99 3.572 7.23 3.723 ;
      RECT 7.025 3.4 7.235 3.693 ;
      RECT 6.985 3.605 7.235 3.69 ;
      RECT 6.98 3.63 7.235 3.67 ;
      RECT 7.02 3.417 7.245 3.61 ;
      RECT 7.015 3.439 7.255 3.503 ;
      RECT 6.965 2.686 6.98 2.955 ;
      RECT 6.92 2.67 6.965 3 ;
      RECT 6.915 2.658 6.92 3.05 ;
      RECT 6.905 2.654 6.915 3.083 ;
      RECT 6.9 2.651 6.905 3.111 ;
      RECT 6.885 2.653 6.9 3.153 ;
      RECT 6.88 2.657 6.885 3.193 ;
      RECT 6.86 2.662 6.88 3.245 ;
      RECT 6.856 2.667 6.86 3.302 ;
      RECT 6.77 2.686 6.856 3.339 ;
      RECT 6.76 2.707 6.77 3.375 ;
      RECT 6.755 2.715 6.76 3.376 ;
      RECT 6.75 2.757 6.755 3.377 ;
      RECT 6.735 2.845 6.75 3.378 ;
      RECT 6.725 2.995 6.735 3.38 ;
      RECT 6.72 3.04 6.725 3.382 ;
      RECT 6.685 3.082 6.72 3.385 ;
      RECT 6.68 3.1 6.685 3.388 ;
      RECT 6.603 3.106 6.68 3.394 ;
      RECT 6.517 3.12 6.603 3.407 ;
      RECT 6.431 3.134 6.517 3.421 ;
      RECT 6.345 3.148 6.431 3.434 ;
      RECT 6.285 3.16 6.345 3.446 ;
      RECT 6.26 3.167 6.285 3.453 ;
      RECT 6.246 3.17 6.26 3.458 ;
      RECT 6.16 3.178 6.246 3.474 ;
      RECT 6.155 3.185 6.16 3.489 ;
      RECT 6.131 3.185 6.155 3.496 ;
      RECT 6.045 3.188 6.131 3.524 ;
      RECT 5.96 3.192 6.045 3.568 ;
      RECT 5.895 3.196 5.96 3.605 ;
      RECT 5.87 3.199 5.895 3.621 ;
      RECT 5.795 3.212 5.87 3.625 ;
      RECT 5.77 3.23 5.795 3.629 ;
      RECT 5.76 3.237 5.77 3.631 ;
      RECT 5.745 3.24 5.76 3.632 ;
      RECT 5.685 3.252 5.745 3.636 ;
      RECT 5.675 3.266 5.685 3.64 ;
      RECT 5.62 3.276 5.675 3.628 ;
      RECT 5.595 3.297 5.62 3.611 ;
      RECT 5.575 3.317 5.595 3.602 ;
      RECT 5.57 3.33 5.575 3.597 ;
      RECT 5.555 3.342 5.57 3.593 ;
      RECT 6.79 1.997 6.795 2.02 ;
      RECT 6.785 1.988 6.79 2.06 ;
      RECT 6.78 1.986 6.785 2.103 ;
      RECT 6.775 1.977 6.78 2.138 ;
      RECT 6.77 1.967 6.775 2.21 ;
      RECT 6.765 1.957 6.77 2.275 ;
      RECT 6.76 1.954 6.765 2.315 ;
      RECT 6.735 1.948 6.76 2.405 ;
      RECT 6.7 1.936 6.735 2.43 ;
      RECT 6.69 1.927 6.7 2.43 ;
      RECT 6.555 1.925 6.565 2.413 ;
      RECT 6.545 1.925 6.555 2.38 ;
      RECT 6.54 1.925 6.545 2.355 ;
      RECT 6.535 1.925 6.54 2.343 ;
      RECT 6.53 1.925 6.535 2.325 ;
      RECT 6.52 1.925 6.53 2.29 ;
      RECT 6.515 1.927 6.52 2.268 ;
      RECT 6.51 1.933 6.515 2.253 ;
      RECT 6.505 1.939 6.51 2.238 ;
      RECT 6.49 1.951 6.505 2.211 ;
      RECT 6.485 1.962 6.49 2.179 ;
      RECT 6.48 1.972 6.485 2.163 ;
      RECT 6.47 1.98 6.48 2.132 ;
      RECT 6.465 1.99 6.47 2.106 ;
      RECT 6.46 2.047 6.465 2.089 ;
      RECT 6.565 1.925 6.69 2.43 ;
      RECT 6.28 2.612 6.54 2.91 ;
      RECT 6.275 2.619 6.54 2.908 ;
      RECT 6.28 2.614 6.555 2.903 ;
      RECT 6.27 2.627 6.555 2.9 ;
      RECT 6.27 2.632 6.56 2.893 ;
      RECT 6.265 2.64 6.56 2.89 ;
      RECT 6.265 2.657 6.565 2.688 ;
      RECT 6.28 2.609 6.511 2.91 ;
      RECT 6.335 2.608 6.511 2.91 ;
      RECT 6.335 2.605 6.425 2.91 ;
      RECT 6.335 2.602 6.421 2.91 ;
      RECT 6.025 2.875 6.03 2.888 ;
      RECT 6.02 2.842 6.025 2.893 ;
      RECT 6.015 2.797 6.02 2.9 ;
      RECT 6.01 2.752 6.015 2.908 ;
      RECT 6.005 2.72 6.01 2.916 ;
      RECT 6 2.68 6.005 2.917 ;
      RECT 5.985 2.66 6 2.919 ;
      RECT 5.91 2.642 5.985 2.931 ;
      RECT 5.9 2.635 5.91 2.942 ;
      RECT 5.895 2.635 5.9 2.944 ;
      RECT 5.865 2.641 5.895 2.948 ;
      RECT 5.825 2.654 5.865 2.948 ;
      RECT 5.8 2.665 5.825 2.934 ;
      RECT 5.785 2.671 5.8 2.917 ;
      RECT 5.775 2.673 5.785 2.908 ;
      RECT 5.77 2.674 5.775 2.903 ;
      RECT 5.765 2.675 5.77 2.898 ;
      RECT 5.76 2.676 5.765 2.895 ;
      RECT 5.735 2.681 5.76 2.885 ;
      RECT 5.725 2.697 5.735 2.872 ;
      RECT 5.72 2.717 5.725 2.867 ;
      RECT 5.73 2.11 5.735 2.306 ;
      RECT 5.715 2.074 5.73 2.308 ;
      RECT 5.705 2.056 5.715 2.313 ;
      RECT 5.695 2.042 5.705 2.317 ;
      RECT 5.65 2.026 5.695 2.327 ;
      RECT 5.645 2.016 5.65 2.336 ;
      RECT 5.6 2.005 5.645 2.342 ;
      RECT 5.595 1.993 5.6 2.349 ;
      RECT 5.58 1.988 5.595 2.353 ;
      RECT 5.565 1.98 5.58 2.358 ;
      RECT 5.555 1.973 5.565 2.363 ;
      RECT 5.545 1.97 5.555 2.368 ;
      RECT 5.535 1.97 5.545 2.369 ;
      RECT 5.53 1.967 5.535 2.368 ;
      RECT 5.495 1.962 5.52 2.367 ;
      RECT 5.471 1.958 5.495 2.366 ;
      RECT 5.385 1.949 5.471 2.363 ;
      RECT 5.37 1.941 5.385 2.36 ;
      RECT 5.348 1.94 5.37 2.359 ;
      RECT 5.262 1.94 5.348 2.357 ;
      RECT 5.176 1.94 5.262 2.355 ;
      RECT 5.09 1.94 5.176 2.352 ;
      RECT 5.08 1.94 5.09 2.343 ;
      RECT 5.05 1.94 5.08 2.303 ;
      RECT 5.04 1.95 5.05 2.258 ;
      RECT 5.035 1.99 5.04 2.243 ;
      RECT 5.03 2.005 5.035 2.23 ;
      RECT 5 2.085 5.03 2.192 ;
      RECT 5.52 1.965 5.53 2.368 ;
      RECT 5.345 2.73 5.36 3.335 ;
      RECT 5.35 2.725 5.36 3.335 ;
      RECT 5.515 2.725 5.52 2.908 ;
      RECT 5.505 2.725 5.515 2.938 ;
      RECT 5.49 2.725 5.505 2.998 ;
      RECT 5.485 2.725 5.49 3.043 ;
      RECT 5.48 2.725 5.485 3.073 ;
      RECT 5.475 2.725 5.48 3.093 ;
      RECT 5.465 2.725 5.475 3.128 ;
      RECT 5.45 2.725 5.465 3.16 ;
      RECT 5.405 2.725 5.45 3.188 ;
      RECT 5.4 2.725 5.405 3.218 ;
      RECT 5.395 2.725 5.4 3.23 ;
      RECT 5.39 2.725 5.395 3.238 ;
      RECT 5.38 2.725 5.39 3.253 ;
      RECT 5.375 2.725 5.38 3.275 ;
      RECT 5.365 2.725 5.375 3.298 ;
      RECT 5.36 2.725 5.365 3.318 ;
      RECT 5.325 2.74 5.345 3.335 ;
      RECT 5.3 2.757 5.325 3.335 ;
      RECT 5.295 2.767 5.3 3.335 ;
      RECT 5.265 2.782 5.295 3.335 ;
      RECT 5.19 2.824 5.265 3.335 ;
      RECT 5.185 2.855 5.19 3.318 ;
      RECT 5.18 2.859 5.185 3.3 ;
      RECT 5.175 2.863 5.18 3.263 ;
      RECT 5.17 3.047 5.175 3.23 ;
      RECT 4.655 3.236 4.741 3.801 ;
      RECT 4.61 3.238 4.775 3.795 ;
      RECT 4.741 3.235 4.775 3.795 ;
      RECT 4.655 3.237 4.86 3.789 ;
      RECT 4.61 3.247 4.87 3.785 ;
      RECT 4.585 3.239 4.86 3.781 ;
      RECT 4.58 3.242 4.86 3.776 ;
      RECT 4.555 3.257 4.87 3.77 ;
      RECT 4.555 3.282 4.91 3.765 ;
      RECT 4.515 3.29 4.91 3.74 ;
      RECT 4.515 3.317 4.925 3.738 ;
      RECT 4.515 3.347 4.935 3.725 ;
      RECT 4.51 3.492 4.935 3.713 ;
      RECT 4.515 3.421 4.955 3.71 ;
      RECT 4.515 3.478 4.96 3.518 ;
      RECT 4.705 2.757 4.875 2.935 ;
      RECT 4.655 2.696 4.705 2.92 ;
      RECT 4.39 2.676 4.655 2.905 ;
      RECT 4.35 2.74 4.825 2.905 ;
      RECT 4.35 2.73 4.78 2.905 ;
      RECT 4.35 2.727 4.77 2.905 ;
      RECT 4.35 2.715 4.76 2.905 ;
      RECT 4.35 2.7 4.705 2.905 ;
      RECT 4.39 2.672 4.591 2.905 ;
      RECT 4.4 2.65 4.591 2.905 ;
      RECT 4.425 2.635 4.505 2.905 ;
      RECT 4.18 3.165 4.3 3.61 ;
      RECT 4.165 3.165 4.3 3.609 ;
      RECT 4.12 3.187 4.3 3.604 ;
      RECT 4.08 3.236 4.3 3.598 ;
      RECT 4.08 3.236 4.305 3.573 ;
      RECT 4.08 3.236 4.325 3.463 ;
      RECT 4.075 3.266 4.325 3.46 ;
      RECT 4.165 3.165 4.335 3.355 ;
      RECT 3.825 1.95 3.83 2.395 ;
      RECT 3.635 1.95 3.655 2.36 ;
      RECT 3.605 1.95 3.61 2.335 ;
      RECT 4.285 2.257 4.3 2.445 ;
      RECT 4.28 2.242 4.285 2.451 ;
      RECT 4.26 2.215 4.28 2.454 ;
      RECT 4.21 2.182 4.26 2.463 ;
      RECT 4.18 2.162 4.21 2.467 ;
      RECT 4.161 2.15 4.18 2.463 ;
      RECT 4.075 2.122 4.161 2.453 ;
      RECT 4.065 2.097 4.075 2.443 ;
      RECT 3.995 2.065 4.065 2.435 ;
      RECT 3.97 2.025 3.995 2.427 ;
      RECT 3.95 2.007 3.97 2.421 ;
      RECT 3.94 1.997 3.95 2.418 ;
      RECT 3.93 1.99 3.94 2.416 ;
      RECT 3.91 1.977 3.93 2.413 ;
      RECT 3.9 1.967 3.91 2.41 ;
      RECT 3.89 1.96 3.9 2.408 ;
      RECT 3.84 1.952 3.89 2.402 ;
      RECT 3.83 1.95 3.84 2.396 ;
      RECT 3.8 1.95 3.825 2.393 ;
      RECT 3.771 1.95 3.8 2.388 ;
      RECT 3.685 1.95 3.771 2.378 ;
      RECT 3.655 1.95 3.685 2.365 ;
      RECT 3.61 1.95 3.635 2.348 ;
      RECT 3.595 1.95 3.605 2.33 ;
      RECT 3.575 1.957 3.595 2.315 ;
      RECT 3.57 1.972 3.575 2.303 ;
      RECT 3.565 1.977 3.57 2.243 ;
      RECT 3.56 1.982 3.565 2.085 ;
      RECT 3.555 1.985 3.56 2.003 ;
      RECT 3.82 2.67 3.906 2.991 ;
      RECT 3.82 2.67 3.94 2.984 ;
      RECT 3.77 2.67 3.94 2.98 ;
      RECT 3.77 2.672 4.026 2.978 ;
      RECT 3.77 2.674 4.05 2.972 ;
      RECT 3.77 2.681 4.06 2.971 ;
      RECT 3.77 2.69 4.065 2.968 ;
      RECT 3.77 2.696 4.07 2.963 ;
      RECT 3.77 2.74 4.075 2.96 ;
      RECT 3.77 2.832 4.08 2.957 ;
      RECT 3.295 3.275 3.33 3.595 ;
      RECT 3.88 3.46 3.885 3.642 ;
      RECT 3.835 3.342 3.88 3.661 ;
      RECT 3.82 3.319 3.835 3.684 ;
      RECT 3.81 3.309 3.82 3.694 ;
      RECT 3.79 3.304 3.81 3.707 ;
      RECT 3.765 3.302 3.79 3.728 ;
      RECT 3.746 3.301 3.765 3.74 ;
      RECT 3.66 3.298 3.746 3.74 ;
      RECT 3.59 3.293 3.66 3.728 ;
      RECT 3.515 3.289 3.59 3.703 ;
      RECT 3.45 3.285 3.515 3.67 ;
      RECT 3.38 3.282 3.45 3.63 ;
      RECT 3.35 3.278 3.38 3.605 ;
      RECT 3.33 3.276 3.35 3.598 ;
      RECT 3.246 3.274 3.295 3.596 ;
      RECT 3.16 3.271 3.246 3.597 ;
      RECT 3.085 3.27 3.16 3.599 ;
      RECT 3 3.27 3.085 3.625 ;
      RECT 2.923 3.271 3 3.65 ;
      RECT 2.837 3.272 2.923 3.65 ;
      RECT 2.751 3.272 2.837 3.65 ;
      RECT 2.665 3.273 2.751 3.65 ;
      RECT 2.645 3.274 2.665 3.642 ;
      RECT 2.63 3.28 2.645 3.627 ;
      RECT 2.595 3.3 2.63 3.607 ;
      RECT 2.585 3.32 2.595 3.589 ;
      RECT 3.555 2.625 3.56 2.895 ;
      RECT 3.55 2.616 3.555 2.9 ;
      RECT 3.54 2.606 3.55 2.912 ;
      RECT 3.535 2.595 3.54 2.923 ;
      RECT 3.515 2.589 3.535 2.941 ;
      RECT 3.47 2.586 3.515 2.99 ;
      RECT 3.455 2.585 3.47 3.035 ;
      RECT 3.45 2.585 3.455 3.048 ;
      RECT 3.44 2.585 3.45 3.06 ;
      RECT 3.435 2.586 3.44 3.075 ;
      RECT 3.415 2.594 3.435 3.08 ;
      RECT 3.385 2.61 3.415 3.08 ;
      RECT 3.375 2.622 3.38 3.08 ;
      RECT 3.34 2.637 3.375 3.08 ;
      RECT 3.31 2.657 3.34 3.08 ;
      RECT 3.3 2.682 3.31 3.08 ;
      RECT 3.295 2.71 3.3 3.08 ;
      RECT 3.29 2.74 3.295 3.08 ;
      RECT 3.285 2.757 3.29 3.08 ;
      RECT 3.275 2.785 3.285 3.08 ;
      RECT 3.265 2.82 3.275 3.08 ;
      RECT 3.26 2.855 3.265 3.08 ;
      RECT 3.38 2.62 3.385 3.08 ;
      RECT 2.895 2.722 3.08 2.895 ;
      RECT 2.855 2.64 3.04 2.893 ;
      RECT 2.816 2.645 3.04 2.889 ;
      RECT 2.73 2.654 3.04 2.884 ;
      RECT 2.646 2.67 3.045 2.879 ;
      RECT 2.56 2.69 3.07 2.873 ;
      RECT 2.56 2.71 3.075 2.873 ;
      RECT 2.646 2.68 3.07 2.879 ;
      RECT 2.73 2.655 3.045 2.884 ;
      RECT 2.895 2.637 3.04 2.895 ;
      RECT 2.895 2.632 2.995 2.895 ;
      RECT 2.981 2.626 2.995 2.895 ;
      RECT 2.37 1.95 2.375 2.349 ;
      RECT 2.115 1.95 2.15 2.347 ;
      RECT 1.71 1.985 1.715 2.341 ;
      RECT 2.455 1.988 2.46 2.243 ;
      RECT 2.45 1.986 2.455 2.249 ;
      RECT 2.445 1.985 2.45 2.256 ;
      RECT 2.42 1.978 2.445 2.28 ;
      RECT 2.415 1.971 2.42 2.304 ;
      RECT 2.41 1.967 2.415 2.313 ;
      RECT 2.4 1.962 2.41 2.326 ;
      RECT 2.395 1.959 2.4 2.335 ;
      RECT 2.39 1.957 2.395 2.34 ;
      RECT 2.375 1.953 2.39 2.35 ;
      RECT 2.36 1.947 2.37 2.349 ;
      RECT 2.322 1.945 2.36 2.349 ;
      RECT 2.236 1.947 2.322 2.349 ;
      RECT 2.15 1.949 2.236 2.348 ;
      RECT 2.079 1.95 2.115 2.347 ;
      RECT 1.993 1.952 2.079 2.347 ;
      RECT 1.907 1.954 1.993 2.346 ;
      RECT 1.821 1.956 1.907 2.346 ;
      RECT 1.735 1.959 1.821 2.345 ;
      RECT 1.725 1.965 1.735 2.344 ;
      RECT 1.715 1.977 1.725 2.342 ;
      RECT 1.655 2.012 1.71 2.338 ;
      RECT 1.65 2.042 1.655 2.1 ;
      RECT 2.395 3.122 2.41 3.315 ;
      RECT 2.39 3.09 2.395 3.315 ;
      RECT 2.38 3.065 2.39 3.315 ;
      RECT 2.375 3.037 2.38 3.315 ;
      RECT 2.345 2.96 2.375 3.315 ;
      RECT 2.32 2.842 2.345 3.315 ;
      RECT 2.315 2.78 2.32 3.315 ;
      RECT 2.305 2.767 2.315 3.315 ;
      RECT 2.285 2.757 2.305 3.315 ;
      RECT 2.27 2.74 2.285 3.315 ;
      RECT 2.24 2.728 2.27 3.315 ;
      RECT 2.235 2.727 2.24 3.26 ;
      RECT 2.23 2.727 2.235 3.218 ;
      RECT 2.215 2.726 2.23 3.17 ;
      RECT 2.2 2.726 2.215 3.108 ;
      RECT 2.18 2.726 2.2 3.068 ;
      RECT 2.175 2.726 2.18 3.053 ;
      RECT 2.15 2.725 2.175 3.048 ;
      RECT 2.08 2.724 2.15 3.035 ;
      RECT 2.065 2.723 2.08 3.02 ;
      RECT 2.035 2.722 2.065 3.003 ;
      RECT 2.03 2.722 2.035 2.988 ;
      RECT 1.98 2.721 2.03 2.968 ;
      RECT 1.915 2.72 1.98 2.923 ;
      RECT 1.91 2.72 1.915 2.895 ;
      RECT 1.995 3.257 2 3.514 ;
      RECT 1.975 3.176 1.995 3.531 ;
      RECT 1.955 3.17 1.975 3.56 ;
      RECT 1.895 3.157 1.955 3.58 ;
      RECT 1.85 3.141 1.895 3.581 ;
      RECT 1.766 3.129 1.85 3.569 ;
      RECT 1.68 3.116 1.766 3.553 ;
      RECT 1.67 3.109 1.68 3.545 ;
      RECT 1.625 3.106 1.67 3.485 ;
      RECT 1.605 3.102 1.625 3.4 ;
      RECT 1.59 3.1 1.605 3.353 ;
      RECT 1.56 3.097 1.59 3.323 ;
      RECT 1.525 3.093 1.56 3.3 ;
      RECT 1.482 3.088 1.525 3.288 ;
      RECT 1.396 3.079 1.482 3.297 ;
      RECT 1.31 3.068 1.396 3.309 ;
      RECT 1.245 3.059 1.31 3.318 ;
      RECT 1.225 3.05 1.245 3.323 ;
      RECT 1.22 3.043 1.225 3.325 ;
      RECT 1.18 3.028 1.22 3.322 ;
      RECT 1.16 3.007 1.18 3.317 ;
      RECT 1.145 2.995 1.16 3.31 ;
      RECT 1.14 2.987 1.145 3.303 ;
      RECT 1.125 2.967 1.14 3.296 ;
      RECT 1.12 2.83 1.125 3.29 ;
      RECT 1.04 2.719 1.12 3.262 ;
      RECT 1.031 2.712 1.04 3.228 ;
      RECT 0.945 2.706 1.031 3.153 ;
      RECT 0.92 2.697 0.945 3.065 ;
      RECT 0.89 2.692 0.92 3.04 ;
      RECT 0.825 2.701 0.89 3.025 ;
      RECT 0.805 2.717 0.825 3 ;
      RECT 0.795 2.723 0.805 2.948 ;
      RECT 0.775 2.745 0.795 2.83 ;
      RECT 1.43 2.71 1.6 2.895 ;
      RECT 1.43 2.71 1.635 2.893 ;
      RECT 1.48 2.62 1.65 2.884 ;
      RECT 1.43 2.777 1.655 2.877 ;
      RECT 1.445 2.655 1.65 2.884 ;
      RECT 0.645 3.388 0.71 3.831 ;
      RECT 0.585 3.413 0.71 3.829 ;
      RECT 0.585 3.413 0.765 3.823 ;
      RECT 0.57 3.438 0.765 3.822 ;
      RECT 0.71 3.375 0.785 3.819 ;
      RECT 0.645 3.4 0.865 3.813 ;
      RECT 0.57 3.439 0.91 3.807 ;
      RECT 0.555 3.466 0.91 3.798 ;
      RECT 0.57 3.459 0.93 3.79 ;
      RECT 0.555 3.468 0.935 3.773 ;
      RECT 0.55 3.485 0.935 3.6 ;
      RECT 0.555 2.207 0.59 2.445 ;
      RECT 0.555 2.207 0.62 2.444 ;
      RECT 0.555 2.207 0.735 2.44 ;
      RECT 0.555 2.207 0.79 2.418 ;
      RECT 0.565 2.15 0.845 2.318 ;
      RECT 0.67 1.99 0.7 2.441 ;
      RECT 0.7 1.985 0.88 2.198 ;
      RECT 0.57 2.126 0.88 2.198 ;
      RECT 0.62 2.022 0.67 2.442 ;
      RECT 0.59 2.078 0.88 2.198 ;
      RECT 89.065 0.575 89.235 1.085 ;
      RECT 89.065 2.395 89.235 3.865 ;
      RECT 89.065 5.015 89.235 6.485 ;
      RECT 89.065 7.795 89.235 8.305 ;
      RECT 88.075 0.575 88.245 1.085 ;
      RECT 88.075 2.395 88.245 3.865 ;
      RECT 88.075 5.015 88.245 6.485 ;
      RECT 88.075 7.795 88.245 8.305 ;
      RECT 86.71 0.575 86.88 3.865 ;
      RECT 86.71 5.015 86.88 8.305 ;
      RECT 86.28 0.575 86.45 1.085 ;
      RECT 86.28 1.655 86.45 3.865 ;
      RECT 86.28 5.015 86.45 7.225 ;
      RECT 86.28 7.795 86.45 8.305 ;
      RECT 84.91 1.66 85.08 2.935 ;
      RECT 84.91 5.945 85.08 7.22 ;
      RECT 71.145 0.575 71.315 1.085 ;
      RECT 71.145 2.395 71.315 3.865 ;
      RECT 71.145 5.015 71.315 6.485 ;
      RECT 71.145 7.795 71.315 8.305 ;
      RECT 70.155 0.575 70.325 1.085 ;
      RECT 70.155 2.395 70.325 3.865 ;
      RECT 70.155 5.015 70.325 6.485 ;
      RECT 70.155 7.795 70.325 8.305 ;
      RECT 68.79 0.575 68.96 3.865 ;
      RECT 68.79 5.015 68.96 8.305 ;
      RECT 68.36 0.575 68.53 1.085 ;
      RECT 68.36 1.655 68.53 3.865 ;
      RECT 68.36 5.015 68.53 7.225 ;
      RECT 68.36 7.795 68.53 8.305 ;
      RECT 66.99 1.66 67.16 2.935 ;
      RECT 66.99 5.945 67.16 7.22 ;
      RECT 53.225 0.575 53.395 1.085 ;
      RECT 53.225 2.395 53.395 3.865 ;
      RECT 53.225 5.015 53.395 6.485 ;
      RECT 53.225 7.795 53.395 8.305 ;
      RECT 52.235 0.575 52.405 1.085 ;
      RECT 52.235 2.395 52.405 3.865 ;
      RECT 52.235 5.015 52.405 6.485 ;
      RECT 52.235 7.795 52.405 8.305 ;
      RECT 50.87 0.575 51.04 3.865 ;
      RECT 50.87 5.015 51.04 8.305 ;
      RECT 50.44 0.575 50.61 1.085 ;
      RECT 50.44 1.655 50.61 3.865 ;
      RECT 50.44 5.015 50.61 7.225 ;
      RECT 50.44 7.795 50.61 8.305 ;
      RECT 49.07 1.66 49.24 2.935 ;
      RECT 49.07 5.945 49.24 7.22 ;
      RECT 35.31 0.575 35.48 1.085 ;
      RECT 35.31 2.395 35.48 3.865 ;
      RECT 35.31 5.015 35.48 6.485 ;
      RECT 35.31 7.795 35.48 8.305 ;
      RECT 34.32 0.575 34.49 1.085 ;
      RECT 34.32 2.395 34.49 3.865 ;
      RECT 34.32 5.015 34.49 6.485 ;
      RECT 34.32 7.795 34.49 8.305 ;
      RECT 32.955 0.575 33.125 3.865 ;
      RECT 32.955 5.015 33.125 8.305 ;
      RECT 32.525 0.575 32.695 1.085 ;
      RECT 32.525 1.655 32.695 3.865 ;
      RECT 32.525 5.015 32.695 7.225 ;
      RECT 32.525 7.795 32.695 8.305 ;
      RECT 31.155 1.66 31.325 2.935 ;
      RECT 31.155 5.945 31.325 7.22 ;
      RECT 17.39 0.575 17.56 1.085 ;
      RECT 17.39 2.395 17.56 3.865 ;
      RECT 17.39 5.015 17.56 6.485 ;
      RECT 17.39 7.795 17.56 8.305 ;
      RECT 16.4 0.575 16.57 1.085 ;
      RECT 16.4 2.395 16.57 3.865 ;
      RECT 16.4 5.015 16.57 6.485 ;
      RECT 16.4 7.795 16.57 8.305 ;
      RECT 15.035 0.575 15.205 3.865 ;
      RECT 15.035 5.015 15.205 8.305 ;
      RECT 14.605 0.575 14.775 1.085 ;
      RECT 14.605 1.655 14.775 3.865 ;
      RECT 14.605 5.015 14.775 7.225 ;
      RECT 14.605 7.795 14.775 8.305 ;
      RECT 13.235 1.66 13.405 2.935 ;
      RECT 13.235 5.945 13.405 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2at_8

MACRO sky130_osu_ring_oscillator_mpr2ca_8
  CLASS CORE ;
  ORIGIN -4 1.605 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ca_8 4 -1.605 ;
  SIZE 71.165 BY 8.88 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT 67.07 1.13 67.4 1.46 ;
      RECT 67.07 1.145 67.87 1.445 ;
      RECT 67.07 2.15 67.4 2.48 ;
      RECT 67.07 2.165 67.87 2.465 ;
      RECT 67.075 2.1 67.375 2.48 ;
      RECT 66.39 4.19 66.72 4.52 ;
      RECT 66.39 4.205 67.19 4.505 ;
      RECT 66.395 4.185 66.695 4.52 ;
      RECT 66.37 1.47 66.7 1.8 ;
      RECT 65.9 1.485 66.7 1.785 ;
      RECT 66.395 1.455 66.695 1.8 ;
      RECT 65.71 3.17 66.04 3.5 ;
      RECT 65.71 3.185 66.51 3.485 ;
      RECT 65.345 4.19 65.675 4.52 ;
      RECT 64.875 4.205 65.675 4.505 ;
      RECT 65.03 0.785 65.36 1.115 ;
      RECT 64.56 0.805 64.92 1.105 ;
      RECT 64.92 0.8 65.36 1.1 ;
      RECT 64.64 4.885 64.94 5.3 ;
      RECT 64.67 4.87 65 5.2 ;
      RECT 64.2 4.885 65 5.185 ;
      RECT 52.895 1.13 53.225 1.46 ;
      RECT 52.895 1.145 53.695 1.445 ;
      RECT 52.895 2.15 53.225 2.48 ;
      RECT 52.895 2.165 53.695 2.465 ;
      RECT 52.9 2.1 53.2 2.48 ;
      RECT 52.215 4.19 52.545 4.52 ;
      RECT 52.215 4.205 53.015 4.505 ;
      RECT 52.22 4.185 52.52 4.52 ;
      RECT 52.195 1.47 52.525 1.8 ;
      RECT 51.725 1.485 52.525 1.785 ;
      RECT 52.22 1.455 52.52 1.8 ;
      RECT 51.535 3.17 51.865 3.5 ;
      RECT 51.535 3.185 52.335 3.485 ;
      RECT 51.17 4.19 51.5 4.52 ;
      RECT 50.7 4.205 51.5 4.505 ;
      RECT 50.855 0.785 51.185 1.115 ;
      RECT 50.385 0.805 50.745 1.105 ;
      RECT 50.745 0.8 51.185 1.1 ;
      RECT 50.465 4.885 50.765 5.3 ;
      RECT 50.495 4.87 50.825 5.2 ;
      RECT 50.025 4.885 50.825 5.185 ;
      RECT 38.725 1.13 39.055 1.46 ;
      RECT 38.725 1.145 39.525 1.445 ;
      RECT 38.725 2.15 39.055 2.48 ;
      RECT 38.725 2.165 39.525 2.465 ;
      RECT 38.73 2.1 39.03 2.48 ;
      RECT 38.045 4.19 38.375 4.52 ;
      RECT 38.045 4.205 38.845 4.505 ;
      RECT 38.05 4.185 38.35 4.52 ;
      RECT 38.025 1.47 38.355 1.8 ;
      RECT 37.555 1.485 38.355 1.785 ;
      RECT 38.05 1.455 38.35 1.8 ;
      RECT 37.365 3.17 37.695 3.5 ;
      RECT 37.365 3.185 38.165 3.485 ;
      RECT 37 4.19 37.33 4.52 ;
      RECT 36.53 4.205 37.33 4.505 ;
      RECT 36.685 0.785 37.015 1.115 ;
      RECT 36.215 0.805 36.575 1.105 ;
      RECT 36.575 0.8 37.015 1.1 ;
      RECT 36.295 4.885 36.595 5.3 ;
      RECT 36.325 4.87 36.655 5.2 ;
      RECT 35.855 4.885 36.655 5.185 ;
      RECT 24.55 1.13 24.88 1.46 ;
      RECT 24.55 1.145 25.35 1.445 ;
      RECT 24.55 2.15 24.88 2.48 ;
      RECT 24.55 2.165 25.35 2.465 ;
      RECT 24.555 2.1 24.855 2.48 ;
      RECT 23.87 4.19 24.2 4.52 ;
      RECT 23.87 4.205 24.67 4.505 ;
      RECT 23.875 4.185 24.175 4.52 ;
      RECT 23.85 1.47 24.18 1.8 ;
      RECT 23.38 1.485 24.18 1.785 ;
      RECT 23.875 1.455 24.175 1.8 ;
      RECT 23.19 3.17 23.52 3.5 ;
      RECT 23.19 3.185 23.99 3.485 ;
      RECT 22.825 4.19 23.155 4.52 ;
      RECT 22.355 4.205 23.155 4.505 ;
      RECT 22.51 0.785 22.84 1.115 ;
      RECT 22.04 0.805 22.4 1.105 ;
      RECT 22.4 0.8 22.84 1.1 ;
      RECT 22.12 4.885 22.42 5.3 ;
      RECT 22.15 4.87 22.48 5.2 ;
      RECT 21.68 4.885 22.48 5.185 ;
      RECT 10.38 1.13 10.71 1.46 ;
      RECT 10.38 1.145 11.18 1.445 ;
      RECT 10.38 2.15 10.71 2.48 ;
      RECT 10.38 2.165 11.18 2.465 ;
      RECT 10.385 2.1 10.685 2.48 ;
      RECT 9.7 4.19 10.03 4.52 ;
      RECT 9.7 4.205 10.5 4.505 ;
      RECT 9.705 4.185 10.005 4.52 ;
      RECT 9.68 1.47 10.01 1.8 ;
      RECT 9.21 1.485 10.01 1.785 ;
      RECT 9.705 1.455 10.005 1.8 ;
      RECT 9.02 3.17 9.35 3.5 ;
      RECT 9.02 3.185 9.82 3.485 ;
      RECT 8.655 4.19 8.985 4.52 ;
      RECT 8.185 4.205 8.985 4.505 ;
      RECT 8.34 0.785 8.67 1.115 ;
      RECT 7.87 0.805 8.23 1.105 ;
      RECT 8.23 0.8 8.67 1.1 ;
      RECT 7.95 4.885 8.25 5.3 ;
      RECT 7.98 4.87 8.31 5.2 ;
      RECT 7.51 4.885 8.31 5.185 ;
    LAYER via2 ;
      RECT 67.135 1.195 67.335 1.395 ;
      RECT 67.135 2.215 67.335 2.415 ;
      RECT 66.455 4.255 66.655 4.455 ;
      RECT 66.435 1.535 66.635 1.735 ;
      RECT 65.775 3.235 65.975 3.435 ;
      RECT 65.41 4.255 65.61 4.455 ;
      RECT 65.095 0.85 65.295 1.05 ;
      RECT 64.735 4.935 64.935 5.135 ;
      RECT 52.96 1.195 53.16 1.395 ;
      RECT 52.96 2.215 53.16 2.415 ;
      RECT 52.28 4.255 52.48 4.455 ;
      RECT 52.26 1.535 52.46 1.735 ;
      RECT 51.6 3.235 51.8 3.435 ;
      RECT 51.235 4.255 51.435 4.455 ;
      RECT 50.92 0.85 51.12 1.05 ;
      RECT 50.56 4.935 50.76 5.135 ;
      RECT 38.79 1.195 38.99 1.395 ;
      RECT 38.79 2.215 38.99 2.415 ;
      RECT 38.11 4.255 38.31 4.455 ;
      RECT 38.09 1.535 38.29 1.735 ;
      RECT 37.43 3.235 37.63 3.435 ;
      RECT 37.065 4.255 37.265 4.455 ;
      RECT 36.75 0.85 36.95 1.05 ;
      RECT 36.39 4.935 36.59 5.135 ;
      RECT 24.615 1.195 24.815 1.395 ;
      RECT 24.615 2.215 24.815 2.415 ;
      RECT 23.935 4.255 24.135 4.455 ;
      RECT 23.915 1.535 24.115 1.735 ;
      RECT 23.255 3.235 23.455 3.435 ;
      RECT 22.89 4.255 23.09 4.455 ;
      RECT 22.575 0.85 22.775 1.05 ;
      RECT 22.215 4.935 22.415 5.135 ;
      RECT 10.445 1.195 10.645 1.395 ;
      RECT 10.445 2.215 10.645 2.415 ;
      RECT 9.765 4.255 9.965 4.455 ;
      RECT 9.745 1.535 9.945 1.735 ;
      RECT 9.085 3.235 9.285 3.435 ;
      RECT 8.72 4.255 8.92 4.455 ;
      RECT 8.405 0.85 8.605 1.05 ;
      RECT 8.045 4.935 8.245 5.135 ;
    LAYER met2 ;
      RECT 14.745 4.675 15.065 5 ;
      RECT 14.775 4.09 14.945 5 ;
      RECT 14.775 4.09 14.95 4.44 ;
      RECT 14.775 4.09 15.75 4.265 ;
      RECT 15.575 0.36 15.75 4.265 ;
      RECT 13.075 0.39 13.4 0.715 ;
      RECT 15.52 0.36 15.87 0.71 ;
      RECT 13.075 0.42 15.87 0.59 ;
      RECT 13.135 -1.355 13.3 0.715 ;
      RECT 74.605 -0.51 74.955 -0.16 ;
      RECT 74.64 -1.355 74.805 -0.16 ;
      RECT 13.135 -1.355 74.805 -1.19 ;
      RECT 71.435 4.675 71.755 5 ;
      RECT 71.465 4.09 71.635 5 ;
      RECT 71.465 4.09 71.64 4.44 ;
      RECT 71.465 4.09 72.44 4.265 ;
      RECT 72.265 0.36 72.44 4.265 ;
      RECT 69.765 0.39 70.09 0.715 ;
      RECT 72.21 0.36 72.56 0.71 ;
      RECT 69.765 0.42 72.56 0.59 ;
      RECT 70.67 -0.48 70.83 0.59 ;
      RECT 60.42 -0.51 60.77 -0.16 ;
      RECT 60.42 -0.48 70.83 -0.32 ;
      RECT 60.455 -0.515 60.62 -0.16 ;
      RECT 72.235 5.05 72.56 5.375 ;
      RECT 71.12 5.14 72.56 5.31 ;
      RECT 71.12 0.79 71.28 5.31 ;
      RECT 69.18 1.58 69.505 1.905 ;
      RECT 69.18 1.62 71.28 1.795 ;
      RECT 69.225 0 69.425 1.905 ;
      RECT 65.055 0.765 65.335 1.135 ;
      RECT 71.435 0.76 71.755 1.08 ;
      RECT 71.12 0.79 71.755 0.96 ;
      RECT 65.075 0 65.275 1.135 ;
      RECT 65.075 0 69.425 0.2 ;
      RECT 70.395 4.26 70.72 4.585 ;
      RECT 70.46 2.03 70.635 4.585 ;
      RECT 70.39 2.03 70.715 2.355 ;
      RECT 64.695 4.85 64.975 5.22 ;
      RECT 64.695 5.02 69.97 5.185 ;
      RECT 69.805 2.05 69.97 5.185 ;
      RECT 69.68 2.05 70.005 2.375 ;
      RECT 68.795 3.175 69.055 3.495 ;
      RECT 68.855 1.135 68.995 3.495 ;
      RECT 68.795 1.135 69.055 1.455 ;
      RECT 67.775 4.195 68.035 4.515 ;
      RECT 67.155 4.285 68.035 4.425 ;
      RECT 67.155 2.13 67.295 4.425 ;
      RECT 67.095 2.13 67.375 2.5 ;
      RECT 66.415 4.17 66.695 4.54 ;
      RECT 66.475 2.245 66.615 4.54 ;
      RECT 66.475 2.245 66.955 2.385 ;
      RECT 66.815 0.455 66.955 2.385 ;
      RECT 66.755 0.455 67.015 0.775 ;
      RECT 65.735 3.15 66.015 3.52 ;
      RECT 65.795 0.795 65.935 3.52 ;
      RECT 65.735 0.795 65.995 1.115 ;
      RECT 65.37 4.17 65.65 4.54 ;
      RECT 65.37 4.195 65.655 4.515 ;
      RECT 57.26 4.675 57.58 5 ;
      RECT 57.29 4.09 57.46 5 ;
      RECT 57.29 4.09 57.465 4.44 ;
      RECT 57.29 4.09 58.265 4.265 ;
      RECT 58.09 0.36 58.265 4.265 ;
      RECT 55.59 0.39 55.915 0.715 ;
      RECT 58.035 0.36 58.385 0.71 ;
      RECT 55.59 0.42 58.385 0.59 ;
      RECT 56.385 -0.475 56.535 0.59 ;
      RECT 46.25 -0.505 46.6 -0.155 ;
      RECT 46.25 -0.475 56.535 -0.325 ;
      RECT 46.285 -0.51 46.45 -0.155 ;
      RECT 58.06 5.05 58.385 5.375 ;
      RECT 56.945 5.14 58.385 5.31 ;
      RECT 56.945 0.79 57.105 5.31 ;
      RECT 55.005 1.58 55.33 1.905 ;
      RECT 55.005 1.62 57.105 1.795 ;
      RECT 55.05 0 55.25 1.905 ;
      RECT 50.88 0.765 51.16 1.135 ;
      RECT 57.26 0.76 57.58 1.08 ;
      RECT 56.945 0.79 57.58 0.96 ;
      RECT 50.9 0 51.1 1.135 ;
      RECT 50.9 0 55.25 0.2 ;
      RECT 56.22 4.26 56.545 4.585 ;
      RECT 56.285 2.03 56.46 4.585 ;
      RECT 56.215 2.03 56.54 2.355 ;
      RECT 50.52 4.85 50.8 5.22 ;
      RECT 50.52 5.02 55.795 5.185 ;
      RECT 55.63 2.05 55.795 5.185 ;
      RECT 55.505 2.05 55.83 2.375 ;
      RECT 54.62 3.175 54.88 3.495 ;
      RECT 54.68 1.135 54.82 3.495 ;
      RECT 54.62 1.135 54.88 1.455 ;
      RECT 53.6 4.195 53.86 4.515 ;
      RECT 52.98 4.285 53.86 4.425 ;
      RECT 52.98 2.13 53.12 4.425 ;
      RECT 52.92 2.13 53.2 2.5 ;
      RECT 52.24 4.17 52.52 4.54 ;
      RECT 52.3 2.245 52.44 4.54 ;
      RECT 52.3 2.245 52.78 2.385 ;
      RECT 52.64 0.455 52.78 2.385 ;
      RECT 52.58 0.455 52.84 0.775 ;
      RECT 51.56 3.15 51.84 3.52 ;
      RECT 51.62 0.795 51.76 3.52 ;
      RECT 51.56 0.795 51.82 1.115 ;
      RECT 51.195 4.17 51.475 4.54 ;
      RECT 51.195 4.195 51.48 4.515 ;
      RECT 43.09 4.675 43.41 5 ;
      RECT 43.12 4.09 43.29 5 ;
      RECT 43.12 4.09 43.295 4.44 ;
      RECT 43.12 4.09 44.095 4.265 ;
      RECT 43.92 0.36 44.095 4.265 ;
      RECT 41.42 0.39 41.745 0.715 ;
      RECT 43.865 0.36 44.215 0.71 ;
      RECT 41.42 0.42 44.215 0.59 ;
      RECT 41.98 -0.49 42.16 0.59 ;
      RECT 32.075 -0.52 32.425 -0.17 ;
      RECT 32.075 -0.49 42.16 -0.31 ;
      RECT 32.11 -0.525 32.275 -0.17 ;
      RECT 43.89 5.05 44.215 5.375 ;
      RECT 42.775 5.14 44.215 5.31 ;
      RECT 42.775 0.79 42.935 5.31 ;
      RECT 40.835 1.58 41.16 1.905 ;
      RECT 40.835 1.62 42.935 1.795 ;
      RECT 40.88 0 41.08 1.905 ;
      RECT 36.71 0.765 36.99 1.135 ;
      RECT 43.09 0.76 43.41 1.08 ;
      RECT 42.775 0.79 43.41 0.96 ;
      RECT 36.73 0 36.93 1.135 ;
      RECT 36.73 0 41.08 0.2 ;
      RECT 42.05 4.26 42.375 4.585 ;
      RECT 42.115 2.03 42.29 4.585 ;
      RECT 42.045 2.03 42.37 2.355 ;
      RECT 36.35 4.85 36.63 5.22 ;
      RECT 36.35 5.02 41.625 5.185 ;
      RECT 41.46 2.05 41.625 5.185 ;
      RECT 41.335 2.05 41.66 2.375 ;
      RECT 40.45 3.175 40.71 3.495 ;
      RECT 40.51 1.135 40.65 3.495 ;
      RECT 40.45 1.135 40.71 1.455 ;
      RECT 39.43 4.195 39.69 4.515 ;
      RECT 38.81 4.285 39.69 4.425 ;
      RECT 38.81 2.13 38.95 4.425 ;
      RECT 38.75 2.13 39.03 2.5 ;
      RECT 38.07 4.17 38.35 4.54 ;
      RECT 38.13 2.245 38.27 4.54 ;
      RECT 38.13 2.245 38.61 2.385 ;
      RECT 38.47 0.455 38.61 2.385 ;
      RECT 38.41 0.455 38.67 0.775 ;
      RECT 37.39 3.15 37.67 3.52 ;
      RECT 37.45 0.795 37.59 3.52 ;
      RECT 37.39 0.795 37.65 1.115 ;
      RECT 37.025 4.17 37.305 4.54 ;
      RECT 37.025 4.195 37.31 4.515 ;
      RECT 28.915 4.675 29.235 5 ;
      RECT 28.945 4.09 29.115 5 ;
      RECT 28.945 4.09 29.12 4.44 ;
      RECT 28.945 4.09 29.92 4.265 ;
      RECT 29.745 0.36 29.92 4.265 ;
      RECT 27.245 0.39 27.57 0.715 ;
      RECT 29.69 0.36 30.04 0.71 ;
      RECT 27.245 0.42 30.04 0.59 ;
      RECT 27.34 -0.48 27.53 0.715 ;
      RECT 17.91 -0.51 18.26 -0.16 ;
      RECT 17.91 -0.48 27.53 -0.29 ;
      RECT 17.945 -0.515 18.11 -0.16 ;
      RECT 29.715 5.05 30.04 5.375 ;
      RECT 28.6 5.14 30.04 5.31 ;
      RECT 28.6 0.79 28.76 5.31 ;
      RECT 26.66 1.58 26.985 1.905 ;
      RECT 26.66 1.62 28.76 1.795 ;
      RECT 26.705 0 26.905 1.905 ;
      RECT 22.535 0.765 22.815 1.135 ;
      RECT 28.915 0.76 29.235 1.08 ;
      RECT 28.6 0.79 29.235 0.96 ;
      RECT 22.555 0 22.755 1.135 ;
      RECT 22.555 0 26.905 0.2 ;
      RECT 27.875 4.26 28.2 4.585 ;
      RECT 27.94 2.03 28.115 4.585 ;
      RECT 27.87 2.03 28.195 2.355 ;
      RECT 22.175 4.85 22.455 5.22 ;
      RECT 22.175 5.02 27.45 5.185 ;
      RECT 27.285 2.05 27.45 5.185 ;
      RECT 27.16 2.05 27.485 2.375 ;
      RECT 26.275 3.175 26.535 3.495 ;
      RECT 26.335 1.135 26.475 3.495 ;
      RECT 26.275 1.135 26.535 1.455 ;
      RECT 25.255 4.195 25.515 4.515 ;
      RECT 24.635 4.285 25.515 4.425 ;
      RECT 24.635 2.13 24.775 4.425 ;
      RECT 24.575 2.13 24.855 2.5 ;
      RECT 23.895 4.17 24.175 4.54 ;
      RECT 23.955 2.245 24.095 4.54 ;
      RECT 23.955 2.245 24.435 2.385 ;
      RECT 24.295 0.455 24.435 2.385 ;
      RECT 24.235 0.455 24.495 0.775 ;
      RECT 23.215 3.15 23.495 3.52 ;
      RECT 23.275 0.795 23.415 3.52 ;
      RECT 23.215 0.795 23.475 1.115 ;
      RECT 22.85 4.17 23.13 4.54 ;
      RECT 22.85 4.195 23.135 4.515 ;
      RECT 15.545 5.05 15.87 5.375 ;
      RECT 14.43 5.14 15.87 5.31 ;
      RECT 14.43 0.79 14.59 5.31 ;
      RECT 12.49 1.58 12.815 1.905 ;
      RECT 12.49 1.62 14.59 1.795 ;
      RECT 12.535 0 12.735 1.905 ;
      RECT 8.365 0.765 8.645 1.135 ;
      RECT 14.745 0.76 15.065 1.08 ;
      RECT 14.43 0.79 15.065 0.96 ;
      RECT 8.385 0 8.585 1.135 ;
      RECT 8.385 0 12.735 0.2 ;
      RECT 13.705 4.26 14.03 4.585 ;
      RECT 13.77 2.03 13.945 4.585 ;
      RECT 13.7 2.03 14.025 2.355 ;
      RECT 8.005 4.85 8.285 5.22 ;
      RECT 8.005 5.02 13.28 5.185 ;
      RECT 13.115 2.05 13.28 5.185 ;
      RECT 12.99 2.05 13.315 2.375 ;
      RECT 12.105 3.175 12.365 3.495 ;
      RECT 12.165 1.135 12.305 3.495 ;
      RECT 12.105 1.135 12.365 1.455 ;
      RECT 11.085 4.195 11.345 4.515 ;
      RECT 10.465 4.285 11.345 4.425 ;
      RECT 10.465 2.13 10.605 4.425 ;
      RECT 10.405 2.13 10.685 2.5 ;
      RECT 9.725 4.17 10.005 4.54 ;
      RECT 9.785 2.245 9.925 4.54 ;
      RECT 9.785 2.245 10.265 2.385 ;
      RECT 10.125 0.455 10.265 2.385 ;
      RECT 10.065 0.455 10.325 0.775 ;
      RECT 9.045 3.15 9.325 3.52 ;
      RECT 9.105 0.795 9.245 3.52 ;
      RECT 9.045 0.795 9.305 1.115 ;
      RECT 8.68 4.17 8.96 4.54 ;
      RECT 8.68 4.195 8.965 4.515 ;
      RECT 67.095 1.11 67.375 1.48 ;
      RECT 66.395 1.45 66.675 1.82 ;
      RECT 52.92 1.11 53.2 1.48 ;
      RECT 52.22 1.45 52.5 1.82 ;
      RECT 38.75 1.11 39.03 1.48 ;
      RECT 38.05 1.45 38.33 1.82 ;
      RECT 24.575 1.11 24.855 1.48 ;
      RECT 23.875 1.45 24.155 1.82 ;
      RECT 10.405 1.11 10.685 1.48 ;
      RECT 9.705 1.45 9.985 1.82 ;
    LAYER via1 ;
      RECT 74.705 -0.41 74.855 -0.26 ;
      RECT 72.325 5.135 72.475 5.285 ;
      RECT 72.31 0.46 72.46 0.61 ;
      RECT 71.52 0.845 71.67 0.995 ;
      RECT 71.52 4.765 71.67 4.915 ;
      RECT 70.485 4.345 70.635 4.495 ;
      RECT 70.48 2.115 70.63 2.265 ;
      RECT 69.855 0.475 70.005 0.625 ;
      RECT 69.77 2.135 69.92 2.285 ;
      RECT 69.27 1.665 69.42 1.815 ;
      RECT 68.85 1.22 69 1.37 ;
      RECT 68.85 3.26 69 3.41 ;
      RECT 67.83 4.28 67.98 4.43 ;
      RECT 67.15 1.22 67.3 1.37 ;
      RECT 67.15 2.24 67.3 2.39 ;
      RECT 66.81 0.54 66.96 0.69 ;
      RECT 66.47 1.56 66.62 1.71 ;
      RECT 66.47 4.28 66.62 4.43 ;
      RECT 65.79 0.88 65.94 1.03 ;
      RECT 65.79 3.26 65.94 3.41 ;
      RECT 65.45 4.28 65.6 4.43 ;
      RECT 65.11 0.875 65.26 1.025 ;
      RECT 64.77 4.96 64.92 5.11 ;
      RECT 60.52 -0.41 60.67 -0.26 ;
      RECT 58.15 5.135 58.3 5.285 ;
      RECT 58.135 0.46 58.285 0.61 ;
      RECT 57.345 0.845 57.495 0.995 ;
      RECT 57.345 4.765 57.495 4.915 ;
      RECT 56.31 4.345 56.46 4.495 ;
      RECT 56.305 2.115 56.455 2.265 ;
      RECT 55.68 0.475 55.83 0.625 ;
      RECT 55.595 2.135 55.745 2.285 ;
      RECT 55.095 1.665 55.245 1.815 ;
      RECT 54.675 1.22 54.825 1.37 ;
      RECT 54.675 3.26 54.825 3.41 ;
      RECT 53.655 4.28 53.805 4.43 ;
      RECT 52.975 1.22 53.125 1.37 ;
      RECT 52.975 2.24 53.125 2.39 ;
      RECT 52.635 0.54 52.785 0.69 ;
      RECT 52.295 1.56 52.445 1.71 ;
      RECT 52.295 4.28 52.445 4.43 ;
      RECT 51.615 0.88 51.765 1.03 ;
      RECT 51.615 3.26 51.765 3.41 ;
      RECT 51.275 4.28 51.425 4.43 ;
      RECT 50.935 0.875 51.085 1.025 ;
      RECT 50.595 4.96 50.745 5.11 ;
      RECT 46.35 -0.405 46.5 -0.255 ;
      RECT 43.98 5.135 44.13 5.285 ;
      RECT 43.965 0.46 44.115 0.61 ;
      RECT 43.175 0.845 43.325 0.995 ;
      RECT 43.175 4.765 43.325 4.915 ;
      RECT 42.14 4.345 42.29 4.495 ;
      RECT 42.135 2.115 42.285 2.265 ;
      RECT 41.51 0.475 41.66 0.625 ;
      RECT 41.425 2.135 41.575 2.285 ;
      RECT 40.925 1.665 41.075 1.815 ;
      RECT 40.505 1.22 40.655 1.37 ;
      RECT 40.505 3.26 40.655 3.41 ;
      RECT 39.485 4.28 39.635 4.43 ;
      RECT 38.805 1.22 38.955 1.37 ;
      RECT 38.805 2.24 38.955 2.39 ;
      RECT 38.465 0.54 38.615 0.69 ;
      RECT 38.125 1.56 38.275 1.71 ;
      RECT 38.125 4.28 38.275 4.43 ;
      RECT 37.445 0.88 37.595 1.03 ;
      RECT 37.445 3.26 37.595 3.41 ;
      RECT 37.105 4.28 37.255 4.43 ;
      RECT 36.765 0.875 36.915 1.025 ;
      RECT 36.425 4.96 36.575 5.11 ;
      RECT 32.175 -0.42 32.325 -0.27 ;
      RECT 29.805 5.135 29.955 5.285 ;
      RECT 29.79 0.46 29.94 0.61 ;
      RECT 29 0.845 29.15 0.995 ;
      RECT 29 4.765 29.15 4.915 ;
      RECT 27.965 4.345 28.115 4.495 ;
      RECT 27.96 2.115 28.11 2.265 ;
      RECT 27.335 0.475 27.485 0.625 ;
      RECT 27.25 2.135 27.4 2.285 ;
      RECT 26.75 1.665 26.9 1.815 ;
      RECT 26.33 1.22 26.48 1.37 ;
      RECT 26.33 3.26 26.48 3.41 ;
      RECT 25.31 4.28 25.46 4.43 ;
      RECT 24.63 1.22 24.78 1.37 ;
      RECT 24.63 2.24 24.78 2.39 ;
      RECT 24.29 0.54 24.44 0.69 ;
      RECT 23.95 1.56 24.1 1.71 ;
      RECT 23.95 4.28 24.1 4.43 ;
      RECT 23.27 0.88 23.42 1.03 ;
      RECT 23.27 3.26 23.42 3.41 ;
      RECT 22.93 4.28 23.08 4.43 ;
      RECT 22.59 0.875 22.74 1.025 ;
      RECT 22.25 4.96 22.4 5.11 ;
      RECT 18.01 -0.41 18.16 -0.26 ;
      RECT 15.635 5.135 15.785 5.285 ;
      RECT 15.62 0.46 15.77 0.61 ;
      RECT 14.83 0.845 14.98 0.995 ;
      RECT 14.83 4.765 14.98 4.915 ;
      RECT 13.795 4.345 13.945 4.495 ;
      RECT 13.79 2.115 13.94 2.265 ;
      RECT 13.165 0.475 13.315 0.625 ;
      RECT 13.08 2.135 13.23 2.285 ;
      RECT 12.58 1.665 12.73 1.815 ;
      RECT 12.16 1.22 12.31 1.37 ;
      RECT 12.16 3.26 12.31 3.41 ;
      RECT 11.14 4.28 11.29 4.43 ;
      RECT 10.46 1.22 10.61 1.37 ;
      RECT 10.46 2.24 10.61 2.39 ;
      RECT 10.12 0.54 10.27 0.69 ;
      RECT 9.78 1.56 9.93 1.71 ;
      RECT 9.78 4.28 9.93 4.43 ;
      RECT 9.1 0.88 9.25 1.03 ;
      RECT 9.1 3.26 9.25 3.41 ;
      RECT 8.76 4.28 8.91 4.43 ;
      RECT 8.42 0.875 8.57 1.025 ;
      RECT 8.08 4.96 8.23 5.11 ;
    LAYER met1 ;
      RECT 62.295 -1.605 69.195 0.345 ;
      RECT 48.12 -1.605 55.02 0.345 ;
      RECT 33.95 -1.605 40.85 0.345 ;
      RECT 19.775 -1.605 26.675 0.345 ;
      RECT 5.605 -1.605 12.505 0.345 ;
      RECT 62.295 -1.605 69.385 0.19 ;
      RECT 48.12 -1.605 55.21 0.19 ;
      RECT 33.95 -1.605 41.04 0.19 ;
      RECT 19.775 -1.605 26.865 0.19 ;
      RECT 5.605 -1.605 12.695 0.19 ;
      RECT 62.04 -1.605 69.385 0.05 ;
      RECT 47.865 -1.605 55.21 0.05 ;
      RECT 33.695 -1.605 41.04 0.05 ;
      RECT 19.52 -1.605 26.865 0.05 ;
      RECT 5.35 -1.605 12.695 0.05 ;
      RECT 4.005 -1.605 75.165 -1.3 ;
      RECT 69.225 2.545 75.165 3.14 ;
      RECT 69.685 2.53 75.165 3.14 ;
      RECT 55.05 2.545 60.99 3.14 ;
      RECT 40.88 2.545 46.82 3.14 ;
      RECT 26.705 2.545 32.645 3.14 ;
      RECT 12.535 2.545 18.475 3.14 ;
      RECT 60.695 2.525 62.155 3.135 ;
      RECT 46.52 2.525 47.98 3.135 ;
      RECT 32.35 2.525 33.81 3.135 ;
      RECT 18.175 2.525 19.635 3.135 ;
      RECT 4.005 2.525 5.465 3.135 ;
      RECT 4.005 2.585 75.165 3.065 ;
      RECT 69.095 2.545 75.165 3.065 ;
      RECT 54.92 2.545 62.155 3.065 ;
      RECT 40.75 2.545 47.98 3.065 ;
      RECT 26.575 2.545 33.81 3.065 ;
      RECT 12.405 2.545 19.635 3.065 ;
      RECT 55.51 2.53 62.155 3.135 ;
      RECT 41.34 2.53 47.98 3.135 ;
      RECT 27.165 2.53 33.81 3.135 ;
      RECT 12.995 2.53 19.635 3.135 ;
      RECT 4.005 6.97 75.165 7.275 ;
      RECT 62 5.575 69.2 7.275 ;
      RECT 47.825 5.575 55.025 7.275 ;
      RECT 33.655 5.575 40.855 7.275 ;
      RECT 19.48 5.575 26.68 7.275 ;
      RECT 5.31 5.575 12.51 7.275 ;
      RECT 62.295 5.305 69.195 7.275 ;
      RECT 48.12 5.305 55.02 7.275 ;
      RECT 33.95 5.305 40.85 7.275 ;
      RECT 19.775 5.305 26.675 7.275 ;
      RECT 5.605 5.305 12.505 7.275 ;
      RECT 74.565 0.76 74.855 0.99 ;
      RECT 74.625 -0.72 74.795 0.99 ;
      RECT 74.605 -0.51 74.955 -0.16 ;
      RECT 74.565 -0.72 74.855 -0.49 ;
      RECT 74.565 6.16 74.855 6.39 ;
      RECT 74.625 4.68 74.795 6.39 ;
      RECT 74.565 4.68 74.855 4.91 ;
      RECT 74.155 1.13 74.485 1.36 ;
      RECT 74.155 1.16 74.655 1.33 ;
      RECT 74.155 0.79 74.345 1.36 ;
      RECT 73.575 0.76 73.865 0.99 ;
      RECT 73.575 0.79 74.345 0.96 ;
      RECT 73.635 -0.72 73.805 0.99 ;
      RECT 73.575 -0.72 73.865 -0.49 ;
      RECT 73.575 6.16 73.865 6.39 ;
      RECT 73.635 4.68 73.805 6.39 ;
      RECT 73.575 4.68 73.865 4.91 ;
      RECT 73.575 4.72 74.425 4.88 ;
      RECT 74.255 4.31 74.425 4.88 ;
      RECT 73.575 4.715 73.965 4.88 ;
      RECT 74.195 4.31 74.485 4.54 ;
      RECT 74.195 4.34 74.655 4.51 ;
      RECT 73.205 1.13 73.495 1.36 ;
      RECT 73.205 1.16 73.665 1.33 ;
      RECT 73.265 0.05 73.43 1.36 ;
      RECT 71.78 0.02 72.07 0.25 ;
      RECT 71.78 0.05 73.43 0.22 ;
      RECT 71.84 -0.72 72.01 0.25 ;
      RECT 71.78 -0.72 72.07 -0.49 ;
      RECT 71.78 6.16 72.07 6.39 ;
      RECT 71.84 5.42 72.01 6.39 ;
      RECT 71.84 5.515 73.43 5.685 ;
      RECT 73.26 4.31 73.43 5.685 ;
      RECT 71.78 5.42 72.07 5.65 ;
      RECT 73.205 4.31 73.495 4.54 ;
      RECT 73.205 4.34 73.665 4.51 ;
      RECT 72.21 0.36 72.56 0.71 ;
      RECT 72.04 0.42 72.56 0.59 ;
      RECT 72.235 5.05 72.56 5.375 ;
      RECT 72.21 5.05 72.56 5.28 ;
      RECT 72.04 5.08 72.56 5.25 ;
      RECT 71.435 0.76 71.755 1.08 ;
      RECT 71.405 0.76 71.755 0.99 ;
      RECT 71.12 0.79 71.755 0.96 ;
      RECT 71.435 4.675 71.755 5 ;
      RECT 71.405 4.68 71.755 4.91 ;
      RECT 71.235 4.71 71.755 4.88 ;
      RECT 70.39 2.03 70.715 2.355 ;
      RECT 70.465 1.13 70.645 2.355 ;
      RECT 70.41 1.13 70.7 1.36 ;
      RECT 70.41 1.16 70.87 1.33 ;
      RECT 70.395 4.26 70.72 4.585 ;
      RECT 70.395 4.34 70.87 4.51 ;
      RECT 69.685 2.05 70.005 2.39 ;
      RECT 69.68 2.05 70.005 2.065 ;
      RECT 69.805 0.39 69.97 2.39 ;
      RECT 69.765 0.39 70.09 0.715 ;
      RECT 68.765 1.165 69.085 1.425 ;
      RECT 68.49 1.225 69.085 1.365 ;
      RECT 66.385 1.505 66.705 1.765 ;
      RECT 68.36 1.52 68.65 1.75 ;
      RECT 66.385 1.565 68.65 1.705 ;
      RECT 67.745 4.225 68.065 4.485 ;
      RECT 67.745 4.285 68.34 4.425 ;
      RECT 67.065 1.165 67.385 1.425 ;
      RECT 62.325 1.18 62.615 1.41 ;
      RECT 62.325 1.225 67.385 1.365 ;
      RECT 67.155 0.885 67.295 1.425 ;
      RECT 67.155 0.885 67.635 1.025 ;
      RECT 67.495 0.5 67.635 1.025 ;
      RECT 67.42 0.5 67.71 0.73 ;
      RECT 67.065 2.185 67.385 2.445 ;
      RECT 66.4 2.2 66.69 2.43 ;
      RECT 64.19 2.2 64.48 2.43 ;
      RECT 64.19 2.245 67.385 2.385 ;
      RECT 65.365 4.225 65.685 4.485 ;
      RECT 67.08 4.24 67.37 4.47 ;
      RECT 64.7 4.24 64.99 4.47 ;
      RECT 64.7 4.285 65.685 4.425 ;
      RECT 67.155 3.945 67.295 4.47 ;
      RECT 65.455 3.945 65.595 4.485 ;
      RECT 65.455 3.945 67.295 4.085 ;
      RECT 64.36 0.84 64.65 1.07 ;
      RECT 64.435 0.545 64.575 1.07 ;
      RECT 66.725 0.485 67.045 0.745 ;
      RECT 66.625 0.5 67.045 0.73 ;
      RECT 64.435 0.545 67.045 0.685 ;
      RECT 65.705 0.825 66.025 1.085 ;
      RECT 65.705 0.885 66.3 1.025 ;
      RECT 64.685 4.905 65.005 5.165 ;
      RECT 63.755 4.965 66.105 5.105 ;
      RECT 65.965 4.24 66.105 5.105 ;
      RECT 63.755 4.24 63.895 5.105 ;
      RECT 65.89 4.24 66.18 4.47 ;
      RECT 63.68 4.24 63.97 4.47 ;
      RECT 65.705 3.205 66.025 3.465 ;
      RECT 63 3.22 63.29 3.45 ;
      RECT 63 3.265 66.025 3.405 ;
      RECT 65.03 0.785 65.36 1.115 ;
      RECT 65.025 0.82 65.36 1.08 ;
      RECT 65.375 0.84 65.49 1.07 ;
      RECT 65.025 0.835 65.375 1.065 ;
      RECT 65.025 0.885 65.505 1.025 ;
      RECT 64.91 0.885 64.92 1.025 ;
      RECT 64.92 0.88 65.49 1.02 ;
      RECT 60.39 0.76 60.68 0.99 ;
      RECT 60.45 -0.72 60.62 0.99 ;
      RECT 60.42 -0.51 60.77 -0.16 ;
      RECT 60.39 -0.72 60.68 -0.49 ;
      RECT 60.39 6.16 60.68 6.39 ;
      RECT 60.45 4.68 60.62 6.39 ;
      RECT 60.39 4.68 60.68 4.91 ;
      RECT 59.98 1.13 60.31 1.36 ;
      RECT 59.98 1.16 60.48 1.33 ;
      RECT 59.98 0.79 60.17 1.36 ;
      RECT 59.4 0.76 59.69 0.99 ;
      RECT 59.4 0.79 60.17 0.96 ;
      RECT 59.46 -0.72 59.63 0.99 ;
      RECT 59.4 -0.72 59.69 -0.49 ;
      RECT 59.4 6.16 59.69 6.39 ;
      RECT 59.46 4.68 59.63 6.39 ;
      RECT 59.4 4.68 59.69 4.91 ;
      RECT 59.4 4.72 60.25 4.88 ;
      RECT 60.08 4.31 60.25 4.88 ;
      RECT 59.4 4.715 59.79 4.88 ;
      RECT 60.02 4.31 60.31 4.54 ;
      RECT 60.02 4.34 60.48 4.51 ;
      RECT 59.03 1.13 59.32 1.36 ;
      RECT 59.03 1.16 59.49 1.33 ;
      RECT 59.09 0.05 59.255 1.36 ;
      RECT 57.605 0.02 57.895 0.25 ;
      RECT 57.605 0.05 59.255 0.22 ;
      RECT 57.665 -0.72 57.835 0.25 ;
      RECT 57.605 -0.72 57.895 -0.49 ;
      RECT 57.605 6.16 57.895 6.39 ;
      RECT 57.665 5.42 57.835 6.39 ;
      RECT 57.665 5.515 59.255 5.685 ;
      RECT 59.085 4.31 59.255 5.685 ;
      RECT 57.605 5.42 57.895 5.65 ;
      RECT 59.03 4.31 59.32 4.54 ;
      RECT 59.03 4.34 59.49 4.51 ;
      RECT 58.035 0.36 58.385 0.71 ;
      RECT 57.865 0.42 58.385 0.59 ;
      RECT 58.06 5.05 58.385 5.375 ;
      RECT 58.035 5.05 58.385 5.28 ;
      RECT 57.865 5.08 58.385 5.25 ;
      RECT 57.26 0.76 57.58 1.08 ;
      RECT 57.23 0.76 57.58 0.99 ;
      RECT 56.945 0.79 57.58 0.96 ;
      RECT 57.26 4.675 57.58 5 ;
      RECT 57.23 4.68 57.58 4.91 ;
      RECT 57.06 4.71 57.58 4.88 ;
      RECT 56.215 2.03 56.54 2.355 ;
      RECT 56.29 1.13 56.47 2.355 ;
      RECT 56.235 1.13 56.525 1.36 ;
      RECT 56.235 1.16 56.695 1.33 ;
      RECT 56.22 4.26 56.545 4.585 ;
      RECT 56.22 4.34 56.695 4.51 ;
      RECT 55.51 2.05 55.83 2.39 ;
      RECT 55.505 2.05 55.83 2.065 ;
      RECT 55.63 0.39 55.795 2.39 ;
      RECT 55.59 0.39 55.915 0.715 ;
      RECT 54.59 1.165 54.91 1.425 ;
      RECT 54.315 1.225 54.91 1.365 ;
      RECT 52.21 1.505 52.53 1.765 ;
      RECT 54.185 1.52 54.475 1.75 ;
      RECT 52.21 1.565 54.475 1.705 ;
      RECT 53.57 4.225 53.89 4.485 ;
      RECT 53.57 4.285 54.165 4.425 ;
      RECT 52.89 1.165 53.21 1.425 ;
      RECT 48.15 1.18 48.44 1.41 ;
      RECT 48.15 1.225 53.21 1.365 ;
      RECT 52.98 0.885 53.12 1.425 ;
      RECT 52.98 0.885 53.46 1.025 ;
      RECT 53.32 0.5 53.46 1.025 ;
      RECT 53.245 0.5 53.535 0.73 ;
      RECT 52.89 2.185 53.21 2.445 ;
      RECT 52.225 2.2 52.515 2.43 ;
      RECT 50.015 2.2 50.305 2.43 ;
      RECT 50.015 2.245 53.21 2.385 ;
      RECT 51.19 4.225 51.51 4.485 ;
      RECT 52.905 4.24 53.195 4.47 ;
      RECT 50.525 4.24 50.815 4.47 ;
      RECT 50.525 4.285 51.51 4.425 ;
      RECT 52.98 3.945 53.12 4.47 ;
      RECT 51.28 3.945 51.42 4.485 ;
      RECT 51.28 3.945 53.12 4.085 ;
      RECT 50.185 0.84 50.475 1.07 ;
      RECT 50.26 0.545 50.4 1.07 ;
      RECT 52.55 0.485 52.87 0.745 ;
      RECT 52.45 0.5 52.87 0.73 ;
      RECT 50.26 0.545 52.87 0.685 ;
      RECT 51.53 0.825 51.85 1.085 ;
      RECT 51.53 0.885 52.125 1.025 ;
      RECT 50.51 4.905 50.83 5.165 ;
      RECT 49.58 4.965 51.93 5.105 ;
      RECT 51.79 4.24 51.93 5.105 ;
      RECT 49.58 4.24 49.72 5.105 ;
      RECT 51.715 4.24 52.005 4.47 ;
      RECT 49.505 4.24 49.795 4.47 ;
      RECT 51.53 3.205 51.85 3.465 ;
      RECT 48.825 3.22 49.115 3.45 ;
      RECT 48.825 3.265 51.85 3.405 ;
      RECT 50.855 0.785 51.185 1.115 ;
      RECT 50.85 0.82 51.185 1.08 ;
      RECT 51.2 0.84 51.315 1.07 ;
      RECT 50.85 0.835 51.2 1.065 ;
      RECT 50.85 0.885 51.33 1.025 ;
      RECT 50.735 0.885 50.745 1.025 ;
      RECT 50.745 0.88 51.315 1.02 ;
      RECT 46.22 0.76 46.51 0.99 ;
      RECT 46.28 -0.72 46.45 0.99 ;
      RECT 46.25 -0.505 46.6 -0.155 ;
      RECT 46.22 -0.72 46.51 -0.49 ;
      RECT 46.22 6.16 46.51 6.39 ;
      RECT 46.28 4.68 46.45 6.39 ;
      RECT 46.22 4.68 46.51 4.91 ;
      RECT 45.81 1.13 46.14 1.36 ;
      RECT 45.81 1.16 46.31 1.33 ;
      RECT 45.81 0.79 46 1.36 ;
      RECT 45.23 0.76 45.52 0.99 ;
      RECT 45.23 0.79 46 0.96 ;
      RECT 45.29 -0.72 45.46 0.99 ;
      RECT 45.23 -0.72 45.52 -0.49 ;
      RECT 45.23 6.16 45.52 6.39 ;
      RECT 45.29 4.68 45.46 6.39 ;
      RECT 45.23 4.68 45.52 4.91 ;
      RECT 45.23 4.72 46.08 4.88 ;
      RECT 45.91 4.31 46.08 4.88 ;
      RECT 45.23 4.715 45.62 4.88 ;
      RECT 45.85 4.31 46.14 4.54 ;
      RECT 45.85 4.34 46.31 4.51 ;
      RECT 44.86 1.13 45.15 1.36 ;
      RECT 44.86 1.16 45.32 1.33 ;
      RECT 44.92 0.05 45.085 1.36 ;
      RECT 43.435 0.02 43.725 0.25 ;
      RECT 43.435 0.05 45.085 0.22 ;
      RECT 43.495 -0.72 43.665 0.25 ;
      RECT 43.435 -0.72 43.725 -0.49 ;
      RECT 43.435 6.16 43.725 6.39 ;
      RECT 43.495 5.42 43.665 6.39 ;
      RECT 43.495 5.515 45.085 5.685 ;
      RECT 44.915 4.31 45.085 5.685 ;
      RECT 43.435 5.42 43.725 5.65 ;
      RECT 44.86 4.31 45.15 4.54 ;
      RECT 44.86 4.34 45.32 4.51 ;
      RECT 43.865 0.36 44.215 0.71 ;
      RECT 43.695 0.42 44.215 0.59 ;
      RECT 43.89 5.05 44.215 5.375 ;
      RECT 43.865 5.05 44.215 5.28 ;
      RECT 43.695 5.08 44.215 5.25 ;
      RECT 43.09 0.76 43.41 1.08 ;
      RECT 43.06 0.76 43.41 0.99 ;
      RECT 42.775 0.79 43.41 0.96 ;
      RECT 43.09 4.675 43.41 5 ;
      RECT 43.06 4.68 43.41 4.91 ;
      RECT 42.89 4.71 43.41 4.88 ;
      RECT 42.045 2.03 42.37 2.355 ;
      RECT 42.12 1.13 42.3 2.355 ;
      RECT 42.065 1.13 42.355 1.36 ;
      RECT 42.065 1.16 42.525 1.33 ;
      RECT 42.05 4.26 42.375 4.585 ;
      RECT 42.05 4.34 42.525 4.51 ;
      RECT 41.34 2.05 41.66 2.39 ;
      RECT 41.335 2.05 41.66 2.065 ;
      RECT 41.46 0.39 41.625 2.39 ;
      RECT 41.42 0.39 41.745 0.715 ;
      RECT 40.42 1.165 40.74 1.425 ;
      RECT 40.145 1.225 40.74 1.365 ;
      RECT 38.04 1.505 38.36 1.765 ;
      RECT 40.015 1.52 40.305 1.75 ;
      RECT 38.04 1.565 40.305 1.705 ;
      RECT 39.4 4.225 39.72 4.485 ;
      RECT 39.4 4.285 39.995 4.425 ;
      RECT 38.72 1.165 39.04 1.425 ;
      RECT 33.98 1.18 34.27 1.41 ;
      RECT 33.98 1.225 39.04 1.365 ;
      RECT 38.81 0.885 38.95 1.425 ;
      RECT 38.81 0.885 39.29 1.025 ;
      RECT 39.15 0.5 39.29 1.025 ;
      RECT 39.075 0.5 39.365 0.73 ;
      RECT 38.72 2.185 39.04 2.445 ;
      RECT 38.055 2.2 38.345 2.43 ;
      RECT 35.845 2.2 36.135 2.43 ;
      RECT 35.845 2.245 39.04 2.385 ;
      RECT 37.02 4.225 37.34 4.485 ;
      RECT 38.735 4.24 39.025 4.47 ;
      RECT 36.355 4.24 36.645 4.47 ;
      RECT 36.355 4.285 37.34 4.425 ;
      RECT 38.81 3.945 38.95 4.47 ;
      RECT 37.11 3.945 37.25 4.485 ;
      RECT 37.11 3.945 38.95 4.085 ;
      RECT 36.015 0.84 36.305 1.07 ;
      RECT 36.09 0.545 36.23 1.07 ;
      RECT 38.38 0.485 38.7 0.745 ;
      RECT 38.28 0.5 38.7 0.73 ;
      RECT 36.09 0.545 38.7 0.685 ;
      RECT 37.36 0.825 37.68 1.085 ;
      RECT 37.36 0.885 37.955 1.025 ;
      RECT 36.34 4.905 36.66 5.165 ;
      RECT 35.41 4.965 37.76 5.105 ;
      RECT 37.62 4.24 37.76 5.105 ;
      RECT 35.41 4.24 35.55 5.105 ;
      RECT 37.545 4.24 37.835 4.47 ;
      RECT 35.335 4.24 35.625 4.47 ;
      RECT 37.36 3.205 37.68 3.465 ;
      RECT 34.655 3.22 34.945 3.45 ;
      RECT 34.655 3.265 37.68 3.405 ;
      RECT 36.685 0.785 37.015 1.115 ;
      RECT 36.68 0.82 37.015 1.08 ;
      RECT 37.03 0.84 37.145 1.07 ;
      RECT 36.68 0.835 37.03 1.065 ;
      RECT 36.68 0.885 37.16 1.025 ;
      RECT 36.565 0.885 36.575 1.025 ;
      RECT 36.575 0.88 37.145 1.02 ;
      RECT 32.045 0.76 32.335 0.99 ;
      RECT 32.105 -0.72 32.275 0.99 ;
      RECT 32.075 -0.52 32.425 -0.17 ;
      RECT 32.045 -0.72 32.335 -0.49 ;
      RECT 32.045 6.16 32.335 6.39 ;
      RECT 32.105 4.68 32.275 6.39 ;
      RECT 32.045 4.68 32.335 4.91 ;
      RECT 31.635 1.13 31.965 1.36 ;
      RECT 31.635 1.16 32.135 1.33 ;
      RECT 31.635 0.79 31.825 1.36 ;
      RECT 31.055 0.76 31.345 0.99 ;
      RECT 31.055 0.79 31.825 0.96 ;
      RECT 31.115 -0.72 31.285 0.99 ;
      RECT 31.055 -0.72 31.345 -0.49 ;
      RECT 31.055 6.16 31.345 6.39 ;
      RECT 31.115 4.68 31.285 6.39 ;
      RECT 31.055 4.68 31.345 4.91 ;
      RECT 31.055 4.72 31.905 4.88 ;
      RECT 31.735 4.31 31.905 4.88 ;
      RECT 31.055 4.715 31.445 4.88 ;
      RECT 31.675 4.31 31.965 4.54 ;
      RECT 31.675 4.34 32.135 4.51 ;
      RECT 30.685 1.13 30.975 1.36 ;
      RECT 30.685 1.16 31.145 1.33 ;
      RECT 30.745 0.05 30.91 1.36 ;
      RECT 29.26 0.02 29.55 0.25 ;
      RECT 29.26 0.05 30.91 0.22 ;
      RECT 29.32 -0.72 29.49 0.25 ;
      RECT 29.26 -0.72 29.55 -0.49 ;
      RECT 29.26 6.16 29.55 6.39 ;
      RECT 29.32 5.42 29.49 6.39 ;
      RECT 29.32 5.515 30.91 5.685 ;
      RECT 30.74 4.31 30.91 5.685 ;
      RECT 29.26 5.42 29.55 5.65 ;
      RECT 30.685 4.31 30.975 4.54 ;
      RECT 30.685 4.34 31.145 4.51 ;
      RECT 29.69 0.36 30.04 0.71 ;
      RECT 29.52 0.42 30.04 0.59 ;
      RECT 29.715 5.05 30.04 5.375 ;
      RECT 29.69 5.05 30.04 5.28 ;
      RECT 29.52 5.08 30.04 5.25 ;
      RECT 28.915 0.76 29.235 1.08 ;
      RECT 28.885 0.76 29.235 0.99 ;
      RECT 28.6 0.79 29.235 0.96 ;
      RECT 28.915 4.675 29.235 5 ;
      RECT 28.885 4.68 29.235 4.91 ;
      RECT 28.715 4.71 29.235 4.88 ;
      RECT 27.87 2.03 28.195 2.355 ;
      RECT 27.945 1.13 28.125 2.355 ;
      RECT 27.89 1.13 28.18 1.36 ;
      RECT 27.89 1.16 28.35 1.33 ;
      RECT 27.875 4.26 28.2 4.585 ;
      RECT 27.875 4.34 28.35 4.51 ;
      RECT 27.165 2.05 27.485 2.39 ;
      RECT 27.16 2.05 27.485 2.065 ;
      RECT 27.285 0.39 27.45 2.39 ;
      RECT 27.245 0.39 27.57 0.715 ;
      RECT 26.245 1.165 26.565 1.425 ;
      RECT 25.97 1.225 26.565 1.365 ;
      RECT 23.865 1.505 24.185 1.765 ;
      RECT 25.84 1.52 26.13 1.75 ;
      RECT 23.865 1.565 26.13 1.705 ;
      RECT 25.225 4.225 25.545 4.485 ;
      RECT 25.225 4.285 25.82 4.425 ;
      RECT 24.545 1.165 24.865 1.425 ;
      RECT 19.805 1.18 20.095 1.41 ;
      RECT 19.805 1.225 24.865 1.365 ;
      RECT 24.635 0.885 24.775 1.425 ;
      RECT 24.635 0.885 25.115 1.025 ;
      RECT 24.975 0.5 25.115 1.025 ;
      RECT 24.9 0.5 25.19 0.73 ;
      RECT 24.545 2.185 24.865 2.445 ;
      RECT 23.88 2.2 24.17 2.43 ;
      RECT 21.67 2.2 21.96 2.43 ;
      RECT 21.67 2.245 24.865 2.385 ;
      RECT 22.845 4.225 23.165 4.485 ;
      RECT 24.56 4.24 24.85 4.47 ;
      RECT 22.18 4.24 22.47 4.47 ;
      RECT 22.18 4.285 23.165 4.425 ;
      RECT 24.635 3.945 24.775 4.47 ;
      RECT 22.935 3.945 23.075 4.485 ;
      RECT 22.935 3.945 24.775 4.085 ;
      RECT 21.84 0.84 22.13 1.07 ;
      RECT 21.915 0.545 22.055 1.07 ;
      RECT 24.205 0.485 24.525 0.745 ;
      RECT 24.105 0.5 24.525 0.73 ;
      RECT 21.915 0.545 24.525 0.685 ;
      RECT 23.185 0.825 23.505 1.085 ;
      RECT 23.185 0.885 23.78 1.025 ;
      RECT 22.165 4.905 22.485 5.165 ;
      RECT 21.235 4.965 23.585 5.105 ;
      RECT 23.445 4.24 23.585 5.105 ;
      RECT 21.235 4.24 21.375 5.105 ;
      RECT 23.37 4.24 23.66 4.47 ;
      RECT 21.16 4.24 21.45 4.47 ;
      RECT 23.185 3.205 23.505 3.465 ;
      RECT 20.48 3.22 20.77 3.45 ;
      RECT 20.48 3.265 23.505 3.405 ;
      RECT 22.51 0.785 22.84 1.115 ;
      RECT 22.505 0.82 22.84 1.08 ;
      RECT 22.855 0.84 22.97 1.07 ;
      RECT 22.505 0.835 22.855 1.065 ;
      RECT 22.505 0.885 22.985 1.025 ;
      RECT 22.39 0.885 22.4 1.025 ;
      RECT 22.4 0.88 22.97 1.02 ;
      RECT 17.875 0.76 18.165 0.99 ;
      RECT 17.935 -0.72 18.105 0.99 ;
      RECT 17.91 -0.51 18.26 -0.16 ;
      RECT 17.875 -0.72 18.165 -0.49 ;
      RECT 17.875 -0.515 18.17 -0.49 ;
      RECT 17.875 6.16 18.165 6.39 ;
      RECT 17.935 4.68 18.105 6.39 ;
      RECT 17.875 4.68 18.165 4.91 ;
      RECT 17.465 1.13 17.795 1.36 ;
      RECT 17.465 1.16 17.965 1.33 ;
      RECT 17.465 0.79 17.655 1.36 ;
      RECT 16.885 0.76 17.175 0.99 ;
      RECT 16.885 0.79 17.655 0.96 ;
      RECT 16.945 -0.72 17.115 0.99 ;
      RECT 16.885 -0.72 17.175 -0.49 ;
      RECT 16.885 6.16 17.175 6.39 ;
      RECT 16.945 4.68 17.115 6.39 ;
      RECT 16.885 4.68 17.175 4.91 ;
      RECT 16.885 4.72 17.735 4.88 ;
      RECT 17.565 4.31 17.735 4.88 ;
      RECT 16.885 4.715 17.275 4.88 ;
      RECT 17.505 4.31 17.795 4.54 ;
      RECT 17.505 4.34 17.965 4.51 ;
      RECT 16.515 1.13 16.805 1.36 ;
      RECT 16.515 1.16 16.975 1.33 ;
      RECT 16.575 0.05 16.74 1.36 ;
      RECT 15.09 0.02 15.38 0.25 ;
      RECT 15.09 0.05 16.74 0.22 ;
      RECT 15.15 -0.72 15.32 0.25 ;
      RECT 15.09 -0.72 15.38 -0.49 ;
      RECT 15.09 6.16 15.38 6.39 ;
      RECT 15.15 5.42 15.32 6.39 ;
      RECT 15.15 5.515 16.74 5.685 ;
      RECT 16.57 4.31 16.74 5.685 ;
      RECT 15.09 5.42 15.38 5.65 ;
      RECT 16.515 4.31 16.805 4.54 ;
      RECT 16.515 4.34 16.975 4.51 ;
      RECT 15.52 0.36 15.87 0.71 ;
      RECT 15.35 0.42 15.87 0.59 ;
      RECT 15.545 5.05 15.87 5.375 ;
      RECT 15.52 5.05 15.87 5.28 ;
      RECT 15.35 5.08 15.87 5.25 ;
      RECT 14.745 0.76 15.065 1.08 ;
      RECT 14.715 0.76 15.065 0.99 ;
      RECT 14.43 0.79 15.065 0.96 ;
      RECT 14.745 4.675 15.065 5 ;
      RECT 14.715 4.68 15.065 4.91 ;
      RECT 14.545 4.71 15.065 4.88 ;
      RECT 13.7 2.03 14.025 2.355 ;
      RECT 13.775 1.13 13.955 2.355 ;
      RECT 13.72 1.13 14.01 1.36 ;
      RECT 13.72 1.16 14.18 1.33 ;
      RECT 13.705 4.26 14.03 4.585 ;
      RECT 13.705 4.34 14.18 4.51 ;
      RECT 12.995 2.05 13.315 2.39 ;
      RECT 12.99 2.05 13.315 2.065 ;
      RECT 13.115 0.39 13.28 2.39 ;
      RECT 13.075 0.39 13.4 0.715 ;
      RECT 12.075 1.165 12.395 1.425 ;
      RECT 11.8 1.225 12.395 1.365 ;
      RECT 9.695 1.505 10.015 1.765 ;
      RECT 11.67 1.52 11.96 1.75 ;
      RECT 9.695 1.565 11.96 1.705 ;
      RECT 11.055 4.225 11.375 4.485 ;
      RECT 11.055 4.285 11.65 4.425 ;
      RECT 10.375 1.165 10.695 1.425 ;
      RECT 5.635 1.18 5.925 1.41 ;
      RECT 5.635 1.225 10.695 1.365 ;
      RECT 10.465 0.885 10.605 1.425 ;
      RECT 10.465 0.885 10.945 1.025 ;
      RECT 10.805 0.5 10.945 1.025 ;
      RECT 10.73 0.5 11.02 0.73 ;
      RECT 10.375 2.185 10.695 2.445 ;
      RECT 9.71 2.2 10 2.43 ;
      RECT 7.5 2.2 7.79 2.43 ;
      RECT 7.5 2.245 10.695 2.385 ;
      RECT 8.675 4.225 8.995 4.485 ;
      RECT 10.39 4.24 10.68 4.47 ;
      RECT 8.01 4.24 8.3 4.47 ;
      RECT 8.01 4.285 8.995 4.425 ;
      RECT 10.465 3.945 10.605 4.47 ;
      RECT 8.765 3.945 8.905 4.485 ;
      RECT 8.765 3.945 10.605 4.085 ;
      RECT 7.67 0.84 7.96 1.07 ;
      RECT 7.745 0.545 7.885 1.07 ;
      RECT 10.035 0.485 10.355 0.745 ;
      RECT 9.935 0.5 10.355 0.73 ;
      RECT 7.745 0.545 10.355 0.685 ;
      RECT 9.015 0.825 9.335 1.085 ;
      RECT 9.015 0.885 9.61 1.025 ;
      RECT 7.995 4.905 8.315 5.165 ;
      RECT 7.065 4.965 9.415 5.105 ;
      RECT 9.275 4.24 9.415 5.105 ;
      RECT 7.065 4.24 7.205 5.105 ;
      RECT 9.2 4.24 9.49 4.47 ;
      RECT 6.99 4.24 7.28 4.47 ;
      RECT 9.015 3.205 9.335 3.465 ;
      RECT 6.31 3.22 6.6 3.45 ;
      RECT 6.31 3.265 9.335 3.405 ;
      RECT 8.34 0.785 8.67 1.115 ;
      RECT 8.335 0.82 8.67 1.08 ;
      RECT 8.685 0.84 8.8 1.07 ;
      RECT 8.335 0.835 8.685 1.065 ;
      RECT 8.335 0.885 8.815 1.025 ;
      RECT 8.22 0.885 8.23 1.025 ;
      RECT 8.23 0.88 8.8 1.02 ;
      RECT 69.18 1.58 69.505 1.905 ;
      RECT 68.44 3.205 69.085 3.465 ;
      RECT 66.385 4.225 66.705 4.485 ;
      RECT 55.005 1.58 55.33 1.905 ;
      RECT 54.265 3.205 54.91 3.465 ;
      RECT 52.21 4.225 52.53 4.485 ;
      RECT 40.835 1.58 41.16 1.905 ;
      RECT 40.095 3.205 40.74 3.465 ;
      RECT 38.04 4.225 38.36 4.485 ;
      RECT 26.66 1.58 26.985 1.905 ;
      RECT 25.92 3.205 26.565 3.465 ;
      RECT 23.865 4.225 24.185 4.485 ;
      RECT 12.49 1.58 12.815 1.905 ;
      RECT 11.75 3.205 12.395 3.465 ;
      RECT 9.695 4.225 10.015 4.485 ;
    LAYER mcon ;
      RECT 74.625 -0.69 74.795 -0.52 ;
      RECT 74.625 0.79 74.795 0.96 ;
      RECT 74.625 4.71 74.795 4.88 ;
      RECT 74.625 6.19 74.795 6.36 ;
      RECT 74.275 -1.5 74.445 -1.33 ;
      RECT 74.275 2.56 74.445 2.73 ;
      RECT 74.275 2.94 74.445 3.11 ;
      RECT 74.275 7 74.445 7.17 ;
      RECT 74.255 1.16 74.425 1.33 ;
      RECT 74.255 4.34 74.425 4.51 ;
      RECT 73.635 -0.69 73.805 -0.52 ;
      RECT 73.635 0.79 73.805 0.96 ;
      RECT 73.635 4.71 73.805 4.88 ;
      RECT 73.635 6.19 73.805 6.36 ;
      RECT 73.285 -1.5 73.455 -1.33 ;
      RECT 73.285 2.56 73.455 2.73 ;
      RECT 73.285 2.94 73.455 3.11 ;
      RECT 73.285 7 73.455 7.17 ;
      RECT 73.265 1.16 73.435 1.33 ;
      RECT 73.265 4.34 73.435 4.51 ;
      RECT 72.58 -1.5 72.75 -1.33 ;
      RECT 72.58 2.56 72.75 2.73 ;
      RECT 72.58 2.94 72.75 3.11 ;
      RECT 72.58 7 72.75 7.17 ;
      RECT 72.27 0.42 72.44 0.59 ;
      RECT 72.27 5.08 72.44 5.25 ;
      RECT 71.9 -1.5 72.07 -1.33 ;
      RECT 71.9 7 72.07 7.17 ;
      RECT 71.84 -0.69 72.01 -0.52 ;
      RECT 71.84 0.05 72.01 0.22 ;
      RECT 71.84 5.45 72.01 5.62 ;
      RECT 71.84 6.19 72.01 6.36 ;
      RECT 71.465 0.79 71.635 0.96 ;
      RECT 71.465 4.71 71.635 4.88 ;
      RECT 71.22 -1.5 71.39 -1.33 ;
      RECT 71.22 7 71.39 7.17 ;
      RECT 70.54 -1.5 70.71 -1.33 ;
      RECT 70.54 7 70.71 7.17 ;
      RECT 70.47 1.16 70.64 1.33 ;
      RECT 70.47 4.34 70.64 4.51 ;
      RECT 68.88 0.02 69.05 0.19 ;
      RECT 68.88 2.74 69.05 2.91 ;
      RECT 68.88 5.46 69.05 5.63 ;
      RECT 68.84 1.21 69.01 1.38 ;
      RECT 68.5 3.25 68.67 3.42 ;
      RECT 68.42 0.02 68.59 0.19 ;
      RECT 68.42 1.55 68.59 1.72 ;
      RECT 68.42 2.74 68.59 2.91 ;
      RECT 68.42 5.46 68.59 5.63 ;
      RECT 67.96 0.02 68.13 0.19 ;
      RECT 67.96 2.74 68.13 2.91 ;
      RECT 67.96 5.46 68.13 5.63 ;
      RECT 67.82 4.27 67.99 4.44 ;
      RECT 67.5 0.02 67.67 0.19 ;
      RECT 67.5 2.74 67.67 2.91 ;
      RECT 67.5 5.46 67.67 5.63 ;
      RECT 67.48 0.53 67.65 0.7 ;
      RECT 67.14 4.27 67.31 4.44 ;
      RECT 67.04 0.02 67.21 0.19 ;
      RECT 67.04 2.74 67.21 2.91 ;
      RECT 67.04 5.46 67.21 5.63 ;
      RECT 66.685 0.53 66.855 0.7 ;
      RECT 66.58 0.02 66.75 0.19 ;
      RECT 66.58 2.74 66.75 2.91 ;
      RECT 66.58 5.46 66.75 5.63 ;
      RECT 66.46 2.23 66.63 2.4 ;
      RECT 66.46 4.27 66.63 4.44 ;
      RECT 66.12 0.02 66.29 0.19 ;
      RECT 66.12 2.74 66.29 2.91 ;
      RECT 66.12 5.46 66.29 5.63 ;
      RECT 65.95 4.27 66.12 4.44 ;
      RECT 65.78 0.87 65.95 1.04 ;
      RECT 65.66 0.02 65.83 0.19 ;
      RECT 65.66 2.74 65.83 2.91 ;
      RECT 65.66 5.46 65.83 5.63 ;
      RECT 65.2 0.02 65.37 0.19 ;
      RECT 65.2 2.74 65.37 2.91 ;
      RECT 65.2 5.46 65.37 5.63 ;
      RECT 64.76 4.27 64.93 4.44 ;
      RECT 64.74 0.02 64.91 0.19 ;
      RECT 64.74 2.74 64.91 2.91 ;
      RECT 64.74 5.46 64.91 5.63 ;
      RECT 64.42 0.87 64.59 1.04 ;
      RECT 64.28 0.02 64.45 0.19 ;
      RECT 64.28 2.74 64.45 2.91 ;
      RECT 64.28 5.46 64.45 5.63 ;
      RECT 64.25 2.23 64.42 2.4 ;
      RECT 63.82 0.02 63.99 0.19 ;
      RECT 63.82 2.74 63.99 2.91 ;
      RECT 63.82 5.46 63.99 5.63 ;
      RECT 63.74 4.27 63.91 4.44 ;
      RECT 63.36 0.02 63.53 0.19 ;
      RECT 63.36 2.74 63.53 2.91 ;
      RECT 63.36 5.46 63.53 5.63 ;
      RECT 63.06 3.25 63.23 3.42 ;
      RECT 62.9 0.02 63.07 0.19 ;
      RECT 62.9 2.74 63.07 2.91 ;
      RECT 62.9 5.46 63.07 5.63 ;
      RECT 62.44 0.02 62.61 0.19 ;
      RECT 62.44 2.74 62.61 2.91 ;
      RECT 62.44 5.46 62.61 5.63 ;
      RECT 62.385 1.21 62.555 1.38 ;
      RECT 60.45 -0.69 60.62 -0.52 ;
      RECT 60.45 0.79 60.62 0.96 ;
      RECT 60.45 4.71 60.62 4.88 ;
      RECT 60.45 6.19 60.62 6.36 ;
      RECT 60.1 -1.5 60.27 -1.33 ;
      RECT 60.1 2.56 60.27 2.73 ;
      RECT 60.1 2.94 60.27 3.11 ;
      RECT 60.1 7 60.27 7.17 ;
      RECT 60.08 1.16 60.25 1.33 ;
      RECT 60.08 4.34 60.25 4.51 ;
      RECT 59.46 -0.69 59.63 -0.52 ;
      RECT 59.46 0.79 59.63 0.96 ;
      RECT 59.46 4.71 59.63 4.88 ;
      RECT 59.46 6.19 59.63 6.36 ;
      RECT 59.11 -1.5 59.28 -1.33 ;
      RECT 59.11 2.56 59.28 2.73 ;
      RECT 59.11 2.94 59.28 3.11 ;
      RECT 59.11 7 59.28 7.17 ;
      RECT 59.09 1.16 59.26 1.33 ;
      RECT 59.09 4.34 59.26 4.51 ;
      RECT 58.405 -1.5 58.575 -1.33 ;
      RECT 58.405 2.56 58.575 2.73 ;
      RECT 58.405 2.94 58.575 3.11 ;
      RECT 58.405 7 58.575 7.17 ;
      RECT 58.095 0.42 58.265 0.59 ;
      RECT 58.095 5.08 58.265 5.25 ;
      RECT 57.725 -1.5 57.895 -1.33 ;
      RECT 57.725 7 57.895 7.17 ;
      RECT 57.665 -0.69 57.835 -0.52 ;
      RECT 57.665 0.05 57.835 0.22 ;
      RECT 57.665 5.45 57.835 5.62 ;
      RECT 57.665 6.19 57.835 6.36 ;
      RECT 57.29 0.79 57.46 0.96 ;
      RECT 57.29 4.71 57.46 4.88 ;
      RECT 57.045 -1.5 57.215 -1.33 ;
      RECT 57.045 7 57.215 7.17 ;
      RECT 56.365 -1.5 56.535 -1.33 ;
      RECT 56.365 7 56.535 7.17 ;
      RECT 56.295 1.16 56.465 1.33 ;
      RECT 56.295 4.34 56.465 4.51 ;
      RECT 54.705 0.02 54.875 0.19 ;
      RECT 54.705 2.74 54.875 2.91 ;
      RECT 54.705 5.46 54.875 5.63 ;
      RECT 54.665 1.21 54.835 1.38 ;
      RECT 54.325 3.25 54.495 3.42 ;
      RECT 54.245 0.02 54.415 0.19 ;
      RECT 54.245 1.55 54.415 1.72 ;
      RECT 54.245 2.74 54.415 2.91 ;
      RECT 54.245 5.46 54.415 5.63 ;
      RECT 53.785 0.02 53.955 0.19 ;
      RECT 53.785 2.74 53.955 2.91 ;
      RECT 53.785 5.46 53.955 5.63 ;
      RECT 53.645 4.27 53.815 4.44 ;
      RECT 53.325 0.02 53.495 0.19 ;
      RECT 53.325 2.74 53.495 2.91 ;
      RECT 53.325 5.46 53.495 5.63 ;
      RECT 53.305 0.53 53.475 0.7 ;
      RECT 52.965 4.27 53.135 4.44 ;
      RECT 52.865 0.02 53.035 0.19 ;
      RECT 52.865 2.74 53.035 2.91 ;
      RECT 52.865 5.46 53.035 5.63 ;
      RECT 52.51 0.53 52.68 0.7 ;
      RECT 52.405 0.02 52.575 0.19 ;
      RECT 52.405 2.74 52.575 2.91 ;
      RECT 52.405 5.46 52.575 5.63 ;
      RECT 52.285 2.23 52.455 2.4 ;
      RECT 52.285 4.27 52.455 4.44 ;
      RECT 51.945 0.02 52.115 0.19 ;
      RECT 51.945 2.74 52.115 2.91 ;
      RECT 51.945 5.46 52.115 5.63 ;
      RECT 51.775 4.27 51.945 4.44 ;
      RECT 51.605 0.87 51.775 1.04 ;
      RECT 51.485 0.02 51.655 0.19 ;
      RECT 51.485 2.74 51.655 2.91 ;
      RECT 51.485 5.46 51.655 5.63 ;
      RECT 51.025 0.02 51.195 0.19 ;
      RECT 51.025 2.74 51.195 2.91 ;
      RECT 51.025 5.46 51.195 5.63 ;
      RECT 50.585 4.27 50.755 4.44 ;
      RECT 50.565 0.02 50.735 0.19 ;
      RECT 50.565 2.74 50.735 2.91 ;
      RECT 50.565 5.46 50.735 5.63 ;
      RECT 50.245 0.87 50.415 1.04 ;
      RECT 50.105 0.02 50.275 0.19 ;
      RECT 50.105 2.74 50.275 2.91 ;
      RECT 50.105 5.46 50.275 5.63 ;
      RECT 50.075 2.23 50.245 2.4 ;
      RECT 49.645 0.02 49.815 0.19 ;
      RECT 49.645 2.74 49.815 2.91 ;
      RECT 49.645 5.46 49.815 5.63 ;
      RECT 49.565 4.27 49.735 4.44 ;
      RECT 49.185 0.02 49.355 0.19 ;
      RECT 49.185 2.74 49.355 2.91 ;
      RECT 49.185 5.46 49.355 5.63 ;
      RECT 48.885 3.25 49.055 3.42 ;
      RECT 48.725 0.02 48.895 0.19 ;
      RECT 48.725 2.74 48.895 2.91 ;
      RECT 48.725 5.46 48.895 5.63 ;
      RECT 48.265 0.02 48.435 0.19 ;
      RECT 48.265 2.74 48.435 2.91 ;
      RECT 48.265 5.46 48.435 5.63 ;
      RECT 48.21 1.21 48.38 1.38 ;
      RECT 46.28 -0.69 46.45 -0.52 ;
      RECT 46.28 0.79 46.45 0.96 ;
      RECT 46.28 4.71 46.45 4.88 ;
      RECT 46.28 6.19 46.45 6.36 ;
      RECT 45.93 -1.5 46.1 -1.33 ;
      RECT 45.93 2.56 46.1 2.73 ;
      RECT 45.93 2.94 46.1 3.11 ;
      RECT 45.93 7 46.1 7.17 ;
      RECT 45.91 1.16 46.08 1.33 ;
      RECT 45.91 4.34 46.08 4.51 ;
      RECT 45.29 -0.69 45.46 -0.52 ;
      RECT 45.29 0.79 45.46 0.96 ;
      RECT 45.29 4.71 45.46 4.88 ;
      RECT 45.29 6.19 45.46 6.36 ;
      RECT 44.94 -1.5 45.11 -1.33 ;
      RECT 44.94 2.56 45.11 2.73 ;
      RECT 44.94 2.94 45.11 3.11 ;
      RECT 44.94 7 45.11 7.17 ;
      RECT 44.92 1.16 45.09 1.33 ;
      RECT 44.92 4.34 45.09 4.51 ;
      RECT 44.235 -1.5 44.405 -1.33 ;
      RECT 44.235 2.56 44.405 2.73 ;
      RECT 44.235 2.94 44.405 3.11 ;
      RECT 44.235 7 44.405 7.17 ;
      RECT 43.925 0.42 44.095 0.59 ;
      RECT 43.925 5.08 44.095 5.25 ;
      RECT 43.555 -1.5 43.725 -1.33 ;
      RECT 43.555 7 43.725 7.17 ;
      RECT 43.495 -0.69 43.665 -0.52 ;
      RECT 43.495 0.05 43.665 0.22 ;
      RECT 43.495 5.45 43.665 5.62 ;
      RECT 43.495 6.19 43.665 6.36 ;
      RECT 43.12 0.79 43.29 0.96 ;
      RECT 43.12 4.71 43.29 4.88 ;
      RECT 42.875 -1.5 43.045 -1.33 ;
      RECT 42.875 7 43.045 7.17 ;
      RECT 42.195 -1.5 42.365 -1.33 ;
      RECT 42.195 7 42.365 7.17 ;
      RECT 42.125 1.16 42.295 1.33 ;
      RECT 42.125 4.34 42.295 4.51 ;
      RECT 40.535 0.02 40.705 0.19 ;
      RECT 40.535 2.74 40.705 2.91 ;
      RECT 40.535 5.46 40.705 5.63 ;
      RECT 40.495 1.21 40.665 1.38 ;
      RECT 40.155 3.25 40.325 3.42 ;
      RECT 40.075 0.02 40.245 0.19 ;
      RECT 40.075 1.55 40.245 1.72 ;
      RECT 40.075 2.74 40.245 2.91 ;
      RECT 40.075 5.46 40.245 5.63 ;
      RECT 39.615 0.02 39.785 0.19 ;
      RECT 39.615 2.74 39.785 2.91 ;
      RECT 39.615 5.46 39.785 5.63 ;
      RECT 39.475 4.27 39.645 4.44 ;
      RECT 39.155 0.02 39.325 0.19 ;
      RECT 39.155 2.74 39.325 2.91 ;
      RECT 39.155 5.46 39.325 5.63 ;
      RECT 39.135 0.53 39.305 0.7 ;
      RECT 38.795 4.27 38.965 4.44 ;
      RECT 38.695 0.02 38.865 0.19 ;
      RECT 38.695 2.74 38.865 2.91 ;
      RECT 38.695 5.46 38.865 5.63 ;
      RECT 38.34 0.53 38.51 0.7 ;
      RECT 38.235 0.02 38.405 0.19 ;
      RECT 38.235 2.74 38.405 2.91 ;
      RECT 38.235 5.46 38.405 5.63 ;
      RECT 38.115 2.23 38.285 2.4 ;
      RECT 38.115 4.27 38.285 4.44 ;
      RECT 37.775 0.02 37.945 0.19 ;
      RECT 37.775 2.74 37.945 2.91 ;
      RECT 37.775 5.46 37.945 5.63 ;
      RECT 37.605 4.27 37.775 4.44 ;
      RECT 37.435 0.87 37.605 1.04 ;
      RECT 37.315 0.02 37.485 0.19 ;
      RECT 37.315 2.74 37.485 2.91 ;
      RECT 37.315 5.46 37.485 5.63 ;
      RECT 36.855 0.02 37.025 0.19 ;
      RECT 36.855 2.74 37.025 2.91 ;
      RECT 36.855 5.46 37.025 5.63 ;
      RECT 36.415 4.27 36.585 4.44 ;
      RECT 36.395 0.02 36.565 0.19 ;
      RECT 36.395 2.74 36.565 2.91 ;
      RECT 36.395 5.46 36.565 5.63 ;
      RECT 36.075 0.87 36.245 1.04 ;
      RECT 35.935 0.02 36.105 0.19 ;
      RECT 35.935 2.74 36.105 2.91 ;
      RECT 35.935 5.46 36.105 5.63 ;
      RECT 35.905 2.23 36.075 2.4 ;
      RECT 35.475 0.02 35.645 0.19 ;
      RECT 35.475 2.74 35.645 2.91 ;
      RECT 35.475 5.46 35.645 5.63 ;
      RECT 35.395 4.27 35.565 4.44 ;
      RECT 35.015 0.02 35.185 0.19 ;
      RECT 35.015 2.74 35.185 2.91 ;
      RECT 35.015 5.46 35.185 5.63 ;
      RECT 34.715 3.25 34.885 3.42 ;
      RECT 34.555 0.02 34.725 0.19 ;
      RECT 34.555 2.74 34.725 2.91 ;
      RECT 34.555 5.46 34.725 5.63 ;
      RECT 34.095 0.02 34.265 0.19 ;
      RECT 34.095 2.74 34.265 2.91 ;
      RECT 34.095 5.46 34.265 5.63 ;
      RECT 34.04 1.21 34.21 1.38 ;
      RECT 32.105 -0.69 32.275 -0.52 ;
      RECT 32.105 0.79 32.275 0.96 ;
      RECT 32.105 4.71 32.275 4.88 ;
      RECT 32.105 6.19 32.275 6.36 ;
      RECT 31.755 -1.5 31.925 -1.33 ;
      RECT 31.755 2.56 31.925 2.73 ;
      RECT 31.755 2.94 31.925 3.11 ;
      RECT 31.755 7 31.925 7.17 ;
      RECT 31.735 1.16 31.905 1.33 ;
      RECT 31.735 4.34 31.905 4.51 ;
      RECT 31.115 -0.69 31.285 -0.52 ;
      RECT 31.115 0.79 31.285 0.96 ;
      RECT 31.115 4.71 31.285 4.88 ;
      RECT 31.115 6.19 31.285 6.36 ;
      RECT 30.765 -1.5 30.935 -1.33 ;
      RECT 30.765 2.56 30.935 2.73 ;
      RECT 30.765 2.94 30.935 3.11 ;
      RECT 30.765 7 30.935 7.17 ;
      RECT 30.745 1.16 30.915 1.33 ;
      RECT 30.745 4.34 30.915 4.51 ;
      RECT 30.06 -1.5 30.23 -1.33 ;
      RECT 30.06 2.56 30.23 2.73 ;
      RECT 30.06 2.94 30.23 3.11 ;
      RECT 30.06 7 30.23 7.17 ;
      RECT 29.75 0.42 29.92 0.59 ;
      RECT 29.75 5.08 29.92 5.25 ;
      RECT 29.38 -1.5 29.55 -1.33 ;
      RECT 29.38 7 29.55 7.17 ;
      RECT 29.32 -0.69 29.49 -0.52 ;
      RECT 29.32 0.05 29.49 0.22 ;
      RECT 29.32 5.45 29.49 5.62 ;
      RECT 29.32 6.19 29.49 6.36 ;
      RECT 28.945 0.79 29.115 0.96 ;
      RECT 28.945 4.71 29.115 4.88 ;
      RECT 28.7 -1.5 28.87 -1.33 ;
      RECT 28.7 7 28.87 7.17 ;
      RECT 28.02 -1.5 28.19 -1.33 ;
      RECT 28.02 7 28.19 7.17 ;
      RECT 27.95 1.16 28.12 1.33 ;
      RECT 27.95 4.34 28.12 4.51 ;
      RECT 26.36 0.02 26.53 0.19 ;
      RECT 26.36 2.74 26.53 2.91 ;
      RECT 26.36 5.46 26.53 5.63 ;
      RECT 26.32 1.21 26.49 1.38 ;
      RECT 25.98 3.25 26.15 3.42 ;
      RECT 25.9 0.02 26.07 0.19 ;
      RECT 25.9 1.55 26.07 1.72 ;
      RECT 25.9 2.74 26.07 2.91 ;
      RECT 25.9 5.46 26.07 5.63 ;
      RECT 25.44 0.02 25.61 0.19 ;
      RECT 25.44 2.74 25.61 2.91 ;
      RECT 25.44 5.46 25.61 5.63 ;
      RECT 25.3 4.27 25.47 4.44 ;
      RECT 24.98 0.02 25.15 0.19 ;
      RECT 24.98 2.74 25.15 2.91 ;
      RECT 24.98 5.46 25.15 5.63 ;
      RECT 24.96 0.53 25.13 0.7 ;
      RECT 24.62 4.27 24.79 4.44 ;
      RECT 24.52 0.02 24.69 0.19 ;
      RECT 24.52 2.74 24.69 2.91 ;
      RECT 24.52 5.46 24.69 5.63 ;
      RECT 24.165 0.53 24.335 0.7 ;
      RECT 24.06 0.02 24.23 0.19 ;
      RECT 24.06 2.74 24.23 2.91 ;
      RECT 24.06 5.46 24.23 5.63 ;
      RECT 23.94 2.23 24.11 2.4 ;
      RECT 23.94 4.27 24.11 4.44 ;
      RECT 23.6 0.02 23.77 0.19 ;
      RECT 23.6 2.74 23.77 2.91 ;
      RECT 23.6 5.46 23.77 5.63 ;
      RECT 23.43 4.27 23.6 4.44 ;
      RECT 23.26 0.87 23.43 1.04 ;
      RECT 23.14 0.02 23.31 0.19 ;
      RECT 23.14 2.74 23.31 2.91 ;
      RECT 23.14 5.46 23.31 5.63 ;
      RECT 22.68 0.02 22.85 0.19 ;
      RECT 22.68 2.74 22.85 2.91 ;
      RECT 22.68 5.46 22.85 5.63 ;
      RECT 22.24 4.27 22.41 4.44 ;
      RECT 22.22 0.02 22.39 0.19 ;
      RECT 22.22 2.74 22.39 2.91 ;
      RECT 22.22 5.46 22.39 5.63 ;
      RECT 21.9 0.87 22.07 1.04 ;
      RECT 21.76 0.02 21.93 0.19 ;
      RECT 21.76 2.74 21.93 2.91 ;
      RECT 21.76 5.46 21.93 5.63 ;
      RECT 21.73 2.23 21.9 2.4 ;
      RECT 21.3 0.02 21.47 0.19 ;
      RECT 21.3 2.74 21.47 2.91 ;
      RECT 21.3 5.46 21.47 5.63 ;
      RECT 21.22 4.27 21.39 4.44 ;
      RECT 20.84 0.02 21.01 0.19 ;
      RECT 20.84 2.74 21.01 2.91 ;
      RECT 20.84 5.46 21.01 5.63 ;
      RECT 20.54 3.25 20.71 3.42 ;
      RECT 20.38 0.02 20.55 0.19 ;
      RECT 20.38 2.74 20.55 2.91 ;
      RECT 20.38 5.46 20.55 5.63 ;
      RECT 19.92 0.02 20.09 0.19 ;
      RECT 19.92 2.74 20.09 2.91 ;
      RECT 19.92 5.46 20.09 5.63 ;
      RECT 19.865 1.21 20.035 1.38 ;
      RECT 17.935 -0.69 18.105 -0.52 ;
      RECT 17.935 0.79 18.105 0.96 ;
      RECT 17.935 4.71 18.105 4.88 ;
      RECT 17.935 6.19 18.105 6.36 ;
      RECT 17.585 -1.5 17.755 -1.33 ;
      RECT 17.585 2.56 17.755 2.73 ;
      RECT 17.585 2.94 17.755 3.11 ;
      RECT 17.585 7 17.755 7.17 ;
      RECT 17.565 1.16 17.735 1.33 ;
      RECT 17.565 4.34 17.735 4.51 ;
      RECT 16.945 -0.69 17.115 -0.52 ;
      RECT 16.945 0.79 17.115 0.96 ;
      RECT 16.945 4.71 17.115 4.88 ;
      RECT 16.945 6.19 17.115 6.36 ;
      RECT 16.595 -1.5 16.765 -1.33 ;
      RECT 16.595 2.56 16.765 2.73 ;
      RECT 16.595 2.94 16.765 3.11 ;
      RECT 16.595 7 16.765 7.17 ;
      RECT 16.575 1.16 16.745 1.33 ;
      RECT 16.575 4.34 16.745 4.51 ;
      RECT 15.89 -1.5 16.06 -1.33 ;
      RECT 15.89 2.56 16.06 2.73 ;
      RECT 15.89 2.94 16.06 3.11 ;
      RECT 15.89 7 16.06 7.17 ;
      RECT 15.58 0.42 15.75 0.59 ;
      RECT 15.58 5.08 15.75 5.25 ;
      RECT 15.21 -1.5 15.38 -1.33 ;
      RECT 15.21 7 15.38 7.17 ;
      RECT 15.15 -0.69 15.32 -0.52 ;
      RECT 15.15 0.05 15.32 0.22 ;
      RECT 15.15 5.45 15.32 5.62 ;
      RECT 15.15 6.19 15.32 6.36 ;
      RECT 14.775 0.79 14.945 0.96 ;
      RECT 14.775 4.71 14.945 4.88 ;
      RECT 14.53 -1.5 14.7 -1.33 ;
      RECT 14.53 7 14.7 7.17 ;
      RECT 13.85 -1.5 14.02 -1.33 ;
      RECT 13.85 7 14.02 7.17 ;
      RECT 13.78 1.16 13.95 1.33 ;
      RECT 13.78 4.34 13.95 4.51 ;
      RECT 12.19 0.02 12.36 0.19 ;
      RECT 12.19 2.74 12.36 2.91 ;
      RECT 12.19 5.46 12.36 5.63 ;
      RECT 12.15 1.21 12.32 1.38 ;
      RECT 11.81 3.25 11.98 3.42 ;
      RECT 11.73 0.02 11.9 0.19 ;
      RECT 11.73 1.55 11.9 1.72 ;
      RECT 11.73 2.74 11.9 2.91 ;
      RECT 11.73 5.46 11.9 5.63 ;
      RECT 11.27 0.02 11.44 0.19 ;
      RECT 11.27 2.74 11.44 2.91 ;
      RECT 11.27 5.46 11.44 5.63 ;
      RECT 11.13 4.27 11.3 4.44 ;
      RECT 10.81 0.02 10.98 0.19 ;
      RECT 10.81 2.74 10.98 2.91 ;
      RECT 10.81 5.46 10.98 5.63 ;
      RECT 10.79 0.53 10.96 0.7 ;
      RECT 10.45 4.27 10.62 4.44 ;
      RECT 10.35 0.02 10.52 0.19 ;
      RECT 10.35 2.74 10.52 2.91 ;
      RECT 10.35 5.46 10.52 5.63 ;
      RECT 9.995 0.53 10.165 0.7 ;
      RECT 9.89 0.02 10.06 0.19 ;
      RECT 9.89 2.74 10.06 2.91 ;
      RECT 9.89 5.46 10.06 5.63 ;
      RECT 9.77 2.23 9.94 2.4 ;
      RECT 9.77 4.27 9.94 4.44 ;
      RECT 9.43 0.02 9.6 0.19 ;
      RECT 9.43 2.74 9.6 2.91 ;
      RECT 9.43 5.46 9.6 5.63 ;
      RECT 9.26 4.27 9.43 4.44 ;
      RECT 9.09 0.87 9.26 1.04 ;
      RECT 8.97 0.02 9.14 0.19 ;
      RECT 8.97 2.74 9.14 2.91 ;
      RECT 8.97 5.46 9.14 5.63 ;
      RECT 8.51 0.02 8.68 0.19 ;
      RECT 8.51 2.74 8.68 2.91 ;
      RECT 8.51 5.46 8.68 5.63 ;
      RECT 8.07 4.27 8.24 4.44 ;
      RECT 8.05 0.02 8.22 0.19 ;
      RECT 8.05 2.74 8.22 2.91 ;
      RECT 8.05 5.46 8.22 5.63 ;
      RECT 7.73 0.87 7.9 1.04 ;
      RECT 7.59 0.02 7.76 0.19 ;
      RECT 7.59 2.74 7.76 2.91 ;
      RECT 7.59 5.46 7.76 5.63 ;
      RECT 7.56 2.23 7.73 2.4 ;
      RECT 7.13 0.02 7.3 0.19 ;
      RECT 7.13 2.74 7.3 2.91 ;
      RECT 7.13 5.46 7.3 5.63 ;
      RECT 7.05 4.27 7.22 4.44 ;
      RECT 6.67 0.02 6.84 0.19 ;
      RECT 6.67 2.74 6.84 2.91 ;
      RECT 6.67 5.46 6.84 5.63 ;
      RECT 6.37 3.25 6.54 3.42 ;
      RECT 6.21 0.02 6.38 0.19 ;
      RECT 6.21 2.74 6.38 2.91 ;
      RECT 6.21 5.46 6.38 5.63 ;
      RECT 5.75 0.02 5.92 0.19 ;
      RECT 5.75 2.74 5.92 2.91 ;
      RECT 5.75 5.46 5.92 5.63 ;
      RECT 5.695 1.21 5.865 1.38 ;
    LAYER li ;
      RECT 62.38 -1.605 62.64 1.01 ;
      RECT 48.205 -1.605 48.465 1.01 ;
      RECT 34.035 -1.605 34.295 1.01 ;
      RECT 19.86 -1.605 20.12 1.01 ;
      RECT 5.69 -1.605 5.95 1.01 ;
      RECT 68.83 -1.605 69.1 1 ;
      RECT 67.92 -1.605 68.16 1 ;
      RECT 54.655 -1.605 54.925 1 ;
      RECT 53.745 -1.605 53.985 1 ;
      RECT 40.485 -1.605 40.755 1 ;
      RECT 39.575 -1.605 39.815 1 ;
      RECT 26.31 -1.605 26.58 1 ;
      RECT 25.4 -1.605 25.64 1 ;
      RECT 12.14 -1.605 12.41 1 ;
      RECT 11.23 -1.605 11.47 1 ;
      RECT 67.05 -1.605 67.3 0.73 ;
      RECT 52.875 -1.605 53.125 0.73 ;
      RECT 38.705 -1.605 38.955 0.73 ;
      RECT 24.53 -1.605 24.78 0.73 ;
      RECT 10.36 -1.605 10.61 0.73 ;
      RECT 64.67 -1.605 65 0.65 ;
      RECT 50.495 -1.605 50.825 0.65 ;
      RECT 36.325 -1.605 36.655 0.65 ;
      RECT 22.15 -1.605 22.48 0.65 ;
      RECT 7.98 -1.605 8.31 0.65 ;
      RECT 62.295 -1.605 69.385 0.19 ;
      RECT 48.12 -1.605 55.21 0.19 ;
      RECT 33.95 -1.605 41.04 0.19 ;
      RECT 19.775 -1.605 26.865 0.19 ;
      RECT 5.605 -1.605 12.695 0.19 ;
      RECT 62.04 -1.605 69.385 0.05 ;
      RECT 47.865 -1.605 55.21 0.05 ;
      RECT 33.695 -1.605 41.04 0.05 ;
      RECT 19.52 -1.605 26.865 0.05 ;
      RECT 5.35 -1.605 12.695 0.05 ;
      RECT 74.195 -1.605 74.365 -0.67 ;
      RECT 73.205 -1.605 73.375 -0.67 ;
      RECT 70.46 -1.605 70.63 -0.67 ;
      RECT 60.02 -1.605 60.19 -0.67 ;
      RECT 59.03 -1.605 59.2 -0.67 ;
      RECT 56.285 -1.605 56.455 -0.67 ;
      RECT 45.85 -1.605 46.02 -0.67 ;
      RECT 44.86 -1.605 45.03 -0.67 ;
      RECT 42.115 -1.605 42.285 -0.67 ;
      RECT 31.675 -1.605 31.845 -0.67 ;
      RECT 30.685 -1.605 30.855 -0.67 ;
      RECT 27.94 -1.605 28.11 -0.67 ;
      RECT 17.505 -1.605 17.675 -0.67 ;
      RECT 16.515 -1.605 16.685 -0.67 ;
      RECT 13.77 -1.605 13.94 -0.67 ;
      RECT 4.005 -1.605 75.165 -1.3 ;
      RECT 74.195 1.8 74.365 3.87 ;
      RECT 73.205 1.8 73.375 3.87 ;
      RECT 70.46 1.8 70.63 3.87 ;
      RECT 60.02 1.8 60.19 3.87 ;
      RECT 59.03 1.8 59.2 3.87 ;
      RECT 56.285 1.8 56.455 3.87 ;
      RECT 45.85 1.8 46.02 3.87 ;
      RECT 44.86 1.8 45.03 3.87 ;
      RECT 42.115 1.8 42.285 3.87 ;
      RECT 31.675 1.8 31.845 3.87 ;
      RECT 30.685 1.8 30.855 3.87 ;
      RECT 27.94 1.8 28.11 3.87 ;
      RECT 17.505 1.8 17.675 3.87 ;
      RECT 16.515 1.8 16.685 3.87 ;
      RECT 13.77 1.8 13.94 3.87 ;
      RECT 65.65 2.085 65.915 3.69 ;
      RECT 51.475 2.085 51.74 3.69 ;
      RECT 37.305 2.085 37.57 3.69 ;
      RECT 23.13 2.085 23.395 3.69 ;
      RECT 8.96 2.085 9.225 3.69 ;
      RECT 63.49 2.235 63.82 3.63 ;
      RECT 49.315 2.235 49.645 3.63 ;
      RECT 35.145 2.235 35.475 3.63 ;
      RECT 20.97 2.235 21.3 3.63 ;
      RECT 6.8 2.235 7.13 3.63 ;
      RECT 64.49 2.74 64.77 3.58 ;
      RECT 50.315 2.74 50.595 3.58 ;
      RECT 36.145 2.74 36.425 3.58 ;
      RECT 21.97 2.74 22.25 3.58 ;
      RECT 7.8 2.74 8.08 3.58 ;
      RECT 66.465 2.74 66.84 3.29 ;
      RECT 52.29 2.74 52.665 3.29 ;
      RECT 38.12 2.74 38.495 3.29 ;
      RECT 23.945 2.74 24.32 3.29 ;
      RECT 9.775 2.74 10.15 3.29 ;
      RECT 69.225 2.53 75.165 3.14 ;
      RECT 55.05 2.53 60.99 3.14 ;
      RECT 40.88 2.53 46.82 3.14 ;
      RECT 26.705 2.53 32.645 3.14 ;
      RECT 12.535 2.53 18.475 3.14 ;
      RECT 60.695 2.525 62.155 3.135 ;
      RECT 46.52 2.525 47.98 3.135 ;
      RECT 32.35 2.525 33.81 3.135 ;
      RECT 18.175 2.525 19.635 3.135 ;
      RECT 4.005 2.525 5.465 3.135 ;
      RECT 69.095 2.53 75.165 3.065 ;
      RECT 54.92 2.53 62.155 3.065 ;
      RECT 40.75 2.53 47.98 3.065 ;
      RECT 26.575 2.53 33.81 3.065 ;
      RECT 12.405 2.53 19.635 3.065 ;
      RECT 4.005 2.74 75.165 2.91 ;
      RECT 68.77 1.6 69.1 2.91 ;
      RECT 67.03 2.195 67.285 2.91 ;
      RECT 65.6 2.085 66.205 2.91 ;
      RECT 64.73 2.195 64.945 2.91 ;
      RECT 63.3 2.235 63.915 2.91 ;
      RECT 63.72 1.87 63.915 2.91 ;
      RECT 62.38 2.23 62.64 2.91 ;
      RECT 54.595 1.6 54.925 2.91 ;
      RECT 52.855 2.195 53.11 2.91 ;
      RECT 51.425 2.085 52.03 2.91 ;
      RECT 50.555 2.195 50.77 2.91 ;
      RECT 49.125 2.235 49.74 2.91 ;
      RECT 49.545 1.87 49.74 2.91 ;
      RECT 48.205 2.23 48.465 2.91 ;
      RECT 40.425 1.6 40.755 2.91 ;
      RECT 38.685 2.195 38.94 2.91 ;
      RECT 37.255 2.085 37.86 2.91 ;
      RECT 36.385 2.195 36.6 2.91 ;
      RECT 34.955 2.235 35.57 2.91 ;
      RECT 35.375 1.87 35.57 2.91 ;
      RECT 34.035 2.23 34.295 2.91 ;
      RECT 26.25 1.6 26.58 2.91 ;
      RECT 24.51 2.195 24.765 2.91 ;
      RECT 23.08 2.085 23.685 2.91 ;
      RECT 22.21 2.195 22.425 2.91 ;
      RECT 20.78 2.235 21.395 2.91 ;
      RECT 21.2 1.87 21.395 2.91 ;
      RECT 19.86 2.23 20.12 2.91 ;
      RECT 12.08 1.6 12.41 2.91 ;
      RECT 10.34 2.195 10.595 2.91 ;
      RECT 8.91 2.085 9.515 2.91 ;
      RECT 8.04 2.195 8.255 2.91 ;
      RECT 6.61 2.235 7.225 2.91 ;
      RECT 7.03 1.87 7.225 2.91 ;
      RECT 5.69 2.23 5.95 2.91 ;
      RECT 66.03 1.815 66.215 2.185 ;
      RECT 51.855 1.815 52.04 2.185 ;
      RECT 37.685 1.815 37.87 2.185 ;
      RECT 23.51 1.815 23.695 2.185 ;
      RECT 9.34 1.815 9.525 2.185 ;
      RECT 66.03 1.815 66.36 2.06 ;
      RECT 63.72 1.87 64.05 2.06 ;
      RECT 51.855 1.815 52.185 2.06 ;
      RECT 49.545 1.87 49.875 2.06 ;
      RECT 37.685 1.815 38.015 2.06 ;
      RECT 35.375 1.87 35.705 2.06 ;
      RECT 23.51 1.815 23.84 2.06 ;
      RECT 21.2 1.87 21.53 2.06 ;
      RECT 9.34 1.815 9.67 2.06 ;
      RECT 7.03 1.87 7.36 2.06 ;
      RECT 4.005 6.97 75.165 7.275 ;
      RECT 74.195 6.34 74.365 7.275 ;
      RECT 73.205 6.34 73.375 7.275 ;
      RECT 70.46 6.34 70.63 7.275 ;
      RECT 62 5.575 69.2 7.275 ;
      RECT 60.02 6.34 60.19 7.275 ;
      RECT 59.03 6.34 59.2 7.275 ;
      RECT 56.285 6.34 56.455 7.275 ;
      RECT 47.825 5.575 55.025 7.275 ;
      RECT 45.85 6.34 46.02 7.275 ;
      RECT 44.86 6.34 45.03 7.275 ;
      RECT 42.115 6.34 42.285 7.275 ;
      RECT 33.655 5.575 40.855 7.275 ;
      RECT 31.675 6.34 31.845 7.275 ;
      RECT 30.685 6.34 30.855 7.275 ;
      RECT 27.94 6.34 28.11 7.275 ;
      RECT 19.48 5.575 26.68 7.275 ;
      RECT 17.505 6.34 17.675 7.275 ;
      RECT 16.515 6.34 16.685 7.275 ;
      RECT 13.77 6.34 13.94 7.275 ;
      RECT 5.31 5.575 12.51 7.275 ;
      RECT 62.295 5.46 69.195 7.275 ;
      RECT 48.12 5.46 55.02 7.275 ;
      RECT 33.95 5.46 40.85 7.275 ;
      RECT 19.775 5.46 26.675 7.275 ;
      RECT 5.605 5.46 12.505 7.275 ;
      RECT 67.73 4.95 68.18 7.275 ;
      RECT 65.64 5.06 65.97 7.275 ;
      RECT 63.57 5 63.82 7.275 ;
      RECT 53.555 4.95 54.005 7.275 ;
      RECT 51.465 5.06 51.795 7.275 ;
      RECT 49.395 5 49.645 7.275 ;
      RECT 39.385 4.95 39.835 7.275 ;
      RECT 37.295 5.06 37.625 7.275 ;
      RECT 35.225 5 35.475 7.275 ;
      RECT 25.21 4.95 25.66 7.275 ;
      RECT 23.12 5.06 23.45 7.275 ;
      RECT 21.05 5 21.3 7.275 ;
      RECT 11.04 4.95 11.49 7.275 ;
      RECT 8.95 5.06 9.28 7.275 ;
      RECT 6.88 5 7.13 7.275 ;
      RECT 74.255 0.135 74.425 1.33 ;
      RECT 74.255 0.135 74.72 0.305 ;
      RECT 74.255 5.365 74.72 5.535 ;
      RECT 74.255 4.34 74.425 5.535 ;
      RECT 73.265 0.135 73.435 1.33 ;
      RECT 73.265 0.135 73.73 0.305 ;
      RECT 73.265 5.365 73.73 5.535 ;
      RECT 73.265 4.34 73.435 5.535 ;
      RECT 71.41 1.03 71.58 2.26 ;
      RECT 71.465 -0.75 71.635 1.2 ;
      RECT 71.41 -1.03 71.58 -0.58 ;
      RECT 71.41 6.25 71.58 6.7 ;
      RECT 71.465 4.47 71.635 6.42 ;
      RECT 71.41 3.41 71.58 4.64 ;
      RECT 70.89 -1.03 71.06 2.26 ;
      RECT 70.89 0.47 71.295 0.8 ;
      RECT 70.89 -0.37 71.295 -0.04 ;
      RECT 70.89 3.41 71.06 6.7 ;
      RECT 70.89 5.71 71.295 6.04 ;
      RECT 70.89 4.87 71.295 5.2 ;
      RECT 66.15 5.04 67.455 5.29 ;
      RECT 66.15 4.72 66.33 5.29 ;
      RECT 65.6 4.72 66.33 4.89 ;
      RECT 65.6 3.88 65.77 4.89 ;
      RECT 66.435 3.92 68.18 4.1 ;
      RECT 67.85 3.08 68.18 4.1 ;
      RECT 65.6 3.88 66.66 4.05 ;
      RECT 67.85 3.25 68.67 3.42 ;
      RECT 67.01 3.08 67.34 3.29 ;
      RECT 67.01 3.08 68.18 3.25 ;
      RECT 67.91 1.6 68.24 2.555 ;
      RECT 67.91 1.6 68.59 1.77 ;
      RECT 68.42 0.36 68.59 1.77 ;
      RECT 68.33 0.36 68.66 1 ;
      RECT 67.455 1.87 67.73 2.57 ;
      RECT 67.56 0.36 67.73 2.57 ;
      RECT 67.9 1.18 68.25 1.43 ;
      RECT 67.56 1.21 68.25 1.38 ;
      RECT 67.47 0.36 67.73 0.84 ;
      RECT 66.8 3.51 67.68 3.75 ;
      RECT 67.45 3.42 67.68 3.75 ;
      RECT 66.15 3.51 67.68 3.71 ;
      RECT 67.065 3.46 67.68 3.75 ;
      RECT 66.15 3.38 66.32 3.71 ;
      RECT 67.035 4.27 67.285 4.87 ;
      RECT 67.035 4.27 67.51 4.47 ;
      RECT 66.53 1.49 67.285 1.99 ;
      RECT 65.6 1.295 65.86 1.915 ;
      RECT 66.515 1.435 66.53 1.74 ;
      RECT 66.5 1.42 66.52 1.705 ;
      RECT 67.16 1.095 67.39 1.695 ;
      RECT 66.475 1.365 66.495 1.68 ;
      RECT 66.455 1.49 67.39 1.665 ;
      RECT 66.43 1.49 67.39 1.655 ;
      RECT 66.36 1.49 67.39 1.645 ;
      RECT 66.34 1.49 67.39 1.615 ;
      RECT 66.32 0.4 66.49 1.585 ;
      RECT 66.29 1.49 67.39 1.555 ;
      RECT 66.255 1.49 67.39 1.53 ;
      RECT 66.225 1.485 66.615 1.495 ;
      RECT 66.225 1.475 66.59 1.495 ;
      RECT 66.225 1.47 66.575 1.495 ;
      RECT 66.225 1.46 66.56 1.495 ;
      RECT 65.6 1.295 66.49 1.465 ;
      RECT 65.6 1.45 66.55 1.465 ;
      RECT 65.6 1.445 66.54 1.465 ;
      RECT 66.495 1.39 66.505 1.695 ;
      RECT 65.6 1.425 66.525 1.465 ;
      RECT 65.6 1.405 66.51 1.465 ;
      RECT 65.6 0.4 66.49 0.57 ;
      RECT 66.66 0.895 66.99 1.32 ;
      RECT 66.66 0.41 66.88 1.32 ;
      RECT 66.575 4.27 66.785 4.87 ;
      RECT 66.435 4.27 66.785 4.47 ;
      RECT 65.155 1.87 65.43 2.57 ;
      RECT 65.375 0.36 65.43 2.57 ;
      RECT 65.26 1.165 65.43 2.57 ;
      RECT 65.26 0.36 65.43 1.16 ;
      RECT 65.17 0.36 65.43 0.835 ;
      RECT 63.3 1.53 63.55 2.065 ;
      RECT 64.27 1.53 64.985 1.995 ;
      RECT 63.3 1.53 65.09 1.7 ;
      RECT 64.86 1.165 65.09 1.7 ;
      RECT 63.855 0.41 64.11 1.7 ;
      RECT 64.86 1.1 64.92 1.995 ;
      RECT 64.92 1.095 65.09 1.16 ;
      RECT 63.32 0.41 64.11 0.675 ;
      RECT 64.28 4.22 64.955 4.47 ;
      RECT 64.69 3.86 64.955 4.47 ;
      RECT 64.44 4.64 64.77 5.19 ;
      RECT 63.38 4.64 64.77 4.83 ;
      RECT 63.38 3.8 63.55 4.83 ;
      RECT 63.26 4.22 63.55 4.55 ;
      RECT 63.38 3.8 64.32 3.97 ;
      RECT 64.02 3.25 64.32 3.97 ;
      RECT 64.28 0.83 64.69 1.35 ;
      RECT 64.28 0.41 64.48 1.35 ;
      RECT 62.89 0.59 63.06 2.57 ;
      RECT 62.89 1.1 63.685 1.35 ;
      RECT 62.89 0.59 63.14 1.35 ;
      RECT 62.81 0.59 63.14 1.01 ;
      RECT 62.84 5 63.4 5.29 ;
      RECT 62.84 3.08 63.09 5.29 ;
      RECT 62.84 3.08 63.3 3.63 ;
      RECT 60.08 0.135 60.25 1.33 ;
      RECT 60.08 0.135 60.545 0.305 ;
      RECT 60.08 5.365 60.545 5.535 ;
      RECT 60.08 4.34 60.25 5.535 ;
      RECT 59.09 0.135 59.26 1.33 ;
      RECT 59.09 0.135 59.555 0.305 ;
      RECT 59.09 5.365 59.555 5.535 ;
      RECT 59.09 4.34 59.26 5.535 ;
      RECT 57.235 1.03 57.405 2.26 ;
      RECT 57.29 -0.75 57.46 1.2 ;
      RECT 57.235 -1.03 57.405 -0.58 ;
      RECT 57.235 6.25 57.405 6.7 ;
      RECT 57.29 4.47 57.46 6.42 ;
      RECT 57.235 3.41 57.405 4.64 ;
      RECT 56.715 -1.03 56.885 2.26 ;
      RECT 56.715 0.47 57.12 0.8 ;
      RECT 56.715 -0.37 57.12 -0.04 ;
      RECT 56.715 3.41 56.885 6.7 ;
      RECT 56.715 5.71 57.12 6.04 ;
      RECT 56.715 4.87 57.12 5.2 ;
      RECT 51.975 5.04 53.28 5.29 ;
      RECT 51.975 4.72 52.155 5.29 ;
      RECT 51.425 4.72 52.155 4.89 ;
      RECT 51.425 3.88 51.595 4.89 ;
      RECT 52.26 3.92 54.005 4.1 ;
      RECT 53.675 3.08 54.005 4.1 ;
      RECT 51.425 3.88 52.485 4.05 ;
      RECT 53.675 3.25 54.495 3.42 ;
      RECT 52.835 3.08 53.165 3.29 ;
      RECT 52.835 3.08 54.005 3.25 ;
      RECT 53.735 1.6 54.065 2.555 ;
      RECT 53.735 1.6 54.415 1.77 ;
      RECT 54.245 0.36 54.415 1.77 ;
      RECT 54.155 0.36 54.485 1 ;
      RECT 53.28 1.87 53.555 2.57 ;
      RECT 53.385 0.36 53.555 2.57 ;
      RECT 53.725 1.18 54.075 1.43 ;
      RECT 53.385 1.21 54.075 1.38 ;
      RECT 53.295 0.36 53.555 0.84 ;
      RECT 52.625 3.51 53.505 3.75 ;
      RECT 53.275 3.42 53.505 3.75 ;
      RECT 51.975 3.51 53.505 3.71 ;
      RECT 52.89 3.46 53.505 3.75 ;
      RECT 51.975 3.38 52.145 3.71 ;
      RECT 52.86 4.27 53.11 4.87 ;
      RECT 52.86 4.27 53.335 4.47 ;
      RECT 52.355 1.49 53.11 1.99 ;
      RECT 51.425 1.295 51.685 1.915 ;
      RECT 52.34 1.435 52.355 1.74 ;
      RECT 52.325 1.42 52.345 1.705 ;
      RECT 52.985 1.095 53.215 1.695 ;
      RECT 52.3 1.365 52.32 1.68 ;
      RECT 52.28 1.49 53.215 1.665 ;
      RECT 52.255 1.49 53.215 1.655 ;
      RECT 52.185 1.49 53.215 1.645 ;
      RECT 52.165 1.49 53.215 1.615 ;
      RECT 52.145 0.4 52.315 1.585 ;
      RECT 52.115 1.49 53.215 1.555 ;
      RECT 52.08 1.49 53.215 1.53 ;
      RECT 52.05 1.485 52.44 1.495 ;
      RECT 52.05 1.475 52.415 1.495 ;
      RECT 52.05 1.47 52.4 1.495 ;
      RECT 52.05 1.46 52.385 1.495 ;
      RECT 51.425 1.295 52.315 1.465 ;
      RECT 51.425 1.45 52.375 1.465 ;
      RECT 51.425 1.445 52.365 1.465 ;
      RECT 52.32 1.39 52.33 1.695 ;
      RECT 51.425 1.425 52.35 1.465 ;
      RECT 51.425 1.405 52.335 1.465 ;
      RECT 51.425 0.4 52.315 0.57 ;
      RECT 52.485 0.895 52.815 1.32 ;
      RECT 52.485 0.41 52.705 1.32 ;
      RECT 52.4 4.27 52.61 4.87 ;
      RECT 52.26 4.27 52.61 4.47 ;
      RECT 50.98 1.87 51.255 2.57 ;
      RECT 51.2 0.36 51.255 2.57 ;
      RECT 51.085 1.165 51.255 2.57 ;
      RECT 51.085 0.36 51.255 1.16 ;
      RECT 50.995 0.36 51.255 0.835 ;
      RECT 49.125 1.53 49.375 2.065 ;
      RECT 50.095 1.53 50.81 1.995 ;
      RECT 49.125 1.53 50.915 1.7 ;
      RECT 50.685 1.165 50.915 1.7 ;
      RECT 49.68 0.41 49.935 1.7 ;
      RECT 50.685 1.1 50.745 1.995 ;
      RECT 50.745 1.095 50.915 1.16 ;
      RECT 49.145 0.41 49.935 0.675 ;
      RECT 50.105 4.22 50.78 4.47 ;
      RECT 50.515 3.86 50.78 4.47 ;
      RECT 50.265 4.64 50.595 5.19 ;
      RECT 49.205 4.64 50.595 4.83 ;
      RECT 49.205 3.8 49.375 4.83 ;
      RECT 49.085 4.22 49.375 4.55 ;
      RECT 49.205 3.8 50.145 3.97 ;
      RECT 49.845 3.25 50.145 3.97 ;
      RECT 50.105 0.83 50.515 1.35 ;
      RECT 50.105 0.41 50.305 1.35 ;
      RECT 48.715 0.59 48.885 2.57 ;
      RECT 48.715 1.1 49.51 1.35 ;
      RECT 48.715 0.59 48.965 1.35 ;
      RECT 48.635 0.59 48.965 1.01 ;
      RECT 48.665 5 49.225 5.29 ;
      RECT 48.665 3.08 48.915 5.29 ;
      RECT 48.665 3.08 49.125 3.63 ;
      RECT 45.91 0.135 46.08 1.33 ;
      RECT 45.91 0.135 46.375 0.305 ;
      RECT 45.91 5.365 46.375 5.535 ;
      RECT 45.91 4.34 46.08 5.535 ;
      RECT 44.92 0.135 45.09 1.33 ;
      RECT 44.92 0.135 45.385 0.305 ;
      RECT 44.92 5.365 45.385 5.535 ;
      RECT 44.92 4.34 45.09 5.535 ;
      RECT 43.065 1.03 43.235 2.26 ;
      RECT 43.12 -0.75 43.29 1.2 ;
      RECT 43.065 -1.03 43.235 -0.58 ;
      RECT 43.065 6.25 43.235 6.7 ;
      RECT 43.12 4.47 43.29 6.42 ;
      RECT 43.065 3.41 43.235 4.64 ;
      RECT 42.545 -1.03 42.715 2.26 ;
      RECT 42.545 0.47 42.95 0.8 ;
      RECT 42.545 -0.37 42.95 -0.04 ;
      RECT 42.545 3.41 42.715 6.7 ;
      RECT 42.545 5.71 42.95 6.04 ;
      RECT 42.545 4.87 42.95 5.2 ;
      RECT 37.805 5.04 39.11 5.29 ;
      RECT 37.805 4.72 37.985 5.29 ;
      RECT 37.255 4.72 37.985 4.89 ;
      RECT 37.255 3.88 37.425 4.89 ;
      RECT 38.09 3.92 39.835 4.1 ;
      RECT 39.505 3.08 39.835 4.1 ;
      RECT 37.255 3.88 38.315 4.05 ;
      RECT 39.505 3.25 40.325 3.42 ;
      RECT 38.665 3.08 38.995 3.29 ;
      RECT 38.665 3.08 39.835 3.25 ;
      RECT 39.565 1.6 39.895 2.555 ;
      RECT 39.565 1.6 40.245 1.77 ;
      RECT 40.075 0.36 40.245 1.77 ;
      RECT 39.985 0.36 40.315 1 ;
      RECT 39.11 1.87 39.385 2.57 ;
      RECT 39.215 0.36 39.385 2.57 ;
      RECT 39.555 1.18 39.905 1.43 ;
      RECT 39.215 1.21 39.905 1.38 ;
      RECT 39.125 0.36 39.385 0.84 ;
      RECT 38.455 3.51 39.335 3.75 ;
      RECT 39.105 3.42 39.335 3.75 ;
      RECT 37.805 3.51 39.335 3.71 ;
      RECT 38.72 3.46 39.335 3.75 ;
      RECT 37.805 3.38 37.975 3.71 ;
      RECT 38.69 4.27 38.94 4.87 ;
      RECT 38.69 4.27 39.165 4.47 ;
      RECT 38.185 1.49 38.94 1.99 ;
      RECT 37.255 1.295 37.515 1.915 ;
      RECT 38.17 1.435 38.185 1.74 ;
      RECT 38.155 1.42 38.175 1.705 ;
      RECT 38.815 1.095 39.045 1.695 ;
      RECT 38.13 1.365 38.15 1.68 ;
      RECT 38.11 1.49 39.045 1.665 ;
      RECT 38.085 1.49 39.045 1.655 ;
      RECT 38.015 1.49 39.045 1.645 ;
      RECT 37.995 1.49 39.045 1.615 ;
      RECT 37.975 0.4 38.145 1.585 ;
      RECT 37.945 1.49 39.045 1.555 ;
      RECT 37.91 1.49 39.045 1.53 ;
      RECT 37.88 1.485 38.27 1.495 ;
      RECT 37.88 1.475 38.245 1.495 ;
      RECT 37.88 1.47 38.23 1.495 ;
      RECT 37.88 1.46 38.215 1.495 ;
      RECT 37.255 1.295 38.145 1.465 ;
      RECT 37.255 1.45 38.205 1.465 ;
      RECT 37.255 1.445 38.195 1.465 ;
      RECT 38.15 1.39 38.16 1.695 ;
      RECT 37.255 1.425 38.18 1.465 ;
      RECT 37.255 1.405 38.165 1.465 ;
      RECT 37.255 0.4 38.145 0.57 ;
      RECT 38.315 0.895 38.645 1.32 ;
      RECT 38.315 0.41 38.535 1.32 ;
      RECT 38.23 4.27 38.44 4.87 ;
      RECT 38.09 4.27 38.44 4.47 ;
      RECT 36.81 1.87 37.085 2.57 ;
      RECT 37.03 0.36 37.085 2.57 ;
      RECT 36.915 1.165 37.085 2.57 ;
      RECT 36.915 0.36 37.085 1.16 ;
      RECT 36.825 0.36 37.085 0.835 ;
      RECT 34.955 1.53 35.205 2.065 ;
      RECT 35.925 1.53 36.64 1.995 ;
      RECT 34.955 1.53 36.745 1.7 ;
      RECT 36.515 1.165 36.745 1.7 ;
      RECT 35.51 0.41 35.765 1.7 ;
      RECT 36.515 1.1 36.575 1.995 ;
      RECT 36.575 1.095 36.745 1.16 ;
      RECT 34.975 0.41 35.765 0.675 ;
      RECT 35.935 4.22 36.61 4.47 ;
      RECT 36.345 3.86 36.61 4.47 ;
      RECT 36.095 4.64 36.425 5.19 ;
      RECT 35.035 4.64 36.425 4.83 ;
      RECT 35.035 3.8 35.205 4.83 ;
      RECT 34.915 4.22 35.205 4.55 ;
      RECT 35.035 3.8 35.975 3.97 ;
      RECT 35.675 3.25 35.975 3.97 ;
      RECT 35.935 0.83 36.345 1.35 ;
      RECT 35.935 0.41 36.135 1.35 ;
      RECT 34.545 0.59 34.715 2.57 ;
      RECT 34.545 1.1 35.34 1.35 ;
      RECT 34.545 0.59 34.795 1.35 ;
      RECT 34.465 0.59 34.795 1.01 ;
      RECT 34.495 5 35.055 5.29 ;
      RECT 34.495 3.08 34.745 5.29 ;
      RECT 34.495 3.08 34.955 3.63 ;
      RECT 31.735 0.135 31.905 1.33 ;
      RECT 31.735 0.135 32.2 0.305 ;
      RECT 31.735 5.365 32.2 5.535 ;
      RECT 31.735 4.34 31.905 5.535 ;
      RECT 30.745 0.135 30.915 1.33 ;
      RECT 30.745 0.135 31.21 0.305 ;
      RECT 30.745 5.365 31.21 5.535 ;
      RECT 30.745 4.34 30.915 5.535 ;
      RECT 28.89 1.03 29.06 2.26 ;
      RECT 28.945 -0.75 29.115 1.2 ;
      RECT 28.89 -1.03 29.06 -0.58 ;
      RECT 28.89 6.25 29.06 6.7 ;
      RECT 28.945 4.47 29.115 6.42 ;
      RECT 28.89 3.41 29.06 4.64 ;
      RECT 28.37 -1.03 28.54 2.26 ;
      RECT 28.37 0.47 28.775 0.8 ;
      RECT 28.37 -0.37 28.775 -0.04 ;
      RECT 28.37 3.41 28.54 6.7 ;
      RECT 28.37 5.71 28.775 6.04 ;
      RECT 28.37 4.87 28.775 5.2 ;
      RECT 23.63 5.04 24.935 5.29 ;
      RECT 23.63 4.72 23.81 5.29 ;
      RECT 23.08 4.72 23.81 4.89 ;
      RECT 23.08 3.88 23.25 4.89 ;
      RECT 23.915 3.92 25.66 4.1 ;
      RECT 25.33 3.08 25.66 4.1 ;
      RECT 23.08 3.88 24.14 4.05 ;
      RECT 25.33 3.25 26.15 3.42 ;
      RECT 24.49 3.08 24.82 3.29 ;
      RECT 24.49 3.08 25.66 3.25 ;
      RECT 25.39 1.6 25.72 2.555 ;
      RECT 25.39 1.6 26.07 1.77 ;
      RECT 25.9 0.36 26.07 1.77 ;
      RECT 25.81 0.36 26.14 1 ;
      RECT 24.935 1.87 25.21 2.57 ;
      RECT 25.04 0.36 25.21 2.57 ;
      RECT 25.38 1.18 25.73 1.43 ;
      RECT 25.04 1.21 25.73 1.38 ;
      RECT 24.95 0.36 25.21 0.84 ;
      RECT 24.28 3.51 25.16 3.75 ;
      RECT 24.93 3.42 25.16 3.75 ;
      RECT 23.63 3.51 25.16 3.71 ;
      RECT 24.545 3.46 25.16 3.75 ;
      RECT 23.63 3.38 23.8 3.71 ;
      RECT 24.515 4.27 24.765 4.87 ;
      RECT 24.515 4.27 24.99 4.47 ;
      RECT 24.01 1.49 24.765 1.99 ;
      RECT 23.08 1.295 23.34 1.915 ;
      RECT 23.995 1.435 24.01 1.74 ;
      RECT 23.98 1.42 24 1.705 ;
      RECT 24.64 1.095 24.87 1.695 ;
      RECT 23.955 1.365 23.975 1.68 ;
      RECT 23.935 1.49 24.87 1.665 ;
      RECT 23.91 1.49 24.87 1.655 ;
      RECT 23.84 1.49 24.87 1.645 ;
      RECT 23.82 1.49 24.87 1.615 ;
      RECT 23.8 0.4 23.97 1.585 ;
      RECT 23.77 1.49 24.87 1.555 ;
      RECT 23.735 1.49 24.87 1.53 ;
      RECT 23.705 1.485 24.095 1.495 ;
      RECT 23.705 1.475 24.07 1.495 ;
      RECT 23.705 1.47 24.055 1.495 ;
      RECT 23.705 1.46 24.04 1.495 ;
      RECT 23.08 1.295 23.97 1.465 ;
      RECT 23.08 1.45 24.03 1.465 ;
      RECT 23.08 1.445 24.02 1.465 ;
      RECT 23.975 1.39 23.985 1.695 ;
      RECT 23.08 1.425 24.005 1.465 ;
      RECT 23.08 1.405 23.99 1.465 ;
      RECT 23.08 0.4 23.97 0.57 ;
      RECT 24.14 0.895 24.47 1.32 ;
      RECT 24.14 0.41 24.36 1.32 ;
      RECT 24.055 4.27 24.265 4.87 ;
      RECT 23.915 4.27 24.265 4.47 ;
      RECT 22.635 1.87 22.91 2.57 ;
      RECT 22.855 0.36 22.91 2.57 ;
      RECT 22.74 1.165 22.91 2.57 ;
      RECT 22.74 0.36 22.91 1.16 ;
      RECT 22.65 0.36 22.91 0.835 ;
      RECT 20.78 1.53 21.03 2.065 ;
      RECT 21.75 1.53 22.465 1.995 ;
      RECT 20.78 1.53 22.57 1.7 ;
      RECT 22.34 1.165 22.57 1.7 ;
      RECT 21.335 0.41 21.59 1.7 ;
      RECT 22.34 1.1 22.4 1.995 ;
      RECT 22.4 1.095 22.57 1.16 ;
      RECT 20.8 0.41 21.59 0.675 ;
      RECT 21.76 4.22 22.435 4.47 ;
      RECT 22.17 3.86 22.435 4.47 ;
      RECT 21.92 4.64 22.25 5.19 ;
      RECT 20.86 4.64 22.25 4.83 ;
      RECT 20.86 3.8 21.03 4.83 ;
      RECT 20.74 4.22 21.03 4.55 ;
      RECT 20.86 3.8 21.8 3.97 ;
      RECT 21.5 3.25 21.8 3.97 ;
      RECT 21.76 0.83 22.17 1.35 ;
      RECT 21.76 0.41 21.96 1.35 ;
      RECT 20.37 0.59 20.54 2.57 ;
      RECT 20.37 1.1 21.165 1.35 ;
      RECT 20.37 0.59 20.62 1.35 ;
      RECT 20.29 0.59 20.62 1.01 ;
      RECT 20.32 5 20.88 5.29 ;
      RECT 20.32 3.08 20.57 5.29 ;
      RECT 20.32 3.08 20.78 3.63 ;
      RECT 17.565 0.135 17.735 1.33 ;
      RECT 17.565 0.135 18.03 0.305 ;
      RECT 17.565 5.365 18.03 5.535 ;
      RECT 17.565 4.34 17.735 5.535 ;
      RECT 16.575 0.135 16.745 1.33 ;
      RECT 16.575 0.135 17.04 0.305 ;
      RECT 16.575 5.365 17.04 5.535 ;
      RECT 16.575 4.34 16.745 5.535 ;
      RECT 14.72 1.03 14.89 2.26 ;
      RECT 14.775 -0.75 14.945 1.2 ;
      RECT 14.72 -1.03 14.89 -0.58 ;
      RECT 14.72 6.25 14.89 6.7 ;
      RECT 14.775 4.47 14.945 6.42 ;
      RECT 14.72 3.41 14.89 4.64 ;
      RECT 14.2 -1.03 14.37 2.26 ;
      RECT 14.2 0.47 14.605 0.8 ;
      RECT 14.2 -0.37 14.605 -0.04 ;
      RECT 14.2 3.41 14.37 6.7 ;
      RECT 14.2 5.71 14.605 6.04 ;
      RECT 14.2 4.87 14.605 5.2 ;
      RECT 9.46 5.04 10.765 5.29 ;
      RECT 9.46 4.72 9.64 5.29 ;
      RECT 8.91 4.72 9.64 4.89 ;
      RECT 8.91 3.88 9.08 4.89 ;
      RECT 9.745 3.92 11.49 4.1 ;
      RECT 11.16 3.08 11.49 4.1 ;
      RECT 8.91 3.88 9.97 4.05 ;
      RECT 11.16 3.25 11.98 3.42 ;
      RECT 10.32 3.08 10.65 3.29 ;
      RECT 10.32 3.08 11.49 3.25 ;
      RECT 11.22 1.6 11.55 2.555 ;
      RECT 11.22 1.6 11.9 1.77 ;
      RECT 11.73 0.36 11.9 1.77 ;
      RECT 11.64 0.36 11.97 1 ;
      RECT 10.765 1.87 11.04 2.57 ;
      RECT 10.87 0.36 11.04 2.57 ;
      RECT 11.21 1.18 11.56 1.43 ;
      RECT 10.87 1.21 11.56 1.38 ;
      RECT 10.78 0.36 11.04 0.84 ;
      RECT 10.11 3.51 10.99 3.75 ;
      RECT 10.76 3.42 10.99 3.75 ;
      RECT 9.46 3.51 10.99 3.71 ;
      RECT 10.375 3.46 10.99 3.75 ;
      RECT 9.46 3.38 9.63 3.71 ;
      RECT 10.345 4.27 10.595 4.87 ;
      RECT 10.345 4.27 10.82 4.47 ;
      RECT 9.84 1.49 10.595 1.99 ;
      RECT 8.91 1.295 9.17 1.915 ;
      RECT 9.825 1.435 9.84 1.74 ;
      RECT 9.81 1.42 9.83 1.705 ;
      RECT 10.47 1.095 10.7 1.695 ;
      RECT 9.785 1.365 9.805 1.68 ;
      RECT 9.765 1.49 10.7 1.665 ;
      RECT 9.74 1.49 10.7 1.655 ;
      RECT 9.67 1.49 10.7 1.645 ;
      RECT 9.65 1.49 10.7 1.615 ;
      RECT 9.63 0.4 9.8 1.585 ;
      RECT 9.6 1.49 10.7 1.555 ;
      RECT 9.565 1.49 10.7 1.53 ;
      RECT 9.535 1.485 9.925 1.495 ;
      RECT 9.535 1.475 9.9 1.495 ;
      RECT 9.535 1.47 9.885 1.495 ;
      RECT 9.535 1.46 9.87 1.495 ;
      RECT 8.91 1.295 9.8 1.465 ;
      RECT 8.91 1.45 9.86 1.465 ;
      RECT 8.91 1.445 9.85 1.465 ;
      RECT 9.805 1.39 9.815 1.695 ;
      RECT 8.91 1.425 9.835 1.465 ;
      RECT 8.91 1.405 9.82 1.465 ;
      RECT 8.91 0.4 9.8 0.57 ;
      RECT 9.97 0.895 10.3 1.32 ;
      RECT 9.97 0.41 10.19 1.32 ;
      RECT 9.885 4.27 10.095 4.87 ;
      RECT 9.745 4.27 10.095 4.47 ;
      RECT 8.465 1.87 8.74 2.57 ;
      RECT 8.685 0.36 8.74 2.57 ;
      RECT 8.57 1.165 8.74 2.57 ;
      RECT 8.57 0.36 8.74 1.16 ;
      RECT 8.48 0.36 8.74 0.835 ;
      RECT 6.61 1.53 6.86 2.065 ;
      RECT 7.58 1.53 8.295 1.995 ;
      RECT 6.61 1.53 8.4 1.7 ;
      RECT 8.17 1.165 8.4 1.7 ;
      RECT 7.165 0.41 7.42 1.7 ;
      RECT 8.17 1.1 8.23 1.995 ;
      RECT 8.23 1.095 8.4 1.16 ;
      RECT 6.63 0.41 7.42 0.675 ;
      RECT 7.59 4.22 8.265 4.47 ;
      RECT 8 3.86 8.265 4.47 ;
      RECT 7.75 4.64 8.08 5.19 ;
      RECT 6.69 4.64 8.08 4.83 ;
      RECT 6.69 3.8 6.86 4.83 ;
      RECT 6.57 4.22 6.86 4.55 ;
      RECT 6.69 3.8 7.63 3.97 ;
      RECT 7.33 3.25 7.63 3.97 ;
      RECT 7.59 0.83 8 1.35 ;
      RECT 7.59 0.41 7.79 1.35 ;
      RECT 6.2 0.59 6.37 2.57 ;
      RECT 6.2 1.1 6.995 1.35 ;
      RECT 6.2 0.59 6.45 1.35 ;
      RECT 6.12 0.59 6.45 1.01 ;
      RECT 6.15 5 6.71 5.29 ;
      RECT 6.15 3.08 6.4 5.29 ;
      RECT 6.15 3.08 6.61 3.63 ;
      RECT 74.625 -1.03 74.795 -0.52 ;
      RECT 74.625 0.79 74.795 2.26 ;
      RECT 74.625 3.41 74.795 4.88 ;
      RECT 74.625 6.19 74.795 6.7 ;
      RECT 73.635 -1.03 73.805 -0.52 ;
      RECT 73.635 0.79 73.805 2.26 ;
      RECT 73.635 3.41 73.805 4.88 ;
      RECT 73.635 6.19 73.805 6.7 ;
      RECT 72.27 -1.03 72.44 2.26 ;
      RECT 72.27 3.41 72.44 6.7 ;
      RECT 71.84 -1.03 72.01 -0.52 ;
      RECT 71.84 0.05 72.01 2.26 ;
      RECT 71.84 3.41 72.01 5.62 ;
      RECT 71.84 6.19 72.01 6.7 ;
      RECT 70.47 0.055 70.64 1.33 ;
      RECT 70.47 4.34 70.64 5.615 ;
      RECT 68.76 1.18 69.11 1.43 ;
      RECT 67.7 4.27 68.15 4.78 ;
      RECT 66.38 2.23 66.86 2.57 ;
      RECT 65.94 4.22 66.265 4.55 ;
      RECT 65.6 0.74 66.15 1.125 ;
      RECT 64.085 2.23 64.56 2.57 ;
      RECT 63.72 4.22 64.06 4.47 ;
      RECT 62.38 1.18 62.72 2.06 ;
      RECT 60.45 -1.03 60.62 -0.52 ;
      RECT 60.45 0.79 60.62 2.26 ;
      RECT 60.45 3.41 60.62 4.88 ;
      RECT 60.45 6.19 60.62 6.7 ;
      RECT 59.46 -1.03 59.63 -0.52 ;
      RECT 59.46 0.79 59.63 2.26 ;
      RECT 59.46 3.41 59.63 4.88 ;
      RECT 59.46 6.19 59.63 6.7 ;
      RECT 58.095 -1.03 58.265 2.26 ;
      RECT 58.095 3.41 58.265 6.7 ;
      RECT 57.665 -1.03 57.835 -0.52 ;
      RECT 57.665 0.05 57.835 2.26 ;
      RECT 57.665 3.41 57.835 5.62 ;
      RECT 57.665 6.19 57.835 6.7 ;
      RECT 56.295 0.055 56.465 1.33 ;
      RECT 56.295 4.34 56.465 5.615 ;
      RECT 54.585 1.18 54.935 1.43 ;
      RECT 53.525 4.27 53.975 4.78 ;
      RECT 52.205 2.23 52.685 2.57 ;
      RECT 51.765 4.22 52.09 4.55 ;
      RECT 51.425 0.74 51.975 1.125 ;
      RECT 49.91 2.23 50.385 2.57 ;
      RECT 49.545 4.22 49.885 4.47 ;
      RECT 48.205 1.18 48.545 2.06 ;
      RECT 46.28 -1.03 46.45 -0.52 ;
      RECT 46.28 0.79 46.45 2.26 ;
      RECT 46.28 3.41 46.45 4.88 ;
      RECT 46.28 6.19 46.45 6.7 ;
      RECT 45.29 -1.03 45.46 -0.52 ;
      RECT 45.29 0.79 45.46 2.26 ;
      RECT 45.29 3.41 45.46 4.88 ;
      RECT 45.29 6.19 45.46 6.7 ;
      RECT 43.925 -1.03 44.095 2.26 ;
      RECT 43.925 3.41 44.095 6.7 ;
      RECT 43.495 -1.03 43.665 -0.52 ;
      RECT 43.495 0.05 43.665 2.26 ;
      RECT 43.495 3.41 43.665 5.62 ;
      RECT 43.495 6.19 43.665 6.7 ;
      RECT 42.125 0.055 42.295 1.33 ;
      RECT 42.125 4.34 42.295 5.615 ;
      RECT 40.415 1.18 40.765 1.43 ;
      RECT 39.355 4.27 39.805 4.78 ;
      RECT 38.035 2.23 38.515 2.57 ;
      RECT 37.595 4.22 37.92 4.55 ;
      RECT 37.255 0.74 37.805 1.125 ;
      RECT 35.74 2.23 36.215 2.57 ;
      RECT 35.375 4.22 35.715 4.47 ;
      RECT 34.035 1.18 34.375 2.06 ;
      RECT 32.105 -1.03 32.275 -0.52 ;
      RECT 32.105 0.79 32.275 2.26 ;
      RECT 32.105 3.41 32.275 4.88 ;
      RECT 32.105 6.19 32.275 6.7 ;
      RECT 31.115 -1.03 31.285 -0.52 ;
      RECT 31.115 0.79 31.285 2.26 ;
      RECT 31.115 3.41 31.285 4.88 ;
      RECT 31.115 6.19 31.285 6.7 ;
      RECT 29.75 -1.03 29.92 2.26 ;
      RECT 29.75 3.41 29.92 6.7 ;
      RECT 29.32 -1.03 29.49 -0.52 ;
      RECT 29.32 0.05 29.49 2.26 ;
      RECT 29.32 3.41 29.49 5.62 ;
      RECT 29.32 6.19 29.49 6.7 ;
      RECT 27.95 0.055 28.12 1.33 ;
      RECT 27.95 4.34 28.12 5.615 ;
      RECT 26.24 1.18 26.59 1.43 ;
      RECT 25.18 4.27 25.63 4.78 ;
      RECT 23.86 2.23 24.34 2.57 ;
      RECT 23.42 4.22 23.745 4.55 ;
      RECT 23.08 0.74 23.63 1.125 ;
      RECT 21.565 2.23 22.04 2.57 ;
      RECT 21.2 4.22 21.54 4.47 ;
      RECT 19.86 1.18 20.2 2.06 ;
      RECT 17.935 -1.03 18.105 -0.52 ;
      RECT 17.935 0.79 18.105 2.26 ;
      RECT 17.935 3.41 18.105 4.88 ;
      RECT 17.935 6.19 18.105 6.7 ;
      RECT 16.945 -1.03 17.115 -0.52 ;
      RECT 16.945 0.79 17.115 2.26 ;
      RECT 16.945 3.41 17.115 4.88 ;
      RECT 16.945 6.19 17.115 6.7 ;
      RECT 15.58 -1.03 15.75 2.26 ;
      RECT 15.58 3.41 15.75 6.7 ;
      RECT 15.15 -1.03 15.32 -0.52 ;
      RECT 15.15 0.05 15.32 2.26 ;
      RECT 15.15 3.41 15.32 5.62 ;
      RECT 15.15 6.19 15.32 6.7 ;
      RECT 13.78 0.055 13.95 1.33 ;
      RECT 13.78 4.34 13.95 5.615 ;
      RECT 12.07 1.18 12.42 1.43 ;
      RECT 11.01 4.27 11.46 4.78 ;
      RECT 9.69 2.23 10.17 2.57 ;
      RECT 9.25 4.22 9.575 4.55 ;
      RECT 8.91 0.74 9.46 1.125 ;
      RECT 7.395 2.23 7.87 2.57 ;
      RECT 7.03 4.22 7.37 4.47 ;
      RECT 5.69 1.18 6.03 2.06 ;
  END
END sky130_osu_ring_oscillator_mpr2ca_8

MACRO sky130_osu_ring_oscillator_mpr2ct_8
  CLASS CORE ;
  ORIGIN -3.235 5.43 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ct_8 3.235 -5.43 ;
  SIZE 71.16 BY 8.89 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT 66.075 0.37 66.405 0.7 ;
      RECT 66.075 0.385 66.875 0.685 ;
      RECT 66.13 0.345 66.43 0.685 ;
      RECT 65.725 -1.665 66.055 -1.335 ;
      RECT 65.725 -1.65 66.525 -1.35 ;
      RECT 65.74 -1.695 66.04 -1.335 ;
      RECT 65.385 -2.345 65.715 -2.015 ;
      RECT 65.385 -2.33 66.185 -2.03 ;
      RECT 65.47 -2.355 65.77 -2.03 ;
      RECT 65.035 0.37 65.365 0.7 ;
      RECT 64.565 0.385 65.365 0.685 ;
      RECT 65.06 0.325 65.36 0.7 ;
      RECT 64.705 -1.265 65.035 -0.935 ;
      RECT 62.665 -1.265 62.995 -0.935 ;
      RECT 62.665 -1.25 65.035 -0.95 ;
      RECT 64.355 -2.005 64.685 -1.675 ;
      RECT 63.895 -1.99 64.695 -1.69 ;
      RECT 64.025 -3.195 64.355 -2.865 ;
      RECT 63.555 -3.18 64.355 -2.88 ;
      RECT 64.015 -3.185 64.355 -2.88 ;
      RECT 64.025 1.06 64.355 1.39 ;
      RECT 63.555 1.075 64.355 1.375 ;
      RECT 63.935 1.035 64.235 1.375 ;
      RECT 63.345 0.37 63.675 0.7 ;
      RECT 62.875 0.385 63.675 0.685 ;
      RECT 51.9 0.37 52.23 0.7 ;
      RECT 51.9 0.385 52.7 0.685 ;
      RECT 51.955 0.345 52.255 0.685 ;
      RECT 51.55 -1.665 51.88 -1.335 ;
      RECT 51.55 -1.65 52.35 -1.35 ;
      RECT 51.565 -1.695 51.865 -1.335 ;
      RECT 51.21 -2.345 51.54 -2.015 ;
      RECT 51.21 -2.33 52.01 -2.03 ;
      RECT 51.295 -2.355 51.595 -2.03 ;
      RECT 50.86 0.37 51.19 0.7 ;
      RECT 50.39 0.385 51.19 0.685 ;
      RECT 50.885 0.325 51.185 0.7 ;
      RECT 50.53 -1.265 50.86 -0.935 ;
      RECT 48.49 -1.265 48.82 -0.935 ;
      RECT 48.49 -1.25 50.86 -0.95 ;
      RECT 50.18 -2.005 50.51 -1.675 ;
      RECT 49.72 -1.99 50.52 -1.69 ;
      RECT 49.85 -3.195 50.18 -2.865 ;
      RECT 49.38 -3.18 50.18 -2.88 ;
      RECT 49.84 -3.185 50.18 -2.88 ;
      RECT 49.85 1.06 50.18 1.39 ;
      RECT 49.38 1.075 50.18 1.375 ;
      RECT 49.76 1.035 50.06 1.375 ;
      RECT 49.17 0.37 49.5 0.7 ;
      RECT 48.7 0.385 49.5 0.685 ;
      RECT 37.725 0.37 38.055 0.7 ;
      RECT 37.725 0.385 38.525 0.685 ;
      RECT 37.78 0.345 38.08 0.685 ;
      RECT 37.375 -1.665 37.705 -1.335 ;
      RECT 37.375 -1.65 38.175 -1.35 ;
      RECT 37.39 -1.695 37.69 -1.335 ;
      RECT 37.035 -2.345 37.365 -2.015 ;
      RECT 37.035 -2.33 37.835 -2.03 ;
      RECT 37.12 -2.355 37.42 -2.03 ;
      RECT 36.685 0.37 37.015 0.7 ;
      RECT 36.215 0.385 37.015 0.685 ;
      RECT 36.71 0.325 37.01 0.7 ;
      RECT 36.355 -1.265 36.685 -0.935 ;
      RECT 34.315 -1.265 34.645 -0.935 ;
      RECT 34.315 -1.25 36.685 -0.95 ;
      RECT 36.005 -2.005 36.335 -1.675 ;
      RECT 35.545 -1.99 36.345 -1.69 ;
      RECT 35.675 -3.195 36.005 -2.865 ;
      RECT 35.205 -3.18 36.005 -2.88 ;
      RECT 35.665 -3.185 36.005 -2.88 ;
      RECT 35.675 1.06 36.005 1.39 ;
      RECT 35.205 1.075 36.005 1.375 ;
      RECT 35.585 1.035 35.885 1.375 ;
      RECT 34.995 0.37 35.325 0.7 ;
      RECT 34.525 0.385 35.325 0.685 ;
      RECT 23.555 0.36 23.885 0.69 ;
      RECT 23.555 0.375 24.355 0.675 ;
      RECT 23.61 0.335 23.91 0.675 ;
      RECT 23.205 -1.675 23.535 -1.345 ;
      RECT 23.205 -1.66 24.005 -1.36 ;
      RECT 23.22 -1.705 23.52 -1.345 ;
      RECT 22.865 -2.355 23.195 -2.025 ;
      RECT 22.865 -2.34 23.665 -2.04 ;
      RECT 22.95 -2.365 23.25 -2.04 ;
      RECT 22.515 0.36 22.845 0.69 ;
      RECT 22.045 0.375 22.845 0.675 ;
      RECT 22.54 0.315 22.84 0.69 ;
      RECT 22.185 -1.275 22.515 -0.945 ;
      RECT 20.145 -1.275 20.475 -0.945 ;
      RECT 20.145 -1.26 22.515 -0.96 ;
      RECT 21.835 -2.015 22.165 -1.685 ;
      RECT 21.375 -2 22.175 -1.7 ;
      RECT 21.505 -3.205 21.835 -2.875 ;
      RECT 21.035 -3.19 21.835 -2.89 ;
      RECT 21.495 -3.195 21.835 -2.89 ;
      RECT 21.505 1.05 21.835 1.38 ;
      RECT 21.035 1.065 21.835 1.365 ;
      RECT 21.415 1.025 21.715 1.365 ;
      RECT 20.825 0.36 21.155 0.69 ;
      RECT 20.355 0.375 21.155 0.675 ;
      RECT 9.39 0.36 9.72 0.69 ;
      RECT 9.39 0.375 10.19 0.675 ;
      RECT 9.445 0.335 9.745 0.675 ;
      RECT 9.04 -1.675 9.37 -1.345 ;
      RECT 9.04 -1.66 9.84 -1.36 ;
      RECT 9.055 -1.705 9.355 -1.345 ;
      RECT 8.7 -2.355 9.03 -2.025 ;
      RECT 8.7 -2.34 9.5 -2.04 ;
      RECT 8.785 -2.365 9.085 -2.04 ;
      RECT 8.35 0.36 8.68 0.69 ;
      RECT 7.88 0.375 8.68 0.675 ;
      RECT 8.375 0.315 8.675 0.69 ;
      RECT 8.02 -1.275 8.35 -0.945 ;
      RECT 5.98 -1.275 6.31 -0.945 ;
      RECT 5.98 -1.26 8.35 -0.96 ;
      RECT 7.67 -2.015 8 -1.685 ;
      RECT 7.21 -2 8.01 -1.7 ;
      RECT 7.34 -3.205 7.67 -2.875 ;
      RECT 6.87 -3.19 7.67 -2.89 ;
      RECT 7.33 -3.195 7.67 -2.89 ;
      RECT 7.34 1.05 7.67 1.38 ;
      RECT 6.87 1.065 7.67 1.365 ;
      RECT 7.25 1.025 7.55 1.365 ;
      RECT 6.66 0.36 6.99 0.69 ;
      RECT 6.19 0.375 6.99 0.675 ;
    LAYER via2 ;
      RECT 66.14 0.435 66.34 0.635 ;
      RECT 65.79 -1.6 65.99 -1.4 ;
      RECT 65.45 -2.28 65.65 -2.08 ;
      RECT 65.1 0.435 65.3 0.635 ;
      RECT 64.77 -1.2 64.97 -1 ;
      RECT 64.42 -1.94 64.62 -1.74 ;
      RECT 64.09 -3.13 64.29 -2.93 ;
      RECT 64.09 1.125 64.29 1.325 ;
      RECT 63.41 0.435 63.61 0.635 ;
      RECT 62.73 -1.2 62.93 -1 ;
      RECT 51.965 0.435 52.165 0.635 ;
      RECT 51.615 -1.6 51.815 -1.4 ;
      RECT 51.275 -2.28 51.475 -2.08 ;
      RECT 50.925 0.435 51.125 0.635 ;
      RECT 50.595 -1.2 50.795 -1 ;
      RECT 50.245 -1.94 50.445 -1.74 ;
      RECT 49.915 -3.13 50.115 -2.93 ;
      RECT 49.915 1.125 50.115 1.325 ;
      RECT 49.235 0.435 49.435 0.635 ;
      RECT 48.555 -1.2 48.755 -1 ;
      RECT 37.79 0.435 37.99 0.635 ;
      RECT 37.44 -1.6 37.64 -1.4 ;
      RECT 37.1 -2.28 37.3 -2.08 ;
      RECT 36.75 0.435 36.95 0.635 ;
      RECT 36.42 -1.2 36.62 -1 ;
      RECT 36.07 -1.94 36.27 -1.74 ;
      RECT 35.74 -3.13 35.94 -2.93 ;
      RECT 35.74 1.125 35.94 1.325 ;
      RECT 35.06 0.435 35.26 0.635 ;
      RECT 34.38 -1.2 34.58 -1 ;
      RECT 23.62 0.425 23.82 0.625 ;
      RECT 23.27 -1.61 23.47 -1.41 ;
      RECT 22.93 -2.29 23.13 -2.09 ;
      RECT 22.58 0.425 22.78 0.625 ;
      RECT 22.25 -1.21 22.45 -1.01 ;
      RECT 21.9 -1.95 22.1 -1.75 ;
      RECT 21.57 -3.14 21.77 -2.94 ;
      RECT 21.57 1.115 21.77 1.315 ;
      RECT 20.89 0.425 21.09 0.625 ;
      RECT 20.21 -1.21 20.41 -1.01 ;
      RECT 9.455 0.425 9.655 0.625 ;
      RECT 9.105 -1.61 9.305 -1.41 ;
      RECT 8.765 -2.29 8.965 -2.09 ;
      RECT 8.415 0.425 8.615 0.625 ;
      RECT 8.085 -1.21 8.285 -1.01 ;
      RECT 7.735 -1.95 7.935 -1.75 ;
      RECT 7.405 -3.14 7.605 -2.94 ;
      RECT 7.405 1.115 7.605 1.315 ;
      RECT 6.725 0.425 6.925 0.625 ;
      RECT 6.045 -1.21 6.245 -1.01 ;
    LAYER met2 ;
      RECT 13.98 0.85 14.3 1.175 ;
      RECT 14.01 0.265 14.18 1.175 ;
      RECT 14.01 0.265 14.185 0.615 ;
      RECT 14.01 0.265 14.985 0.44 ;
      RECT 14.81 -3.465 14.985 0.44 ;
      RECT 12.31 -3.435 12.635 -3.11 ;
      RECT 14.755 -3.465 15.105 -3.115 ;
      RECT 12.31 -3.405 15.105 -3.235 ;
      RECT 12.375 -5.17 12.54 -3.11 ;
      RECT 73.81 -4.325 74.16 -3.975 ;
      RECT 73.845 -5.17 74.01 -3.975 ;
      RECT 12.375 -5.17 74.01 -5.005 ;
      RECT 70.665 0.86 70.985 1.185 ;
      RECT 70.695 0.275 70.865 1.185 ;
      RECT 70.695 0.275 70.87 0.625 ;
      RECT 70.695 0.275 71.67 0.45 ;
      RECT 71.495 -3.455 71.67 0.45 ;
      RECT 68.995 -3.425 69.32 -3.1 ;
      RECT 71.44 -3.455 71.79 -3.105 ;
      RECT 68.995 -3.395 71.79 -3.225 ;
      RECT 69.07 -4.295 69.21 -3.1 ;
      RECT 59.65 -4.325 60 -3.975 ;
      RECT 59.65 -4.295 69.21 -4.155 ;
      RECT 71.465 1.235 71.79 1.56 ;
      RECT 70.35 1.325 71.79 1.495 ;
      RECT 70.35 -3.025 70.51 1.495 ;
      RECT 68.525 -2.365 70.51 -2.19 ;
      RECT 68.525 -3.075 68.7 -2.19 ;
      RECT 70.665 -3.055 70.985 -2.735 ;
      RECT 64.05 -3.215 64.33 -2.845 ;
      RECT 70.35 -3.025 70.985 -2.855 ;
      RECT 64.05 -3.075 68.7 -2.9 ;
      RECT 69.62 0.435 69.945 0.76 ;
      RECT 69.69 -1.925 69.86 0.76 ;
      RECT 69.62 -1.925 69.945 -1.6 ;
      RECT 63.39 1.875 68.91 2.04 ;
      RECT 68.745 -1.605 68.91 2.04 ;
      RECT 63.39 0.35 63.555 2.04 ;
      RECT 63.37 0.35 63.65 0.72 ;
      RECT 68.91 -1.765 69.235 -1.44 ;
      RECT 67.12 1.06 67.38 1.38 ;
      RECT 67.18 -2.68 67.32 1.38 ;
      RECT 67.12 -2.68 67.38 -2.36 ;
      RECT 66.44 -0.64 66.7 -0.32 ;
      RECT 66.5 -1.66 66.64 -0.32 ;
      RECT 66.44 -1.66 66.7 -1.34 ;
      RECT 65.42 1.06 65.68 1.38 ;
      RECT 65.48 -0.21 65.62 1.38 ;
      RECT 64.8 -0.21 65.62 -0.07 ;
      RECT 64.8 -2.68 64.94 -0.07 ;
      RECT 64.73 -1.285 65.01 -0.915 ;
      RECT 64.74 -2.68 65 -2.36 ;
      RECT 62.69 -1.285 62.97 -0.915 ;
      RECT 62.76 -3.02 62.9 -0.915 ;
      RECT 62.7 -3.02 62.96 -2.7 ;
      RECT 62.02 -0.64 62.28 -0.32 ;
      RECT 62.08 -2.68 62.22 -0.32 ;
      RECT 62.02 -2.68 62.28 -2.36 ;
      RECT 56.49 0.86 56.81 1.185 ;
      RECT 56.52 0.275 56.69 1.185 ;
      RECT 56.52 0.275 56.695 0.625 ;
      RECT 56.52 0.275 57.495 0.45 ;
      RECT 57.32 -3.455 57.495 0.45 ;
      RECT 54.82 -3.425 55.145 -3.1 ;
      RECT 57.265 -3.455 57.615 -3.105 ;
      RECT 54.82 -3.395 57.615 -3.225 ;
      RECT 54.945 -4.295 55.095 -3.1 ;
      RECT 45.47 -4.325 45.82 -3.975 ;
      RECT 45.47 -4.295 55.095 -4.145 ;
      RECT 57.29 1.235 57.615 1.56 ;
      RECT 56.175 1.325 57.615 1.495 ;
      RECT 56.175 -3.025 56.335 1.495 ;
      RECT 54.35 -2.365 56.335 -2.19 ;
      RECT 54.35 -3.075 54.525 -2.19 ;
      RECT 56.49 -3.055 56.81 -2.735 ;
      RECT 49.875 -3.215 50.155 -2.845 ;
      RECT 56.175 -3.025 56.81 -2.855 ;
      RECT 49.875 -3.075 54.525 -2.9 ;
      RECT 55.445 0.435 55.77 0.76 ;
      RECT 55.515 -1.925 55.685 0.76 ;
      RECT 55.445 -1.925 55.77 -1.6 ;
      RECT 49.215 1.875 54.735 2.04 ;
      RECT 54.57 -1.605 54.735 2.04 ;
      RECT 49.215 0.35 49.38 2.04 ;
      RECT 49.195 0.35 49.475 0.72 ;
      RECT 54.735 -1.765 55.06 -1.44 ;
      RECT 52.945 1.06 53.205 1.38 ;
      RECT 53.005 -2.68 53.145 1.38 ;
      RECT 52.945 -2.68 53.205 -2.36 ;
      RECT 52.265 -0.64 52.525 -0.32 ;
      RECT 52.325 -1.66 52.465 -0.32 ;
      RECT 52.265 -1.66 52.525 -1.34 ;
      RECT 51.245 1.06 51.505 1.38 ;
      RECT 51.305 -0.21 51.445 1.38 ;
      RECT 50.625 -0.21 51.445 -0.07 ;
      RECT 50.625 -2.68 50.765 -0.07 ;
      RECT 50.555 -1.285 50.835 -0.915 ;
      RECT 50.565 -2.68 50.825 -2.36 ;
      RECT 48.515 -1.285 48.795 -0.915 ;
      RECT 48.585 -3.02 48.725 -0.915 ;
      RECT 48.525 -3.02 48.785 -2.7 ;
      RECT 47.845 -0.64 48.105 -0.32 ;
      RECT 47.905 -2.68 48.045 -0.32 ;
      RECT 47.845 -2.68 48.105 -2.36 ;
      RECT 42.315 0.86 42.635 1.185 ;
      RECT 42.345 0.275 42.515 1.185 ;
      RECT 42.345 0.275 42.52 0.625 ;
      RECT 42.345 0.275 43.32 0.45 ;
      RECT 43.145 -3.455 43.32 0.45 ;
      RECT 40.645 -3.425 40.97 -3.1 ;
      RECT 43.09 -3.455 43.44 -3.105 ;
      RECT 40.645 -3.395 43.44 -3.225 ;
      RECT 40.76 -4.3 40.9 -3.1 ;
      RECT 31.31 -4.33 31.66 -3.98 ;
      RECT 31.31 -4.3 40.9 -4.16 ;
      RECT 43.115 1.235 43.44 1.56 ;
      RECT 42 1.325 43.44 1.495 ;
      RECT 42 -3.025 42.16 1.495 ;
      RECT 40.175 -2.365 42.16 -2.19 ;
      RECT 40.175 -3.075 40.35 -2.19 ;
      RECT 42.315 -3.055 42.635 -2.735 ;
      RECT 35.7 -3.215 35.98 -2.845 ;
      RECT 42 -3.025 42.635 -2.855 ;
      RECT 35.7 -3.075 40.35 -2.9 ;
      RECT 41.27 0.435 41.595 0.76 ;
      RECT 41.34 -1.925 41.51 0.76 ;
      RECT 41.27 -1.925 41.595 -1.6 ;
      RECT 35.04 1.875 40.56 2.04 ;
      RECT 40.395 -1.605 40.56 2.04 ;
      RECT 35.04 0.35 35.205 2.04 ;
      RECT 35.02 0.35 35.3 0.72 ;
      RECT 40.56 -1.765 40.885 -1.44 ;
      RECT 38.77 1.06 39.03 1.38 ;
      RECT 38.83 -2.68 38.97 1.38 ;
      RECT 38.77 -2.68 39.03 -2.36 ;
      RECT 38.09 -0.64 38.35 -0.32 ;
      RECT 38.15 -1.66 38.29 -0.32 ;
      RECT 38.09 -1.66 38.35 -1.34 ;
      RECT 37.07 1.06 37.33 1.38 ;
      RECT 37.13 -0.21 37.27 1.38 ;
      RECT 36.45 -0.21 37.27 -0.07 ;
      RECT 36.45 -2.68 36.59 -0.07 ;
      RECT 36.38 -1.285 36.66 -0.915 ;
      RECT 36.39 -2.68 36.65 -2.36 ;
      RECT 34.34 -1.285 34.62 -0.915 ;
      RECT 34.41 -3.02 34.55 -0.915 ;
      RECT 34.35 -3.02 34.61 -2.7 ;
      RECT 33.67 -0.64 33.93 -0.32 ;
      RECT 33.73 -2.68 33.87 -0.32 ;
      RECT 33.67 -2.68 33.93 -2.36 ;
      RECT 28.145 0.85 28.465 1.175 ;
      RECT 28.175 0.265 28.345 1.175 ;
      RECT 28.175 0.265 28.35 0.615 ;
      RECT 28.175 0.265 29.15 0.44 ;
      RECT 28.975 -3.465 29.15 0.44 ;
      RECT 26.475 -3.435 26.8 -3.11 ;
      RECT 28.92 -3.465 29.27 -3.115 ;
      RECT 26.475 -3.405 29.27 -3.235 ;
      RECT 26.595 -4.3 26.735 -3.11 ;
      RECT 17.14 -4.33 17.49 -3.98 ;
      RECT 17.14 -4.3 26.735 -4.16 ;
      RECT 28.945 1.225 29.27 1.55 ;
      RECT 27.83 1.315 29.27 1.485 ;
      RECT 27.83 -3.035 27.99 1.485 ;
      RECT 26.005 -2.375 27.99 -2.2 ;
      RECT 26.005 -3.085 26.18 -2.2 ;
      RECT 28.145 -3.065 28.465 -2.745 ;
      RECT 21.53 -3.225 21.81 -2.855 ;
      RECT 27.83 -3.035 28.465 -2.865 ;
      RECT 21.53 -3.085 26.18 -2.91 ;
      RECT 27.1 0.425 27.425 0.75 ;
      RECT 27.17 -1.935 27.34 0.75 ;
      RECT 27.1 -1.935 27.425 -1.61 ;
      RECT 20.87 1.865 26.39 2.03 ;
      RECT 26.225 -1.615 26.39 2.03 ;
      RECT 20.87 0.34 21.035 2.03 ;
      RECT 20.85 0.34 21.13 0.71 ;
      RECT 26.39 -1.775 26.715 -1.45 ;
      RECT 24.6 1.05 24.86 1.37 ;
      RECT 24.66 -2.69 24.8 1.37 ;
      RECT 24.6 -2.69 24.86 -2.37 ;
      RECT 23.92 -0.65 24.18 -0.33 ;
      RECT 23.98 -1.67 24.12 -0.33 ;
      RECT 23.92 -1.67 24.18 -1.35 ;
      RECT 22.9 1.05 23.16 1.37 ;
      RECT 22.96 -0.22 23.1 1.37 ;
      RECT 22.28 -0.22 23.1 -0.08 ;
      RECT 22.28 -2.69 22.42 -0.08 ;
      RECT 22.21 -1.295 22.49 -0.925 ;
      RECT 22.22 -2.69 22.48 -2.37 ;
      RECT 20.17 -1.295 20.45 -0.925 ;
      RECT 20.24 -3.03 20.38 -0.925 ;
      RECT 20.18 -3.03 20.44 -2.71 ;
      RECT 19.5 -0.65 19.76 -0.33 ;
      RECT 19.56 -2.69 19.7 -0.33 ;
      RECT 19.5 -2.69 19.76 -2.37 ;
      RECT 14.78 1.225 15.105 1.55 ;
      RECT 13.665 1.315 15.105 1.485 ;
      RECT 13.665 -3.035 13.825 1.485 ;
      RECT 11.84 -2.375 13.825 -2.2 ;
      RECT 11.84 -3.085 12.015 -2.2 ;
      RECT 13.98 -3.065 14.3 -2.745 ;
      RECT 7.365 -3.225 7.645 -2.855 ;
      RECT 13.665 -3.035 14.3 -2.865 ;
      RECT 7.365 -3.085 12.015 -2.91 ;
      RECT 12.935 0.425 13.26 0.75 ;
      RECT 13.005 -1.935 13.175 0.75 ;
      RECT 12.935 -1.935 13.26 -1.61 ;
      RECT 6.705 1.865 12.225 2.03 ;
      RECT 12.06 -1.615 12.225 2.03 ;
      RECT 6.705 0.34 6.87 2.03 ;
      RECT 6.685 0.34 6.965 0.71 ;
      RECT 12.225 -1.775 12.55 -1.45 ;
      RECT 10.435 1.05 10.695 1.37 ;
      RECT 10.495 -2.69 10.635 1.37 ;
      RECT 10.435 -2.69 10.695 -2.37 ;
      RECT 9.755 -0.65 10.015 -0.33 ;
      RECT 9.815 -1.67 9.955 -0.33 ;
      RECT 9.755 -1.67 10.015 -1.35 ;
      RECT 8.735 1.05 8.995 1.37 ;
      RECT 8.795 -0.22 8.935 1.37 ;
      RECT 8.115 -0.22 8.935 -0.08 ;
      RECT 8.115 -2.69 8.255 -0.08 ;
      RECT 8.045 -1.295 8.325 -0.925 ;
      RECT 8.055 -2.69 8.315 -2.37 ;
      RECT 6.005 -1.295 6.285 -0.925 ;
      RECT 6.075 -3.03 6.215 -0.925 ;
      RECT 6.015 -3.03 6.275 -2.71 ;
      RECT 5.335 -0.65 5.595 -0.33 ;
      RECT 5.395 -2.69 5.535 -0.33 ;
      RECT 5.335 -2.69 5.595 -2.37 ;
      RECT 66.1 0.35 66.38 0.72 ;
      RECT 65.75 -1.685 66.03 -1.315 ;
      RECT 65.41 -2.365 65.69 -1.995 ;
      RECT 65.06 0.35 65.34 0.72 ;
      RECT 64.38 -2.025 64.66 -1.655 ;
      RECT 64.05 1.04 64.33 1.41 ;
      RECT 51.925 0.35 52.205 0.72 ;
      RECT 51.575 -1.685 51.855 -1.315 ;
      RECT 51.235 -2.365 51.515 -1.995 ;
      RECT 50.885 0.35 51.165 0.72 ;
      RECT 50.205 -2.025 50.485 -1.655 ;
      RECT 49.875 1.04 50.155 1.41 ;
      RECT 37.75 0.35 38.03 0.72 ;
      RECT 37.4 -1.685 37.68 -1.315 ;
      RECT 37.06 -2.365 37.34 -1.995 ;
      RECT 36.71 0.35 36.99 0.72 ;
      RECT 36.03 -2.025 36.31 -1.655 ;
      RECT 35.7 1.04 35.98 1.41 ;
      RECT 23.58 0.34 23.86 0.71 ;
      RECT 23.23 -1.695 23.51 -1.325 ;
      RECT 22.89 -2.375 23.17 -2.005 ;
      RECT 22.54 0.34 22.82 0.71 ;
      RECT 21.86 -2.035 22.14 -1.665 ;
      RECT 21.53 1.03 21.81 1.4 ;
      RECT 9.415 0.34 9.695 0.71 ;
      RECT 9.065 -1.695 9.345 -1.325 ;
      RECT 8.725 -2.375 9.005 -2.005 ;
      RECT 8.375 0.34 8.655 0.71 ;
      RECT 7.695 -2.035 7.975 -1.665 ;
      RECT 7.365 1.03 7.645 1.4 ;
    LAYER via1 ;
      RECT 73.91 -4.225 74.06 -4.075 ;
      RECT 71.555 1.32 71.705 1.47 ;
      RECT 71.54 -3.355 71.69 -3.205 ;
      RECT 70.75 -2.97 70.9 -2.82 ;
      RECT 70.75 0.95 70.9 1.1 ;
      RECT 69.71 -1.84 69.86 -1.69 ;
      RECT 69.71 0.52 69.86 0.67 ;
      RECT 69.085 -3.34 69.235 -3.19 ;
      RECT 69 -1.68 69.15 -1.53 ;
      RECT 67.175 -2.595 67.325 -2.445 ;
      RECT 67.175 1.145 67.325 1.295 ;
      RECT 66.495 -1.575 66.645 -1.425 ;
      RECT 66.495 -0.555 66.645 -0.405 ;
      RECT 66.155 0.465 66.305 0.615 ;
      RECT 65.815 -1.575 65.965 -1.425 ;
      RECT 65.475 -2.255 65.625 -2.105 ;
      RECT 65.475 1.145 65.625 1.295 ;
      RECT 65.125 0.465 65.275 0.615 ;
      RECT 64.795 -2.595 64.945 -2.445 ;
      RECT 64.455 -1.915 64.605 -1.765 ;
      RECT 64.115 -3.105 64.265 -2.955 ;
      RECT 64.115 1.145 64.265 1.295 ;
      RECT 63.435 0.465 63.585 0.615 ;
      RECT 62.755 -2.935 62.905 -2.785 ;
      RECT 62.075 -2.595 62.225 -2.445 ;
      RECT 62.075 -0.555 62.225 -0.405 ;
      RECT 59.75 -4.225 59.9 -4.075 ;
      RECT 57.38 1.32 57.53 1.47 ;
      RECT 57.365 -3.355 57.515 -3.205 ;
      RECT 56.575 -2.97 56.725 -2.82 ;
      RECT 56.575 0.95 56.725 1.1 ;
      RECT 55.535 -1.84 55.685 -1.69 ;
      RECT 55.535 0.52 55.685 0.67 ;
      RECT 54.91 -3.34 55.06 -3.19 ;
      RECT 54.825 -1.68 54.975 -1.53 ;
      RECT 53 -2.595 53.15 -2.445 ;
      RECT 53 1.145 53.15 1.295 ;
      RECT 52.32 -1.575 52.47 -1.425 ;
      RECT 52.32 -0.555 52.47 -0.405 ;
      RECT 51.98 0.465 52.13 0.615 ;
      RECT 51.64 -1.575 51.79 -1.425 ;
      RECT 51.3 -2.255 51.45 -2.105 ;
      RECT 51.3 1.145 51.45 1.295 ;
      RECT 50.95 0.465 51.1 0.615 ;
      RECT 50.62 -2.595 50.77 -2.445 ;
      RECT 50.28 -1.915 50.43 -1.765 ;
      RECT 49.94 -3.105 50.09 -2.955 ;
      RECT 49.94 1.145 50.09 1.295 ;
      RECT 49.26 0.465 49.41 0.615 ;
      RECT 48.58 -2.935 48.73 -2.785 ;
      RECT 47.9 -2.595 48.05 -2.445 ;
      RECT 47.9 -0.555 48.05 -0.405 ;
      RECT 45.57 -4.225 45.72 -4.075 ;
      RECT 43.205 1.32 43.355 1.47 ;
      RECT 43.19 -3.355 43.34 -3.205 ;
      RECT 42.4 -2.97 42.55 -2.82 ;
      RECT 42.4 0.95 42.55 1.1 ;
      RECT 41.36 -1.84 41.51 -1.69 ;
      RECT 41.36 0.52 41.51 0.67 ;
      RECT 40.735 -3.34 40.885 -3.19 ;
      RECT 40.65 -1.68 40.8 -1.53 ;
      RECT 38.825 -2.595 38.975 -2.445 ;
      RECT 38.825 1.145 38.975 1.295 ;
      RECT 38.145 -1.575 38.295 -1.425 ;
      RECT 38.145 -0.555 38.295 -0.405 ;
      RECT 37.805 0.465 37.955 0.615 ;
      RECT 37.465 -1.575 37.615 -1.425 ;
      RECT 37.125 -2.255 37.275 -2.105 ;
      RECT 37.125 1.145 37.275 1.295 ;
      RECT 36.775 0.465 36.925 0.615 ;
      RECT 36.445 -2.595 36.595 -2.445 ;
      RECT 36.105 -1.915 36.255 -1.765 ;
      RECT 35.765 -3.105 35.915 -2.955 ;
      RECT 35.765 1.145 35.915 1.295 ;
      RECT 35.085 0.465 35.235 0.615 ;
      RECT 34.405 -2.935 34.555 -2.785 ;
      RECT 33.725 -2.595 33.875 -2.445 ;
      RECT 33.725 -0.555 33.875 -0.405 ;
      RECT 31.41 -4.23 31.56 -4.08 ;
      RECT 29.035 1.31 29.185 1.46 ;
      RECT 29.02 -3.365 29.17 -3.215 ;
      RECT 28.23 -2.98 28.38 -2.83 ;
      RECT 28.23 0.94 28.38 1.09 ;
      RECT 27.19 -1.85 27.34 -1.7 ;
      RECT 27.19 0.51 27.34 0.66 ;
      RECT 26.565 -3.35 26.715 -3.2 ;
      RECT 26.48 -1.69 26.63 -1.54 ;
      RECT 24.655 -2.605 24.805 -2.455 ;
      RECT 24.655 1.135 24.805 1.285 ;
      RECT 23.975 -1.585 24.125 -1.435 ;
      RECT 23.975 -0.565 24.125 -0.415 ;
      RECT 23.635 0.455 23.785 0.605 ;
      RECT 23.295 -1.585 23.445 -1.435 ;
      RECT 22.955 -2.265 23.105 -2.115 ;
      RECT 22.955 1.135 23.105 1.285 ;
      RECT 22.605 0.455 22.755 0.605 ;
      RECT 22.275 -2.605 22.425 -2.455 ;
      RECT 21.935 -1.925 22.085 -1.775 ;
      RECT 21.595 -3.115 21.745 -2.965 ;
      RECT 21.595 1.135 21.745 1.285 ;
      RECT 20.915 0.455 21.065 0.605 ;
      RECT 20.235 -2.945 20.385 -2.795 ;
      RECT 19.555 -2.605 19.705 -2.455 ;
      RECT 19.555 -0.565 19.705 -0.415 ;
      RECT 17.24 -4.23 17.39 -4.08 ;
      RECT 14.87 1.31 15.02 1.46 ;
      RECT 14.855 -3.365 15.005 -3.215 ;
      RECT 14.065 -2.98 14.215 -2.83 ;
      RECT 14.065 0.94 14.215 1.09 ;
      RECT 13.025 -1.85 13.175 -1.7 ;
      RECT 13.025 0.51 13.175 0.66 ;
      RECT 12.4 -3.35 12.55 -3.2 ;
      RECT 12.315 -1.69 12.465 -1.54 ;
      RECT 10.49 -2.605 10.64 -2.455 ;
      RECT 10.49 1.135 10.64 1.285 ;
      RECT 9.81 -1.585 9.96 -1.435 ;
      RECT 9.81 -0.565 9.96 -0.415 ;
      RECT 9.47 0.455 9.62 0.605 ;
      RECT 9.13 -1.585 9.28 -1.435 ;
      RECT 8.79 -2.265 8.94 -2.115 ;
      RECT 8.79 1.135 8.94 1.285 ;
      RECT 8.44 0.455 8.59 0.605 ;
      RECT 8.11 -2.605 8.26 -2.455 ;
      RECT 7.77 -1.925 7.92 -1.775 ;
      RECT 7.43 -3.115 7.58 -2.965 ;
      RECT 7.43 1.135 7.58 1.285 ;
      RECT 6.75 0.455 6.9 0.605 ;
      RECT 6.07 -2.945 6.22 -2.795 ;
      RECT 5.39 -2.605 5.54 -2.455 ;
      RECT 5.39 -0.565 5.54 -0.415 ;
    LAYER met1 ;
      RECT 60.96 -5.42 68.32 -3.47 ;
      RECT 46.785 -5.42 54.145 -3.47 ;
      RECT 32.61 -5.42 39.97 -3.47 ;
      RECT 18.44 -5.43 25.8 -3.48 ;
      RECT 4.275 -5.43 11.635 -3.48 ;
      RECT 60.96 -5.42 68.615 -3.625 ;
      RECT 46.785 -5.42 54.44 -3.625 ;
      RECT 32.61 -5.42 40.265 -3.625 ;
      RECT 18.44 -5.43 26.095 -3.635 ;
      RECT 4.275 -5.43 11.93 -3.635 ;
      RECT 60.955 -5.42 68.615 -3.785 ;
      RECT 46.78 -5.42 54.44 -3.785 ;
      RECT 32.605 -5.42 40.265 -3.785 ;
      RECT 18.435 -5.43 26.095 -3.795 ;
      RECT 4.27 -5.43 11.93 -3.795 ;
      RECT 31.575 -5.42 74.395 -5.115 ;
      RECT 3.24 -5.43 31.875 -5.125 ;
      RECT 68.41 -1.285 74.395 -0.675 ;
      RECT 54.235 -1.285 60.22 -0.675 ;
      RECT 40.06 -1.285 46.045 -0.675 ;
      RECT 54.235 -1.23 61.335 -0.68 ;
      RECT 40.06 -1.23 47.16 -0.68 ;
      RECT 31.575 -1.23 32.985 -0.68 ;
      RECT 25.89 -1.23 32.985 -0.685 ;
      RECT 11.725 -1.295 17.71 -0.685 ;
      RECT 11.725 -1.24 18.815 -0.69 ;
      RECT 3.24 -1.24 4.65 -0.69 ;
      RECT 25.89 -1.23 74.395 -0.75 ;
      RECT 68.405 -1.285 74.395 -0.75 ;
      RECT 25.885 -1.295 31.875 -0.76 ;
      RECT 54.23 -1.285 61.315 -0.75 ;
      RECT 59.925 -1.29 61.315 -0.68 ;
      RECT 40.055 -1.285 47.14 -0.75 ;
      RECT 45.75 -1.29 47.14 -0.68 ;
      RECT 3.24 -1.24 32.965 -0.76 ;
      RECT 31.575 -1.29 32.965 -0.68 ;
      RECT 11.72 -1.295 18.795 -0.76 ;
      RECT 17.405 -1.3 18.795 -0.69 ;
      RECT 3.24 -1.3 4.63 -0.69 ;
      RECT 31.575 3.155 74.395 3.46 ;
      RECT 3.24 3.145 31.875 3.45 ;
      RECT 61.23 1.76 68.43 3.46 ;
      RECT 47.055 1.76 54.255 3.46 ;
      RECT 32.88 1.76 40.08 3.46 ;
      RECT 18.71 1.75 25.91 3.45 ;
      RECT 4.545 1.75 11.745 3.45 ;
      RECT 60.96 1.49 68.32 1.97 ;
      RECT 46.785 1.49 54.145 1.97 ;
      RECT 32.61 1.49 39.97 1.97 ;
      RECT 18.44 1.48 25.8 1.96 ;
      RECT 4.275 1.48 11.635 1.96 ;
      RECT 73.795 -3.055 74.085 -2.825 ;
      RECT 73.855 -4.535 74.025 -2.825 ;
      RECT 73.81 -4.325 74.16 -3.975 ;
      RECT 73.795 -4.535 74.085 -4.305 ;
      RECT 73.795 2.345 74.085 2.575 ;
      RECT 73.855 0.865 74.025 2.575 ;
      RECT 73.795 0.865 74.085 1.095 ;
      RECT 73.385 -2.685 73.715 -2.455 ;
      RECT 73.385 -2.655 73.885 -2.485 ;
      RECT 73.385 -3.025 73.575 -2.455 ;
      RECT 72.805 -3.055 73.095 -2.825 ;
      RECT 72.805 -3.025 73.575 -2.855 ;
      RECT 72.865 -4.535 73.035 -2.825 ;
      RECT 72.805 -4.535 73.095 -4.305 ;
      RECT 72.805 2.345 73.095 2.575 ;
      RECT 72.865 0.865 73.035 2.575 ;
      RECT 72.805 0.865 73.095 1.095 ;
      RECT 72.805 0.905 73.655 1.065 ;
      RECT 73.485 0.495 73.655 1.065 ;
      RECT 72.805 0.9 73.195 1.065 ;
      RECT 73.425 0.495 73.715 0.725 ;
      RECT 73.425 0.525 73.885 0.695 ;
      RECT 72.435 -2.685 72.725 -2.455 ;
      RECT 72.435 -2.655 72.895 -2.485 ;
      RECT 72.495 -3.765 72.66 -2.455 ;
      RECT 71.01 -3.795 71.3 -3.565 ;
      RECT 71.01 -3.765 72.66 -3.595 ;
      RECT 71.07 -4.535 71.24 -3.565 ;
      RECT 71.01 -4.535 71.3 -4.305 ;
      RECT 71.01 2.345 71.3 2.575 ;
      RECT 71.07 1.605 71.24 2.575 ;
      RECT 71.07 1.7 72.66 1.87 ;
      RECT 72.49 0.495 72.66 1.87 ;
      RECT 71.01 1.605 71.3 1.835 ;
      RECT 72.435 0.495 72.725 0.725 ;
      RECT 72.435 0.525 72.895 0.695 ;
      RECT 71.44 -3.455 71.79 -3.105 ;
      RECT 71.27 -3.395 71.79 -3.225 ;
      RECT 71.465 1.235 71.79 1.56 ;
      RECT 71.44 1.235 71.79 1.465 ;
      RECT 71.27 1.265 71.79 1.435 ;
      RECT 70.665 -3.055 70.985 -2.735 ;
      RECT 70.635 -3.055 70.985 -2.825 ;
      RECT 70.35 -3.025 70.985 -2.855 ;
      RECT 70.665 0.86 70.985 1.185 ;
      RECT 70.635 0.865 70.985 1.095 ;
      RECT 70.465 0.895 70.985 1.065 ;
      RECT 69.62 -1.925 69.945 -1.6 ;
      RECT 69.7 -2.685 69.87 -1.6 ;
      RECT 69.64 -2.685 69.93 -2.455 ;
      RECT 69.64 -2.655 70.1 -2.485 ;
      RECT 69.62 0.435 69.945 0.76 ;
      RECT 69.62 0.525 70.1 0.695 ;
      RECT 68.91 -1.765 69.235 -1.44 ;
      RECT 69.035 -3.425 69.2 -1.44 ;
      RECT 68.995 -3.425 69.32 -3.1 ;
      RECT 66.41 -1.63 66.73 -1.37 ;
      RECT 67.445 -1.615 67.735 -1.385 ;
      RECT 66.41 -1.57 67.735 -1.43 ;
      RECT 66.07 0.41 66.39 0.67 ;
      RECT 67.445 0.425 67.735 0.655 ;
      RECT 67.52 0.13 67.66 0.655 ;
      RECT 66.16 0.13 66.3 0.67 ;
      RECT 66.16 0.13 67.66 0.27 ;
      RECT 67.09 -2.65 67.41 -2.39 ;
      RECT 66.815 -2.59 67.41 -2.45 ;
      RECT 64.03 1.09 64.35 1.35 ;
      RECT 63.025 1.105 63.315 1.335 ;
      RECT 63.025 1.15 64.94 1.29 ;
      RECT 64.8 0.81 64.94 1.29 ;
      RECT 64.8 0.81 66.81 0.95 ;
      RECT 66.67 0.425 66.81 0.95 ;
      RECT 66.595 0.425 66.885 0.655 ;
      RECT 66.41 -0.61 66.73 -0.35 ;
      RECT 64.265 -0.595 64.555 -0.365 ;
      RECT 64.265 -0.55 66.73 -0.41 ;
      RECT 65.73 -1.63 66.05 -1.37 ;
      RECT 63.365 -1.615 63.655 -1.385 ;
      RECT 63.365 -1.57 66.05 -1.43 ;
      RECT 65.39 1.09 65.71 1.35 ;
      RECT 65.39 1.15 65.985 1.29 ;
      RECT 65.39 -2.31 65.71 -2.05 ;
      RECT 65.115 -2.25 65.71 -2.11 ;
      RECT 64.71 -2.65 65.03 -2.39 ;
      RECT 64.435 -2.59 65.03 -2.45 ;
      RECT 64.37 -1.97 64.69 -1.71 ;
      RECT 61.495 -1.955 61.785 -1.725 ;
      RECT 61.495 -1.91 64.69 -1.77 ;
      RECT 63.95 -2.63 64.09 -1.77 ;
      RECT 63.875 -2.63 64.165 -2.4 ;
      RECT 64.03 -3.16 64.35 -2.9 ;
      RECT 64.03 -3.145 64.535 -2.915 ;
      RECT 63.94 -3.1 64.535 -2.96 ;
      RECT 63.35 0.41 63.67 0.67 ;
      RECT 60.985 0.425 61.275 0.655 ;
      RECT 60.985 0.47 63.67 0.61 ;
      RECT 63.365 -2.63 63.655 -2.4 ;
      RECT 62.76 -2.585 63.655 -2.445 ;
      RECT 62.76 -2.99 62.9 -2.445 ;
      RECT 62.67 -2.99 62.99 -2.73 ;
      RECT 61.99 -2.65 62.31 -2.39 ;
      RECT 61.715 -2.59 62.31 -2.45 ;
      RECT 61.99 -0.61 62.31 -0.35 ;
      RECT 61.715 -0.55 62.31 -0.41 ;
      RECT 59.62 -3.055 59.91 -2.825 ;
      RECT 59.68 -4.535 59.85 -2.825 ;
      RECT 59.65 -4.325 60 -3.975 ;
      RECT 59.62 -4.535 59.91 -4.305 ;
      RECT 59.62 2.345 59.91 2.575 ;
      RECT 59.68 0.865 59.85 2.575 ;
      RECT 59.62 0.865 59.91 1.095 ;
      RECT 59.21 -2.685 59.54 -2.455 ;
      RECT 59.21 -2.655 59.71 -2.485 ;
      RECT 59.21 -3.025 59.4 -2.455 ;
      RECT 58.63 -3.055 58.92 -2.825 ;
      RECT 58.63 -3.025 59.4 -2.855 ;
      RECT 58.69 -4.535 58.86 -2.825 ;
      RECT 58.63 -4.535 58.92 -4.305 ;
      RECT 58.63 2.345 58.92 2.575 ;
      RECT 58.69 0.865 58.86 2.575 ;
      RECT 58.63 0.865 58.92 1.095 ;
      RECT 58.63 0.905 59.48 1.065 ;
      RECT 59.31 0.495 59.48 1.065 ;
      RECT 58.63 0.9 59.02 1.065 ;
      RECT 59.25 0.495 59.54 0.725 ;
      RECT 59.25 0.525 59.71 0.695 ;
      RECT 58.26 -2.685 58.55 -2.455 ;
      RECT 58.26 -2.655 58.72 -2.485 ;
      RECT 58.32 -3.765 58.485 -2.455 ;
      RECT 56.835 -3.795 57.125 -3.565 ;
      RECT 56.835 -3.765 58.485 -3.595 ;
      RECT 56.895 -4.535 57.065 -3.565 ;
      RECT 56.835 -4.535 57.125 -4.305 ;
      RECT 56.835 2.345 57.125 2.575 ;
      RECT 56.895 1.605 57.065 2.575 ;
      RECT 56.895 1.7 58.485 1.87 ;
      RECT 58.315 0.495 58.485 1.87 ;
      RECT 56.835 1.605 57.125 1.835 ;
      RECT 58.26 0.495 58.55 0.725 ;
      RECT 58.26 0.525 58.72 0.695 ;
      RECT 57.265 -3.455 57.615 -3.105 ;
      RECT 57.095 -3.395 57.615 -3.225 ;
      RECT 57.29 1.235 57.615 1.56 ;
      RECT 57.265 1.235 57.615 1.465 ;
      RECT 57.095 1.265 57.615 1.435 ;
      RECT 56.49 -3.055 56.81 -2.735 ;
      RECT 56.46 -3.055 56.81 -2.825 ;
      RECT 56.175 -3.025 56.81 -2.855 ;
      RECT 56.49 0.86 56.81 1.185 ;
      RECT 56.46 0.865 56.81 1.095 ;
      RECT 56.29 0.895 56.81 1.065 ;
      RECT 55.445 -1.925 55.77 -1.6 ;
      RECT 55.525 -2.685 55.695 -1.6 ;
      RECT 55.465 -2.685 55.755 -2.455 ;
      RECT 55.465 -2.655 55.925 -2.485 ;
      RECT 55.445 0.435 55.77 0.76 ;
      RECT 55.445 0.525 55.925 0.695 ;
      RECT 54.735 -1.765 55.06 -1.44 ;
      RECT 54.86 -3.425 55.025 -1.44 ;
      RECT 54.82 -3.425 55.145 -3.1 ;
      RECT 52.235 -1.63 52.555 -1.37 ;
      RECT 53.27 -1.615 53.56 -1.385 ;
      RECT 52.235 -1.57 53.56 -1.43 ;
      RECT 51.895 0.41 52.215 0.67 ;
      RECT 53.27 0.425 53.56 0.655 ;
      RECT 53.345 0.13 53.485 0.655 ;
      RECT 51.985 0.13 52.125 0.67 ;
      RECT 51.985 0.13 53.485 0.27 ;
      RECT 52.915 -2.65 53.235 -2.39 ;
      RECT 52.64 -2.59 53.235 -2.45 ;
      RECT 49.855 1.09 50.175 1.35 ;
      RECT 48.85 1.105 49.14 1.335 ;
      RECT 48.85 1.15 50.765 1.29 ;
      RECT 50.625 0.81 50.765 1.29 ;
      RECT 50.625 0.81 52.635 0.95 ;
      RECT 52.495 0.425 52.635 0.95 ;
      RECT 52.42 0.425 52.71 0.655 ;
      RECT 52.235 -0.61 52.555 -0.35 ;
      RECT 50.09 -0.595 50.38 -0.365 ;
      RECT 50.09 -0.55 52.555 -0.41 ;
      RECT 51.555 -1.63 51.875 -1.37 ;
      RECT 49.19 -1.615 49.48 -1.385 ;
      RECT 49.19 -1.57 51.875 -1.43 ;
      RECT 51.215 1.09 51.535 1.35 ;
      RECT 51.215 1.15 51.81 1.29 ;
      RECT 51.215 -2.31 51.535 -2.05 ;
      RECT 50.94 -2.25 51.535 -2.11 ;
      RECT 50.535 -2.65 50.855 -2.39 ;
      RECT 50.26 -2.59 50.855 -2.45 ;
      RECT 50.195 -1.97 50.515 -1.71 ;
      RECT 47.32 -1.955 47.61 -1.725 ;
      RECT 47.32 -1.91 50.515 -1.77 ;
      RECT 49.775 -2.63 49.915 -1.77 ;
      RECT 49.7 -2.63 49.99 -2.4 ;
      RECT 49.855 -3.16 50.175 -2.9 ;
      RECT 49.855 -3.145 50.36 -2.915 ;
      RECT 49.765 -3.1 50.36 -2.96 ;
      RECT 49.175 0.41 49.495 0.67 ;
      RECT 46.81 0.425 47.1 0.655 ;
      RECT 46.81 0.47 49.495 0.61 ;
      RECT 49.19 -2.63 49.48 -2.4 ;
      RECT 48.585 -2.585 49.48 -2.445 ;
      RECT 48.585 -2.99 48.725 -2.445 ;
      RECT 48.495 -2.99 48.815 -2.73 ;
      RECT 47.815 -2.65 48.135 -2.39 ;
      RECT 47.54 -2.59 48.135 -2.45 ;
      RECT 47.815 -0.61 48.135 -0.35 ;
      RECT 47.54 -0.55 48.135 -0.41 ;
      RECT 45.445 -3.055 45.735 -2.825 ;
      RECT 45.505 -4.535 45.675 -2.825 ;
      RECT 45.47 -4.325 45.82 -3.975 ;
      RECT 45.445 -4.535 45.735 -4.305 ;
      RECT 45.445 2.345 45.735 2.575 ;
      RECT 45.505 0.865 45.675 2.575 ;
      RECT 45.445 0.865 45.735 1.095 ;
      RECT 45.035 -2.685 45.365 -2.455 ;
      RECT 45.035 -2.655 45.535 -2.485 ;
      RECT 45.035 -3.025 45.225 -2.455 ;
      RECT 44.455 -3.055 44.745 -2.825 ;
      RECT 44.455 -3.025 45.225 -2.855 ;
      RECT 44.515 -4.535 44.685 -2.825 ;
      RECT 44.455 -4.535 44.745 -4.305 ;
      RECT 44.455 2.345 44.745 2.575 ;
      RECT 44.515 0.865 44.685 2.575 ;
      RECT 44.455 0.865 44.745 1.095 ;
      RECT 44.455 0.905 45.305 1.065 ;
      RECT 45.135 0.495 45.305 1.065 ;
      RECT 44.455 0.9 44.845 1.065 ;
      RECT 45.075 0.495 45.365 0.725 ;
      RECT 45.075 0.525 45.535 0.695 ;
      RECT 44.085 -2.685 44.375 -2.455 ;
      RECT 44.085 -2.655 44.545 -2.485 ;
      RECT 44.145 -3.765 44.31 -2.455 ;
      RECT 42.66 -3.795 42.95 -3.565 ;
      RECT 42.66 -3.765 44.31 -3.595 ;
      RECT 42.72 -4.535 42.89 -3.565 ;
      RECT 42.66 -4.535 42.95 -4.305 ;
      RECT 42.66 2.345 42.95 2.575 ;
      RECT 42.72 1.605 42.89 2.575 ;
      RECT 42.72 1.7 44.31 1.87 ;
      RECT 44.14 0.495 44.31 1.87 ;
      RECT 42.66 1.605 42.95 1.835 ;
      RECT 44.085 0.495 44.375 0.725 ;
      RECT 44.085 0.525 44.545 0.695 ;
      RECT 43.09 -3.455 43.44 -3.105 ;
      RECT 42.92 -3.395 43.44 -3.225 ;
      RECT 43.115 1.235 43.44 1.56 ;
      RECT 43.09 1.235 43.44 1.465 ;
      RECT 42.92 1.265 43.44 1.435 ;
      RECT 42.315 -3.055 42.635 -2.735 ;
      RECT 42.285 -3.055 42.635 -2.825 ;
      RECT 42 -3.025 42.635 -2.855 ;
      RECT 42.315 0.86 42.635 1.185 ;
      RECT 42.285 0.865 42.635 1.095 ;
      RECT 42.115 0.895 42.635 1.065 ;
      RECT 41.27 -1.925 41.595 -1.6 ;
      RECT 41.35 -2.685 41.52 -1.6 ;
      RECT 41.29 -2.685 41.58 -2.455 ;
      RECT 41.29 -2.655 41.75 -2.485 ;
      RECT 41.27 0.435 41.595 0.76 ;
      RECT 41.27 0.525 41.75 0.695 ;
      RECT 40.56 -1.765 40.885 -1.44 ;
      RECT 40.685 -3.425 40.85 -1.44 ;
      RECT 40.645 -3.425 40.97 -3.1 ;
      RECT 38.06 -1.63 38.38 -1.37 ;
      RECT 39.095 -1.615 39.385 -1.385 ;
      RECT 38.06 -1.57 39.385 -1.43 ;
      RECT 37.72 0.41 38.04 0.67 ;
      RECT 39.095 0.425 39.385 0.655 ;
      RECT 39.17 0.13 39.31 0.655 ;
      RECT 37.81 0.13 37.95 0.67 ;
      RECT 37.81 0.13 39.31 0.27 ;
      RECT 38.74 -2.65 39.06 -2.39 ;
      RECT 38.465 -2.59 39.06 -2.45 ;
      RECT 35.68 1.09 36 1.35 ;
      RECT 34.675 1.105 34.965 1.335 ;
      RECT 34.675 1.15 36.59 1.29 ;
      RECT 36.45 0.81 36.59 1.29 ;
      RECT 36.45 0.81 38.46 0.95 ;
      RECT 38.32 0.425 38.46 0.95 ;
      RECT 38.245 0.425 38.535 0.655 ;
      RECT 38.06 -0.61 38.38 -0.35 ;
      RECT 35.915 -0.595 36.205 -0.365 ;
      RECT 35.915 -0.55 38.38 -0.41 ;
      RECT 37.38 -1.63 37.7 -1.37 ;
      RECT 35.015 -1.615 35.305 -1.385 ;
      RECT 35.015 -1.57 37.7 -1.43 ;
      RECT 37.04 1.09 37.36 1.35 ;
      RECT 37.04 1.15 37.635 1.29 ;
      RECT 37.04 -2.31 37.36 -2.05 ;
      RECT 36.765 -2.25 37.36 -2.11 ;
      RECT 36.36 -2.65 36.68 -2.39 ;
      RECT 36.085 -2.59 36.68 -2.45 ;
      RECT 36.02 -1.97 36.34 -1.71 ;
      RECT 33.145 -1.955 33.435 -1.725 ;
      RECT 33.145 -1.91 36.34 -1.77 ;
      RECT 35.6 -2.63 35.74 -1.77 ;
      RECT 35.525 -2.63 35.815 -2.4 ;
      RECT 35.68 -3.16 36 -2.9 ;
      RECT 35.68 -3.145 36.185 -2.915 ;
      RECT 35.59 -3.1 36.185 -2.96 ;
      RECT 35 0.41 35.32 0.67 ;
      RECT 32.635 0.425 32.925 0.655 ;
      RECT 32.635 0.47 35.32 0.61 ;
      RECT 35.015 -2.63 35.305 -2.4 ;
      RECT 34.41 -2.585 35.305 -2.445 ;
      RECT 34.41 -2.99 34.55 -2.445 ;
      RECT 34.32 -2.99 34.64 -2.73 ;
      RECT 33.64 -2.65 33.96 -2.39 ;
      RECT 33.365 -2.59 33.96 -2.45 ;
      RECT 33.64 -0.61 33.96 -0.35 ;
      RECT 33.365 -0.55 33.96 -0.41 ;
      RECT 31.275 -3.065 31.565 -2.835 ;
      RECT 31.335 -4.545 31.505 -2.835 ;
      RECT 31.31 -4.33 31.66 -3.98 ;
      RECT 31.275 -4.545 31.565 -4.315 ;
      RECT 31.275 2.335 31.565 2.565 ;
      RECT 31.335 0.855 31.505 2.565 ;
      RECT 31.275 0.855 31.565 1.085 ;
      RECT 30.865 -2.695 31.195 -2.465 ;
      RECT 30.865 -2.665 31.365 -2.495 ;
      RECT 30.865 -3.035 31.055 -2.465 ;
      RECT 30.285 -3.065 30.575 -2.835 ;
      RECT 30.285 -3.035 31.055 -2.865 ;
      RECT 30.345 -4.545 30.515 -2.835 ;
      RECT 30.285 -4.545 30.575 -4.315 ;
      RECT 30.285 2.335 30.575 2.565 ;
      RECT 30.345 0.855 30.515 2.565 ;
      RECT 30.285 0.855 30.575 1.085 ;
      RECT 30.285 0.895 31.135 1.055 ;
      RECT 30.965 0.485 31.135 1.055 ;
      RECT 30.285 0.89 30.675 1.055 ;
      RECT 30.905 0.485 31.195 0.715 ;
      RECT 30.905 0.515 31.365 0.685 ;
      RECT 29.915 -2.695 30.205 -2.465 ;
      RECT 29.915 -2.665 30.375 -2.495 ;
      RECT 29.975 -3.775 30.14 -2.465 ;
      RECT 28.49 -3.805 28.78 -3.575 ;
      RECT 28.49 -3.775 30.14 -3.605 ;
      RECT 28.55 -4.545 28.72 -3.575 ;
      RECT 28.49 -4.545 28.78 -4.315 ;
      RECT 28.49 2.335 28.78 2.565 ;
      RECT 28.55 1.595 28.72 2.565 ;
      RECT 28.55 1.69 30.14 1.86 ;
      RECT 29.97 0.485 30.14 1.86 ;
      RECT 28.49 1.595 28.78 1.825 ;
      RECT 29.915 0.485 30.205 0.715 ;
      RECT 29.915 0.515 30.375 0.685 ;
      RECT 28.92 -3.465 29.27 -3.115 ;
      RECT 28.75 -3.405 29.27 -3.235 ;
      RECT 28.945 1.225 29.27 1.55 ;
      RECT 28.92 1.225 29.27 1.455 ;
      RECT 28.75 1.255 29.27 1.425 ;
      RECT 28.145 -3.065 28.465 -2.745 ;
      RECT 28.115 -3.065 28.465 -2.835 ;
      RECT 27.83 -3.035 28.465 -2.865 ;
      RECT 28.145 0.85 28.465 1.175 ;
      RECT 28.115 0.855 28.465 1.085 ;
      RECT 27.945 0.885 28.465 1.055 ;
      RECT 27.1 -1.935 27.425 -1.61 ;
      RECT 27.18 -2.695 27.35 -1.61 ;
      RECT 27.12 -2.695 27.41 -2.465 ;
      RECT 27.12 -2.665 27.58 -2.495 ;
      RECT 27.1 0.425 27.425 0.75 ;
      RECT 27.1 0.515 27.58 0.685 ;
      RECT 26.39 -1.775 26.715 -1.45 ;
      RECT 26.515 -3.435 26.68 -1.45 ;
      RECT 26.475 -3.435 26.8 -3.11 ;
      RECT 23.89 -1.64 24.21 -1.38 ;
      RECT 24.925 -1.625 25.215 -1.395 ;
      RECT 23.89 -1.58 25.215 -1.44 ;
      RECT 23.55 0.4 23.87 0.66 ;
      RECT 24.925 0.415 25.215 0.645 ;
      RECT 25 0.12 25.14 0.645 ;
      RECT 23.64 0.12 23.78 0.66 ;
      RECT 23.64 0.12 25.14 0.26 ;
      RECT 24.57 -2.66 24.89 -2.4 ;
      RECT 24.295 -2.6 24.89 -2.46 ;
      RECT 21.51 1.08 21.83 1.34 ;
      RECT 20.505 1.095 20.795 1.325 ;
      RECT 20.505 1.14 22.42 1.28 ;
      RECT 22.28 0.8 22.42 1.28 ;
      RECT 22.28 0.8 24.29 0.94 ;
      RECT 24.15 0.415 24.29 0.94 ;
      RECT 24.075 0.415 24.365 0.645 ;
      RECT 23.89 -0.62 24.21 -0.36 ;
      RECT 21.745 -0.605 22.035 -0.375 ;
      RECT 21.745 -0.56 24.21 -0.42 ;
      RECT 23.21 -1.64 23.53 -1.38 ;
      RECT 20.845 -1.625 21.135 -1.395 ;
      RECT 20.845 -1.58 23.53 -1.44 ;
      RECT 22.87 1.08 23.19 1.34 ;
      RECT 22.87 1.14 23.465 1.28 ;
      RECT 22.87 -2.32 23.19 -2.06 ;
      RECT 22.595 -2.26 23.19 -2.12 ;
      RECT 22.19 -2.66 22.51 -2.4 ;
      RECT 21.915 -2.6 22.51 -2.46 ;
      RECT 21.85 -1.98 22.17 -1.72 ;
      RECT 18.975 -1.965 19.265 -1.735 ;
      RECT 18.975 -1.92 22.17 -1.78 ;
      RECT 21.43 -2.64 21.57 -1.78 ;
      RECT 21.355 -2.64 21.645 -2.41 ;
      RECT 21.51 -3.17 21.83 -2.91 ;
      RECT 21.51 -3.155 22.015 -2.925 ;
      RECT 21.42 -3.11 22.015 -2.97 ;
      RECT 20.83 0.4 21.15 0.66 ;
      RECT 18.465 0.415 18.755 0.645 ;
      RECT 18.465 0.46 21.15 0.6 ;
      RECT 20.845 -2.64 21.135 -2.41 ;
      RECT 20.24 -2.595 21.135 -2.455 ;
      RECT 20.24 -3 20.38 -2.455 ;
      RECT 20.15 -3 20.47 -2.74 ;
      RECT 19.47 -2.66 19.79 -2.4 ;
      RECT 19.195 -2.6 19.79 -2.46 ;
      RECT 19.47 -0.62 19.79 -0.36 ;
      RECT 19.195 -0.56 19.79 -0.42 ;
      RECT 17.11 -3.065 17.4 -2.835 ;
      RECT 17.17 -4.545 17.34 -2.835 ;
      RECT 17.14 -4.33 17.49 -3.98 ;
      RECT 17.11 -4.545 17.4 -4.315 ;
      RECT 17.11 2.335 17.4 2.565 ;
      RECT 17.17 0.855 17.34 2.565 ;
      RECT 17.11 0.855 17.4 1.085 ;
      RECT 16.7 -2.695 17.03 -2.465 ;
      RECT 16.7 -2.665 17.2 -2.495 ;
      RECT 16.7 -3.035 16.89 -2.465 ;
      RECT 16.12 -3.065 16.41 -2.835 ;
      RECT 16.12 -3.035 16.89 -2.865 ;
      RECT 16.18 -4.545 16.35 -2.835 ;
      RECT 16.12 -4.545 16.41 -4.315 ;
      RECT 16.12 2.335 16.41 2.565 ;
      RECT 16.18 0.855 16.35 2.565 ;
      RECT 16.12 0.855 16.41 1.085 ;
      RECT 16.12 0.895 16.97 1.055 ;
      RECT 16.8 0.485 16.97 1.055 ;
      RECT 16.12 0.89 16.51 1.055 ;
      RECT 16.74 0.485 17.03 0.715 ;
      RECT 16.74 0.515 17.2 0.685 ;
      RECT 15.75 -2.695 16.04 -2.465 ;
      RECT 15.75 -2.665 16.21 -2.495 ;
      RECT 15.81 -3.775 15.975 -2.465 ;
      RECT 14.325 -3.805 14.615 -3.575 ;
      RECT 14.325 -3.775 15.975 -3.605 ;
      RECT 14.385 -4.545 14.555 -3.575 ;
      RECT 14.325 -4.545 14.615 -4.315 ;
      RECT 14.325 2.335 14.615 2.565 ;
      RECT 14.385 1.595 14.555 2.565 ;
      RECT 14.385 1.69 15.975 1.86 ;
      RECT 15.805 0.485 15.975 1.86 ;
      RECT 14.325 1.595 14.615 1.825 ;
      RECT 15.75 0.485 16.04 0.715 ;
      RECT 15.75 0.515 16.21 0.685 ;
      RECT 14.755 -3.465 15.105 -3.115 ;
      RECT 14.585 -3.405 15.105 -3.235 ;
      RECT 14.78 1.225 15.105 1.55 ;
      RECT 14.755 1.225 15.105 1.455 ;
      RECT 14.585 1.255 15.105 1.425 ;
      RECT 13.98 -3.065 14.3 -2.745 ;
      RECT 13.95 -3.065 14.3 -2.835 ;
      RECT 13.665 -3.035 14.3 -2.865 ;
      RECT 13.98 0.85 14.3 1.175 ;
      RECT 13.95 0.855 14.3 1.085 ;
      RECT 13.78 0.885 14.3 1.055 ;
      RECT 12.935 -1.935 13.26 -1.61 ;
      RECT 13.015 -2.695 13.185 -1.61 ;
      RECT 12.955 -2.695 13.245 -2.465 ;
      RECT 12.955 -2.665 13.415 -2.495 ;
      RECT 12.935 0.425 13.26 0.75 ;
      RECT 12.935 0.515 13.415 0.685 ;
      RECT 12.225 -1.775 12.55 -1.45 ;
      RECT 12.35 -3.435 12.515 -1.45 ;
      RECT 12.31 -3.435 12.635 -3.11 ;
      RECT 9.725 -1.64 10.045 -1.38 ;
      RECT 10.76 -1.625 11.05 -1.395 ;
      RECT 9.725 -1.58 11.05 -1.44 ;
      RECT 9.385 0.4 9.705 0.66 ;
      RECT 10.76 0.415 11.05 0.645 ;
      RECT 10.835 0.12 10.975 0.645 ;
      RECT 9.475 0.12 9.615 0.66 ;
      RECT 9.475 0.12 10.975 0.26 ;
      RECT 10.405 -2.66 10.725 -2.4 ;
      RECT 10.13 -2.6 10.725 -2.46 ;
      RECT 7.345 1.08 7.665 1.34 ;
      RECT 6.34 1.095 6.63 1.325 ;
      RECT 6.34 1.14 8.255 1.28 ;
      RECT 8.115 0.8 8.255 1.28 ;
      RECT 8.115 0.8 10.125 0.94 ;
      RECT 9.985 0.415 10.125 0.94 ;
      RECT 9.91 0.415 10.2 0.645 ;
      RECT 9.725 -0.62 10.045 -0.36 ;
      RECT 7.58 -0.605 7.87 -0.375 ;
      RECT 7.58 -0.56 10.045 -0.42 ;
      RECT 9.045 -1.64 9.365 -1.38 ;
      RECT 6.68 -1.625 6.97 -1.395 ;
      RECT 6.68 -1.58 9.365 -1.44 ;
      RECT 8.705 1.08 9.025 1.34 ;
      RECT 8.705 1.14 9.3 1.28 ;
      RECT 8.705 -2.32 9.025 -2.06 ;
      RECT 8.43 -2.26 9.025 -2.12 ;
      RECT 8.025 -2.66 8.345 -2.4 ;
      RECT 7.75 -2.6 8.345 -2.46 ;
      RECT 7.685 -1.98 8.005 -1.72 ;
      RECT 4.81 -1.965 5.1 -1.735 ;
      RECT 4.81 -1.92 8.005 -1.78 ;
      RECT 7.265 -2.64 7.405 -1.78 ;
      RECT 7.19 -2.64 7.48 -2.41 ;
      RECT 7.345 -3.17 7.665 -2.91 ;
      RECT 7.345 -3.155 7.85 -2.925 ;
      RECT 7.255 -3.11 7.85 -2.97 ;
      RECT 6.665 0.4 6.985 0.66 ;
      RECT 4.3 0.415 4.59 0.645 ;
      RECT 4.3 0.46 6.985 0.6 ;
      RECT 6.68 -2.64 6.97 -2.41 ;
      RECT 6.075 -2.595 6.97 -2.455 ;
      RECT 6.075 -3 6.215 -2.455 ;
      RECT 5.985 -3 6.305 -2.74 ;
      RECT 5.305 -2.66 5.625 -2.4 ;
      RECT 5.03 -2.6 5.625 -2.46 ;
      RECT 5.305 -0.62 5.625 -0.36 ;
      RECT 5.03 -0.56 5.625 -0.42 ;
      RECT 66.765 1.09 67.41 1.35 ;
      RECT 64.715 0.41 65.36 0.67 ;
      RECT 52.59 1.09 53.235 1.35 ;
      RECT 50.54 0.41 51.185 0.67 ;
      RECT 38.415 1.09 39.06 1.35 ;
      RECT 36.365 0.41 37.01 0.67 ;
      RECT 24.245 1.08 24.89 1.34 ;
      RECT 22.195 0.4 22.84 0.66 ;
      RECT 10.08 1.08 10.725 1.34 ;
      RECT 8.03 0.4 8.675 0.66 ;
    LAYER mcon ;
      RECT 73.855 -4.505 74.025 -4.335 ;
      RECT 73.855 -3.025 74.025 -2.855 ;
      RECT 73.855 0.895 74.025 1.065 ;
      RECT 73.855 2.375 74.025 2.545 ;
      RECT 73.505 -5.315 73.675 -5.145 ;
      RECT 73.505 -1.255 73.675 -1.085 ;
      RECT 73.505 -0.875 73.675 -0.705 ;
      RECT 73.505 3.185 73.675 3.355 ;
      RECT 73.485 -2.655 73.655 -2.485 ;
      RECT 73.485 0.525 73.655 0.695 ;
      RECT 72.865 -4.505 73.035 -4.335 ;
      RECT 72.865 -3.025 73.035 -2.855 ;
      RECT 72.865 0.895 73.035 1.065 ;
      RECT 72.865 2.375 73.035 2.545 ;
      RECT 72.515 -5.315 72.685 -5.145 ;
      RECT 72.515 -1.255 72.685 -1.085 ;
      RECT 72.515 -0.875 72.685 -0.705 ;
      RECT 72.515 3.185 72.685 3.355 ;
      RECT 72.495 -2.655 72.665 -2.485 ;
      RECT 72.495 0.525 72.665 0.695 ;
      RECT 71.81 -5.315 71.98 -5.145 ;
      RECT 71.81 -1.255 71.98 -1.085 ;
      RECT 71.81 -0.875 71.98 -0.705 ;
      RECT 71.81 3.185 71.98 3.355 ;
      RECT 71.5 -3.395 71.67 -3.225 ;
      RECT 71.5 1.265 71.67 1.435 ;
      RECT 71.13 -5.315 71.3 -5.145 ;
      RECT 71.13 3.185 71.3 3.355 ;
      RECT 71.07 -4.505 71.24 -4.335 ;
      RECT 71.07 -3.765 71.24 -3.595 ;
      RECT 71.07 1.635 71.24 1.805 ;
      RECT 71.07 2.375 71.24 2.545 ;
      RECT 70.695 -3.025 70.865 -2.855 ;
      RECT 70.695 0.895 70.865 1.065 ;
      RECT 70.45 -5.315 70.62 -5.145 ;
      RECT 70.45 3.185 70.62 3.355 ;
      RECT 69.77 -5.315 69.94 -5.145 ;
      RECT 69.77 3.185 69.94 3.355 ;
      RECT 69.7 -2.655 69.87 -2.485 ;
      RECT 69.7 0.525 69.87 0.695 ;
      RECT 68.005 -3.795 68.175 -3.625 ;
      RECT 68.005 -1.075 68.175 -0.905 ;
      RECT 68.005 1.645 68.175 1.815 ;
      RECT 67.545 -3.795 67.715 -3.625 ;
      RECT 67.545 -1.075 67.715 -0.905 ;
      RECT 67.545 1.645 67.715 1.815 ;
      RECT 67.505 -1.585 67.675 -1.415 ;
      RECT 67.505 0.455 67.675 0.625 ;
      RECT 67.165 -2.605 67.335 -2.435 ;
      RECT 67.085 -3.795 67.255 -3.625 ;
      RECT 67.085 -1.075 67.255 -0.905 ;
      RECT 67.085 1.645 67.255 1.815 ;
      RECT 66.825 1.135 66.995 1.305 ;
      RECT 66.655 0.455 66.825 0.625 ;
      RECT 66.625 -3.795 66.795 -3.625 ;
      RECT 66.625 -1.075 66.795 -0.905 ;
      RECT 66.625 1.645 66.795 1.815 ;
      RECT 66.165 -3.795 66.335 -3.625 ;
      RECT 66.165 -1.075 66.335 -0.905 ;
      RECT 66.165 1.645 66.335 1.815 ;
      RECT 66.145 0.455 66.315 0.625 ;
      RECT 65.705 -3.795 65.875 -3.625 ;
      RECT 65.705 -1.075 65.875 -0.905 ;
      RECT 65.705 1.645 65.875 1.815 ;
      RECT 65.465 -2.265 65.635 -2.095 ;
      RECT 65.465 1.135 65.635 1.305 ;
      RECT 65.245 -3.795 65.415 -3.625 ;
      RECT 65.245 -1.075 65.415 -0.905 ;
      RECT 65.245 1.645 65.415 1.815 ;
      RECT 64.785 -3.795 64.955 -3.625 ;
      RECT 64.785 -2.605 64.955 -2.435 ;
      RECT 64.785 -1.075 64.955 -0.905 ;
      RECT 64.785 1.645 64.955 1.815 ;
      RECT 64.775 0.455 64.945 0.625 ;
      RECT 64.325 -3.795 64.495 -3.625 ;
      RECT 64.325 -1.075 64.495 -0.905 ;
      RECT 64.325 -0.565 64.495 -0.395 ;
      RECT 64.325 1.645 64.495 1.815 ;
      RECT 64.305 -3.115 64.475 -2.945 ;
      RECT 63.935 -2.6 64.105 -2.43 ;
      RECT 63.865 -3.795 64.035 -3.625 ;
      RECT 63.865 -1.075 64.035 -0.905 ;
      RECT 63.865 1.645 64.035 1.815 ;
      RECT 63.425 -2.6 63.595 -2.43 ;
      RECT 63.425 -1.585 63.595 -1.415 ;
      RECT 63.425 0.455 63.595 0.625 ;
      RECT 63.405 -3.795 63.575 -3.625 ;
      RECT 63.405 -1.075 63.575 -0.905 ;
      RECT 63.405 1.645 63.575 1.815 ;
      RECT 63.085 1.135 63.255 1.305 ;
      RECT 62.945 -3.795 63.115 -3.625 ;
      RECT 62.945 -1.075 63.115 -0.905 ;
      RECT 62.945 1.645 63.115 1.815 ;
      RECT 62.485 -3.795 62.655 -3.625 ;
      RECT 62.485 -1.075 62.655 -0.905 ;
      RECT 62.485 1.645 62.655 1.815 ;
      RECT 62.065 -2.605 62.235 -2.435 ;
      RECT 62.065 -0.565 62.235 -0.395 ;
      RECT 62.025 -3.795 62.195 -3.625 ;
      RECT 62.025 -1.075 62.195 -0.905 ;
      RECT 62.025 1.645 62.195 1.815 ;
      RECT 61.565 -3.795 61.735 -3.625 ;
      RECT 61.565 -1.075 61.735 -0.905 ;
      RECT 61.565 1.645 61.735 1.815 ;
      RECT 61.555 -1.925 61.725 -1.755 ;
      RECT 61.105 -3.795 61.275 -3.625 ;
      RECT 61.105 -1.075 61.275 -0.905 ;
      RECT 61.105 1.645 61.275 1.815 ;
      RECT 61.045 0.455 61.215 0.625 ;
      RECT 59.68 -4.505 59.85 -4.335 ;
      RECT 59.68 -3.025 59.85 -2.855 ;
      RECT 59.68 0.895 59.85 1.065 ;
      RECT 59.68 2.375 59.85 2.545 ;
      RECT 59.33 -5.315 59.5 -5.145 ;
      RECT 59.33 -1.255 59.5 -1.085 ;
      RECT 59.33 -0.875 59.5 -0.705 ;
      RECT 59.33 3.185 59.5 3.355 ;
      RECT 59.31 -2.655 59.48 -2.485 ;
      RECT 59.31 0.525 59.48 0.695 ;
      RECT 58.69 -4.505 58.86 -4.335 ;
      RECT 58.69 -3.025 58.86 -2.855 ;
      RECT 58.69 0.895 58.86 1.065 ;
      RECT 58.69 2.375 58.86 2.545 ;
      RECT 58.34 -5.315 58.51 -5.145 ;
      RECT 58.34 -1.255 58.51 -1.085 ;
      RECT 58.34 -0.875 58.51 -0.705 ;
      RECT 58.34 3.185 58.51 3.355 ;
      RECT 58.32 -2.655 58.49 -2.485 ;
      RECT 58.32 0.525 58.49 0.695 ;
      RECT 57.635 -5.315 57.805 -5.145 ;
      RECT 57.635 -1.255 57.805 -1.085 ;
      RECT 57.635 -0.875 57.805 -0.705 ;
      RECT 57.635 3.185 57.805 3.355 ;
      RECT 57.325 -3.395 57.495 -3.225 ;
      RECT 57.325 1.265 57.495 1.435 ;
      RECT 56.955 -5.315 57.125 -5.145 ;
      RECT 56.955 3.185 57.125 3.355 ;
      RECT 56.895 -4.505 57.065 -4.335 ;
      RECT 56.895 -3.765 57.065 -3.595 ;
      RECT 56.895 1.635 57.065 1.805 ;
      RECT 56.895 2.375 57.065 2.545 ;
      RECT 56.52 -3.025 56.69 -2.855 ;
      RECT 56.52 0.895 56.69 1.065 ;
      RECT 56.275 -5.315 56.445 -5.145 ;
      RECT 56.275 3.185 56.445 3.355 ;
      RECT 55.595 -5.315 55.765 -5.145 ;
      RECT 55.595 3.185 55.765 3.355 ;
      RECT 55.525 -2.655 55.695 -2.485 ;
      RECT 55.525 0.525 55.695 0.695 ;
      RECT 53.83 -3.795 54 -3.625 ;
      RECT 53.83 -1.075 54 -0.905 ;
      RECT 53.83 1.645 54 1.815 ;
      RECT 53.37 -3.795 53.54 -3.625 ;
      RECT 53.37 -1.075 53.54 -0.905 ;
      RECT 53.37 1.645 53.54 1.815 ;
      RECT 53.33 -1.585 53.5 -1.415 ;
      RECT 53.33 0.455 53.5 0.625 ;
      RECT 52.99 -2.605 53.16 -2.435 ;
      RECT 52.91 -3.795 53.08 -3.625 ;
      RECT 52.91 -1.075 53.08 -0.905 ;
      RECT 52.91 1.645 53.08 1.815 ;
      RECT 52.65 1.135 52.82 1.305 ;
      RECT 52.48 0.455 52.65 0.625 ;
      RECT 52.45 -3.795 52.62 -3.625 ;
      RECT 52.45 -1.075 52.62 -0.905 ;
      RECT 52.45 1.645 52.62 1.815 ;
      RECT 51.99 -3.795 52.16 -3.625 ;
      RECT 51.99 -1.075 52.16 -0.905 ;
      RECT 51.99 1.645 52.16 1.815 ;
      RECT 51.97 0.455 52.14 0.625 ;
      RECT 51.53 -3.795 51.7 -3.625 ;
      RECT 51.53 -1.075 51.7 -0.905 ;
      RECT 51.53 1.645 51.7 1.815 ;
      RECT 51.29 -2.265 51.46 -2.095 ;
      RECT 51.29 1.135 51.46 1.305 ;
      RECT 51.07 -3.795 51.24 -3.625 ;
      RECT 51.07 -1.075 51.24 -0.905 ;
      RECT 51.07 1.645 51.24 1.815 ;
      RECT 50.61 -3.795 50.78 -3.625 ;
      RECT 50.61 -2.605 50.78 -2.435 ;
      RECT 50.61 -1.075 50.78 -0.905 ;
      RECT 50.61 1.645 50.78 1.815 ;
      RECT 50.6 0.455 50.77 0.625 ;
      RECT 50.15 -3.795 50.32 -3.625 ;
      RECT 50.15 -1.075 50.32 -0.905 ;
      RECT 50.15 -0.565 50.32 -0.395 ;
      RECT 50.15 1.645 50.32 1.815 ;
      RECT 50.13 -3.115 50.3 -2.945 ;
      RECT 49.76 -2.6 49.93 -2.43 ;
      RECT 49.69 -3.795 49.86 -3.625 ;
      RECT 49.69 -1.075 49.86 -0.905 ;
      RECT 49.69 1.645 49.86 1.815 ;
      RECT 49.25 -2.6 49.42 -2.43 ;
      RECT 49.25 -1.585 49.42 -1.415 ;
      RECT 49.25 0.455 49.42 0.625 ;
      RECT 49.23 -3.795 49.4 -3.625 ;
      RECT 49.23 -1.075 49.4 -0.905 ;
      RECT 49.23 1.645 49.4 1.815 ;
      RECT 48.91 1.135 49.08 1.305 ;
      RECT 48.77 -3.795 48.94 -3.625 ;
      RECT 48.77 -1.075 48.94 -0.905 ;
      RECT 48.77 1.645 48.94 1.815 ;
      RECT 48.31 -3.795 48.48 -3.625 ;
      RECT 48.31 -1.075 48.48 -0.905 ;
      RECT 48.31 1.645 48.48 1.815 ;
      RECT 47.89 -2.605 48.06 -2.435 ;
      RECT 47.89 -0.565 48.06 -0.395 ;
      RECT 47.85 -3.795 48.02 -3.625 ;
      RECT 47.85 -1.075 48.02 -0.905 ;
      RECT 47.85 1.645 48.02 1.815 ;
      RECT 47.39 -3.795 47.56 -3.625 ;
      RECT 47.39 -1.075 47.56 -0.905 ;
      RECT 47.39 1.645 47.56 1.815 ;
      RECT 47.38 -1.925 47.55 -1.755 ;
      RECT 46.93 -3.795 47.1 -3.625 ;
      RECT 46.93 -1.075 47.1 -0.905 ;
      RECT 46.93 1.645 47.1 1.815 ;
      RECT 46.87 0.455 47.04 0.625 ;
      RECT 45.505 -4.505 45.675 -4.335 ;
      RECT 45.505 -3.025 45.675 -2.855 ;
      RECT 45.505 0.895 45.675 1.065 ;
      RECT 45.505 2.375 45.675 2.545 ;
      RECT 45.155 -5.315 45.325 -5.145 ;
      RECT 45.155 -1.255 45.325 -1.085 ;
      RECT 45.155 -0.875 45.325 -0.705 ;
      RECT 45.155 3.185 45.325 3.355 ;
      RECT 45.135 -2.655 45.305 -2.485 ;
      RECT 45.135 0.525 45.305 0.695 ;
      RECT 44.515 -4.505 44.685 -4.335 ;
      RECT 44.515 -3.025 44.685 -2.855 ;
      RECT 44.515 0.895 44.685 1.065 ;
      RECT 44.515 2.375 44.685 2.545 ;
      RECT 44.165 -5.315 44.335 -5.145 ;
      RECT 44.165 -1.255 44.335 -1.085 ;
      RECT 44.165 -0.875 44.335 -0.705 ;
      RECT 44.165 3.185 44.335 3.355 ;
      RECT 44.145 -2.655 44.315 -2.485 ;
      RECT 44.145 0.525 44.315 0.695 ;
      RECT 43.46 -5.315 43.63 -5.145 ;
      RECT 43.46 -1.255 43.63 -1.085 ;
      RECT 43.46 -0.875 43.63 -0.705 ;
      RECT 43.46 3.185 43.63 3.355 ;
      RECT 43.15 -3.395 43.32 -3.225 ;
      RECT 43.15 1.265 43.32 1.435 ;
      RECT 42.78 -5.315 42.95 -5.145 ;
      RECT 42.78 3.185 42.95 3.355 ;
      RECT 42.72 -4.505 42.89 -4.335 ;
      RECT 42.72 -3.765 42.89 -3.595 ;
      RECT 42.72 1.635 42.89 1.805 ;
      RECT 42.72 2.375 42.89 2.545 ;
      RECT 42.345 -3.025 42.515 -2.855 ;
      RECT 42.345 0.895 42.515 1.065 ;
      RECT 42.1 -5.315 42.27 -5.145 ;
      RECT 42.1 3.185 42.27 3.355 ;
      RECT 41.42 -5.315 41.59 -5.145 ;
      RECT 41.42 3.185 41.59 3.355 ;
      RECT 41.35 -2.655 41.52 -2.485 ;
      RECT 41.35 0.525 41.52 0.695 ;
      RECT 39.655 -3.795 39.825 -3.625 ;
      RECT 39.655 -1.075 39.825 -0.905 ;
      RECT 39.655 1.645 39.825 1.815 ;
      RECT 39.195 -3.795 39.365 -3.625 ;
      RECT 39.195 -1.075 39.365 -0.905 ;
      RECT 39.195 1.645 39.365 1.815 ;
      RECT 39.155 -1.585 39.325 -1.415 ;
      RECT 39.155 0.455 39.325 0.625 ;
      RECT 38.815 -2.605 38.985 -2.435 ;
      RECT 38.735 -3.795 38.905 -3.625 ;
      RECT 38.735 -1.075 38.905 -0.905 ;
      RECT 38.735 1.645 38.905 1.815 ;
      RECT 38.475 1.135 38.645 1.305 ;
      RECT 38.305 0.455 38.475 0.625 ;
      RECT 38.275 -3.795 38.445 -3.625 ;
      RECT 38.275 -1.075 38.445 -0.905 ;
      RECT 38.275 1.645 38.445 1.815 ;
      RECT 37.815 -3.795 37.985 -3.625 ;
      RECT 37.815 -1.075 37.985 -0.905 ;
      RECT 37.815 1.645 37.985 1.815 ;
      RECT 37.795 0.455 37.965 0.625 ;
      RECT 37.355 -3.795 37.525 -3.625 ;
      RECT 37.355 -1.075 37.525 -0.905 ;
      RECT 37.355 1.645 37.525 1.815 ;
      RECT 37.115 -2.265 37.285 -2.095 ;
      RECT 37.115 1.135 37.285 1.305 ;
      RECT 36.895 -3.795 37.065 -3.625 ;
      RECT 36.895 -1.075 37.065 -0.905 ;
      RECT 36.895 1.645 37.065 1.815 ;
      RECT 36.435 -3.795 36.605 -3.625 ;
      RECT 36.435 -2.605 36.605 -2.435 ;
      RECT 36.435 -1.075 36.605 -0.905 ;
      RECT 36.435 1.645 36.605 1.815 ;
      RECT 36.425 0.455 36.595 0.625 ;
      RECT 35.975 -3.795 36.145 -3.625 ;
      RECT 35.975 -1.075 36.145 -0.905 ;
      RECT 35.975 -0.565 36.145 -0.395 ;
      RECT 35.975 1.645 36.145 1.815 ;
      RECT 35.955 -3.115 36.125 -2.945 ;
      RECT 35.585 -2.6 35.755 -2.43 ;
      RECT 35.515 -3.795 35.685 -3.625 ;
      RECT 35.515 -1.075 35.685 -0.905 ;
      RECT 35.515 1.645 35.685 1.815 ;
      RECT 35.075 -2.6 35.245 -2.43 ;
      RECT 35.075 -1.585 35.245 -1.415 ;
      RECT 35.075 0.455 35.245 0.625 ;
      RECT 35.055 -3.795 35.225 -3.625 ;
      RECT 35.055 -1.075 35.225 -0.905 ;
      RECT 35.055 1.645 35.225 1.815 ;
      RECT 34.735 1.135 34.905 1.305 ;
      RECT 34.595 -3.795 34.765 -3.625 ;
      RECT 34.595 -1.075 34.765 -0.905 ;
      RECT 34.595 1.645 34.765 1.815 ;
      RECT 34.135 -3.795 34.305 -3.625 ;
      RECT 34.135 -1.075 34.305 -0.905 ;
      RECT 34.135 1.645 34.305 1.815 ;
      RECT 33.715 -2.605 33.885 -2.435 ;
      RECT 33.715 -0.565 33.885 -0.395 ;
      RECT 33.675 -3.795 33.845 -3.625 ;
      RECT 33.675 -1.075 33.845 -0.905 ;
      RECT 33.675 1.645 33.845 1.815 ;
      RECT 33.215 -3.795 33.385 -3.625 ;
      RECT 33.215 -1.075 33.385 -0.905 ;
      RECT 33.215 1.645 33.385 1.815 ;
      RECT 33.205 -1.925 33.375 -1.755 ;
      RECT 32.755 -3.795 32.925 -3.625 ;
      RECT 32.755 -1.075 32.925 -0.905 ;
      RECT 32.755 1.645 32.925 1.815 ;
      RECT 32.695 0.455 32.865 0.625 ;
      RECT 31.335 -4.515 31.505 -4.345 ;
      RECT 31.335 -3.035 31.505 -2.865 ;
      RECT 31.335 0.885 31.505 1.055 ;
      RECT 31.335 2.365 31.505 2.535 ;
      RECT 30.985 -5.325 31.155 -5.155 ;
      RECT 30.985 -1.265 31.155 -1.095 ;
      RECT 30.985 -0.885 31.155 -0.715 ;
      RECT 30.985 3.175 31.155 3.345 ;
      RECT 30.965 -2.665 31.135 -2.495 ;
      RECT 30.965 0.515 31.135 0.685 ;
      RECT 30.345 -4.515 30.515 -4.345 ;
      RECT 30.345 -3.035 30.515 -2.865 ;
      RECT 30.345 0.885 30.515 1.055 ;
      RECT 30.345 2.365 30.515 2.535 ;
      RECT 29.995 -5.325 30.165 -5.155 ;
      RECT 29.995 -1.265 30.165 -1.095 ;
      RECT 29.995 -0.885 30.165 -0.715 ;
      RECT 29.995 3.175 30.165 3.345 ;
      RECT 29.975 -2.665 30.145 -2.495 ;
      RECT 29.975 0.515 30.145 0.685 ;
      RECT 29.29 -5.325 29.46 -5.155 ;
      RECT 29.29 -1.265 29.46 -1.095 ;
      RECT 29.29 -0.885 29.46 -0.715 ;
      RECT 29.29 3.175 29.46 3.345 ;
      RECT 28.98 -3.405 29.15 -3.235 ;
      RECT 28.98 1.255 29.15 1.425 ;
      RECT 28.61 -5.325 28.78 -5.155 ;
      RECT 28.61 3.175 28.78 3.345 ;
      RECT 28.55 -4.515 28.72 -4.345 ;
      RECT 28.55 -3.775 28.72 -3.605 ;
      RECT 28.55 1.625 28.72 1.795 ;
      RECT 28.55 2.365 28.72 2.535 ;
      RECT 28.175 -3.035 28.345 -2.865 ;
      RECT 28.175 0.885 28.345 1.055 ;
      RECT 27.93 -5.325 28.1 -5.155 ;
      RECT 27.93 3.175 28.1 3.345 ;
      RECT 27.25 -5.325 27.42 -5.155 ;
      RECT 27.25 3.175 27.42 3.345 ;
      RECT 27.18 -2.665 27.35 -2.495 ;
      RECT 27.18 0.515 27.35 0.685 ;
      RECT 25.485 -3.805 25.655 -3.635 ;
      RECT 25.485 -1.085 25.655 -0.915 ;
      RECT 25.485 1.635 25.655 1.805 ;
      RECT 25.025 -3.805 25.195 -3.635 ;
      RECT 25.025 -1.085 25.195 -0.915 ;
      RECT 25.025 1.635 25.195 1.805 ;
      RECT 24.985 -1.595 25.155 -1.425 ;
      RECT 24.985 0.445 25.155 0.615 ;
      RECT 24.645 -2.615 24.815 -2.445 ;
      RECT 24.565 -3.805 24.735 -3.635 ;
      RECT 24.565 -1.085 24.735 -0.915 ;
      RECT 24.565 1.635 24.735 1.805 ;
      RECT 24.305 1.125 24.475 1.295 ;
      RECT 24.135 0.445 24.305 0.615 ;
      RECT 24.105 -3.805 24.275 -3.635 ;
      RECT 24.105 -1.085 24.275 -0.915 ;
      RECT 24.105 1.635 24.275 1.805 ;
      RECT 23.645 -3.805 23.815 -3.635 ;
      RECT 23.645 -1.085 23.815 -0.915 ;
      RECT 23.645 1.635 23.815 1.805 ;
      RECT 23.625 0.445 23.795 0.615 ;
      RECT 23.185 -3.805 23.355 -3.635 ;
      RECT 23.185 -1.085 23.355 -0.915 ;
      RECT 23.185 1.635 23.355 1.805 ;
      RECT 22.945 -2.275 23.115 -2.105 ;
      RECT 22.945 1.125 23.115 1.295 ;
      RECT 22.725 -3.805 22.895 -3.635 ;
      RECT 22.725 -1.085 22.895 -0.915 ;
      RECT 22.725 1.635 22.895 1.805 ;
      RECT 22.265 -3.805 22.435 -3.635 ;
      RECT 22.265 -2.615 22.435 -2.445 ;
      RECT 22.265 -1.085 22.435 -0.915 ;
      RECT 22.265 1.635 22.435 1.805 ;
      RECT 22.255 0.445 22.425 0.615 ;
      RECT 21.805 -3.805 21.975 -3.635 ;
      RECT 21.805 -1.085 21.975 -0.915 ;
      RECT 21.805 -0.575 21.975 -0.405 ;
      RECT 21.805 1.635 21.975 1.805 ;
      RECT 21.785 -3.125 21.955 -2.955 ;
      RECT 21.415 -2.61 21.585 -2.44 ;
      RECT 21.345 -3.805 21.515 -3.635 ;
      RECT 21.345 -1.085 21.515 -0.915 ;
      RECT 21.345 1.635 21.515 1.805 ;
      RECT 20.905 -2.61 21.075 -2.44 ;
      RECT 20.905 -1.595 21.075 -1.425 ;
      RECT 20.905 0.445 21.075 0.615 ;
      RECT 20.885 -3.805 21.055 -3.635 ;
      RECT 20.885 -1.085 21.055 -0.915 ;
      RECT 20.885 1.635 21.055 1.805 ;
      RECT 20.565 1.125 20.735 1.295 ;
      RECT 20.425 -3.805 20.595 -3.635 ;
      RECT 20.425 -1.085 20.595 -0.915 ;
      RECT 20.425 1.635 20.595 1.805 ;
      RECT 19.965 -3.805 20.135 -3.635 ;
      RECT 19.965 -1.085 20.135 -0.915 ;
      RECT 19.965 1.635 20.135 1.805 ;
      RECT 19.545 -2.615 19.715 -2.445 ;
      RECT 19.545 -0.575 19.715 -0.405 ;
      RECT 19.505 -3.805 19.675 -3.635 ;
      RECT 19.505 -1.085 19.675 -0.915 ;
      RECT 19.505 1.635 19.675 1.805 ;
      RECT 19.045 -3.805 19.215 -3.635 ;
      RECT 19.045 -1.085 19.215 -0.915 ;
      RECT 19.045 1.635 19.215 1.805 ;
      RECT 19.035 -1.935 19.205 -1.765 ;
      RECT 18.585 -3.805 18.755 -3.635 ;
      RECT 18.585 -1.085 18.755 -0.915 ;
      RECT 18.585 1.635 18.755 1.805 ;
      RECT 18.525 0.445 18.695 0.615 ;
      RECT 17.17 -4.515 17.34 -4.345 ;
      RECT 17.17 -3.035 17.34 -2.865 ;
      RECT 17.17 0.885 17.34 1.055 ;
      RECT 17.17 2.365 17.34 2.535 ;
      RECT 16.82 -5.325 16.99 -5.155 ;
      RECT 16.82 -1.265 16.99 -1.095 ;
      RECT 16.82 -0.885 16.99 -0.715 ;
      RECT 16.82 3.175 16.99 3.345 ;
      RECT 16.8 -2.665 16.97 -2.495 ;
      RECT 16.8 0.515 16.97 0.685 ;
      RECT 16.18 -4.515 16.35 -4.345 ;
      RECT 16.18 -3.035 16.35 -2.865 ;
      RECT 16.18 0.885 16.35 1.055 ;
      RECT 16.18 2.365 16.35 2.535 ;
      RECT 15.83 -5.325 16 -5.155 ;
      RECT 15.83 -1.265 16 -1.095 ;
      RECT 15.83 -0.885 16 -0.715 ;
      RECT 15.83 3.175 16 3.345 ;
      RECT 15.81 -2.665 15.98 -2.495 ;
      RECT 15.81 0.515 15.98 0.685 ;
      RECT 15.125 -5.325 15.295 -5.155 ;
      RECT 15.125 -1.265 15.295 -1.095 ;
      RECT 15.125 -0.885 15.295 -0.715 ;
      RECT 15.125 3.175 15.295 3.345 ;
      RECT 14.815 -3.405 14.985 -3.235 ;
      RECT 14.815 1.255 14.985 1.425 ;
      RECT 14.445 -5.325 14.615 -5.155 ;
      RECT 14.445 3.175 14.615 3.345 ;
      RECT 14.385 -4.515 14.555 -4.345 ;
      RECT 14.385 -3.775 14.555 -3.605 ;
      RECT 14.385 1.625 14.555 1.795 ;
      RECT 14.385 2.365 14.555 2.535 ;
      RECT 14.01 -3.035 14.18 -2.865 ;
      RECT 14.01 0.885 14.18 1.055 ;
      RECT 13.765 -5.325 13.935 -5.155 ;
      RECT 13.765 3.175 13.935 3.345 ;
      RECT 13.085 -5.325 13.255 -5.155 ;
      RECT 13.085 3.175 13.255 3.345 ;
      RECT 13.015 -2.665 13.185 -2.495 ;
      RECT 13.015 0.515 13.185 0.685 ;
      RECT 11.32 -3.805 11.49 -3.635 ;
      RECT 11.32 -1.085 11.49 -0.915 ;
      RECT 11.32 1.635 11.49 1.805 ;
      RECT 10.86 -3.805 11.03 -3.635 ;
      RECT 10.86 -1.085 11.03 -0.915 ;
      RECT 10.86 1.635 11.03 1.805 ;
      RECT 10.82 -1.595 10.99 -1.425 ;
      RECT 10.82 0.445 10.99 0.615 ;
      RECT 10.48 -2.615 10.65 -2.445 ;
      RECT 10.4 -3.805 10.57 -3.635 ;
      RECT 10.4 -1.085 10.57 -0.915 ;
      RECT 10.4 1.635 10.57 1.805 ;
      RECT 10.14 1.125 10.31 1.295 ;
      RECT 9.97 0.445 10.14 0.615 ;
      RECT 9.94 -3.805 10.11 -3.635 ;
      RECT 9.94 -1.085 10.11 -0.915 ;
      RECT 9.94 1.635 10.11 1.805 ;
      RECT 9.48 -3.805 9.65 -3.635 ;
      RECT 9.48 -1.085 9.65 -0.915 ;
      RECT 9.48 1.635 9.65 1.805 ;
      RECT 9.46 0.445 9.63 0.615 ;
      RECT 9.02 -3.805 9.19 -3.635 ;
      RECT 9.02 -1.085 9.19 -0.915 ;
      RECT 9.02 1.635 9.19 1.805 ;
      RECT 8.78 -2.275 8.95 -2.105 ;
      RECT 8.78 1.125 8.95 1.295 ;
      RECT 8.56 -3.805 8.73 -3.635 ;
      RECT 8.56 -1.085 8.73 -0.915 ;
      RECT 8.56 1.635 8.73 1.805 ;
      RECT 8.1 -3.805 8.27 -3.635 ;
      RECT 8.1 -2.615 8.27 -2.445 ;
      RECT 8.1 -1.085 8.27 -0.915 ;
      RECT 8.1 1.635 8.27 1.805 ;
      RECT 8.09 0.445 8.26 0.615 ;
      RECT 7.64 -3.805 7.81 -3.635 ;
      RECT 7.64 -1.085 7.81 -0.915 ;
      RECT 7.64 -0.575 7.81 -0.405 ;
      RECT 7.64 1.635 7.81 1.805 ;
      RECT 7.62 -3.125 7.79 -2.955 ;
      RECT 7.25 -2.61 7.42 -2.44 ;
      RECT 7.18 -3.805 7.35 -3.635 ;
      RECT 7.18 -1.085 7.35 -0.915 ;
      RECT 7.18 1.635 7.35 1.805 ;
      RECT 6.74 -2.61 6.91 -2.44 ;
      RECT 6.74 -1.595 6.91 -1.425 ;
      RECT 6.74 0.445 6.91 0.615 ;
      RECT 6.72 -3.805 6.89 -3.635 ;
      RECT 6.72 -1.085 6.89 -0.915 ;
      RECT 6.72 1.635 6.89 1.805 ;
      RECT 6.4 1.125 6.57 1.295 ;
      RECT 6.26 -3.805 6.43 -3.635 ;
      RECT 6.26 -1.085 6.43 -0.915 ;
      RECT 6.26 1.635 6.43 1.805 ;
      RECT 5.8 -3.805 5.97 -3.635 ;
      RECT 5.8 -1.085 5.97 -0.915 ;
      RECT 5.8 1.635 5.97 1.805 ;
      RECT 5.38 -2.615 5.55 -2.445 ;
      RECT 5.38 -0.575 5.55 -0.405 ;
      RECT 5.34 -3.805 5.51 -3.635 ;
      RECT 5.34 -1.085 5.51 -0.915 ;
      RECT 5.34 1.635 5.51 1.805 ;
      RECT 4.88 -3.805 5.05 -3.635 ;
      RECT 4.88 -1.085 5.05 -0.915 ;
      RECT 4.88 1.635 5.05 1.805 ;
      RECT 4.87 -1.935 5.04 -1.765 ;
      RECT 4.42 -3.805 4.59 -3.635 ;
      RECT 4.42 -1.085 4.59 -0.915 ;
      RECT 4.42 1.635 4.59 1.805 ;
      RECT 4.36 0.445 4.53 0.615 ;
    LAYER li ;
      RECT 65.185 -5.42 65.475 -2.79 ;
      RECT 51.01 -5.42 51.3 -2.79 ;
      RECT 36.835 -5.42 37.125 -2.79 ;
      RECT 22.665 -5.43 22.955 -2.8 ;
      RECT 8.5 -5.43 8.79 -2.8 ;
      RECT 61.985 -5.42 62.215 -2.805 ;
      RECT 61.105 -5.42 61.315 -2.805 ;
      RECT 47.81 -5.42 48.04 -2.805 ;
      RECT 46.93 -5.42 47.14 -2.805 ;
      RECT 33.635 -5.42 33.865 -2.805 ;
      RECT 32.755 -5.42 32.965 -2.805 ;
      RECT 64.735 -5.42 65.005 -2.815 ;
      RECT 63.825 -5.42 64.065 -2.815 ;
      RECT 63.375 -5.42 63.615 -2.815 ;
      RECT 62.435 -5.42 62.705 -2.815 ;
      RECT 50.56 -5.42 50.83 -2.815 ;
      RECT 49.65 -5.42 49.89 -2.815 ;
      RECT 49.2 -5.42 49.44 -2.815 ;
      RECT 48.26 -5.42 48.53 -2.815 ;
      RECT 36.385 -5.42 36.655 -2.815 ;
      RECT 35.475 -5.42 35.715 -2.815 ;
      RECT 35.025 -5.42 35.265 -2.815 ;
      RECT 34.085 -5.42 34.355 -2.815 ;
      RECT 19.465 -5.43 19.695 -2.815 ;
      RECT 18.585 -5.43 18.795 -2.815 ;
      RECT 5.3 -5.43 5.53 -2.815 ;
      RECT 4.42 -5.43 4.63 -2.815 ;
      RECT 22.215 -5.43 22.485 -2.825 ;
      RECT 21.305 -5.43 21.545 -2.825 ;
      RECT 20.855 -5.43 21.095 -2.825 ;
      RECT 19.915 -5.43 20.185 -2.825 ;
      RECT 8.05 -5.43 8.32 -2.825 ;
      RECT 7.14 -5.43 7.38 -2.825 ;
      RECT 6.69 -5.43 6.93 -2.825 ;
      RECT 5.75 -5.43 6.02 -2.825 ;
      RECT 67.855 -5.42 68.185 -3.235 ;
      RECT 67.015 -5.42 67.345 -3.235 ;
      RECT 53.68 -5.42 54.01 -3.235 ;
      RECT 52.84 -5.42 53.17 -3.235 ;
      RECT 39.505 -5.42 39.835 -3.235 ;
      RECT 38.665 -5.42 38.995 -3.235 ;
      RECT 25.335 -5.43 25.665 -3.245 ;
      RECT 24.495 -5.43 24.825 -3.245 ;
      RECT 11.17 -5.43 11.5 -3.245 ;
      RECT 10.33 -5.43 10.66 -3.245 ;
      RECT 60.96 -5.42 68.615 -3.625 ;
      RECT 46.785 -5.42 54.44 -3.625 ;
      RECT 32.61 -5.42 40.265 -3.625 ;
      RECT 18.44 -5.43 26.095 -3.635 ;
      RECT 4.275 -5.43 11.93 -3.635 ;
      RECT 60.955 -5.42 68.615 -3.785 ;
      RECT 46.78 -5.42 54.44 -3.785 ;
      RECT 32.605 -5.42 40.265 -3.785 ;
      RECT 18.435 -5.43 26.095 -3.795 ;
      RECT 4.27 -5.43 11.93 -3.795 ;
      RECT 73.425 -5.42 73.595 -4.485 ;
      RECT 72.435 -5.42 72.605 -4.485 ;
      RECT 69.69 -5.42 69.86 -4.485 ;
      RECT 59.25 -5.42 59.42 -4.485 ;
      RECT 58.26 -5.42 58.43 -4.485 ;
      RECT 55.515 -5.42 55.685 -4.485 ;
      RECT 45.075 -5.42 45.245 -4.485 ;
      RECT 44.085 -5.42 44.255 -4.485 ;
      RECT 41.34 -5.42 41.51 -4.485 ;
      RECT 30.905 -5.43 31.075 -4.495 ;
      RECT 29.915 -5.43 30.085 -4.495 ;
      RECT 27.17 -5.43 27.34 -4.495 ;
      RECT 16.74 -5.43 16.91 -4.495 ;
      RECT 15.75 -5.43 15.92 -4.495 ;
      RECT 13.005 -5.43 13.175 -4.495 ;
      RECT 31.575 -5.42 74.395 -5.115 ;
      RECT 3.24 -5.43 31.875 -5.125 ;
      RECT 67.495 -1.075 67.775 0.235 ;
      RECT 66.565 -1.075 66.825 0.235 ;
      RECT 66.115 -1.075 66.395 0.235 ;
      RECT 65.185 -1.075 65.445 0.235 ;
      RECT 64.755 -1.075 65.015 0.235 ;
      RECT 63.805 -1.075 64.085 0.235 ;
      RECT 62.455 -2.215 62.715 0.235 ;
      RECT 61.505 -1.075 61.785 0.235 ;
      RECT 53.32 -1.075 53.6 0.235 ;
      RECT 52.39 -1.075 52.65 0.235 ;
      RECT 51.94 -1.075 52.22 0.235 ;
      RECT 51.01 -1.075 51.27 0.235 ;
      RECT 50.58 -1.075 50.84 0.235 ;
      RECT 49.63 -1.075 49.91 0.235 ;
      RECT 48.28 -2.215 48.54 0.235 ;
      RECT 47.33 -1.075 47.61 0.235 ;
      RECT 39.145 -1.075 39.425 0.235 ;
      RECT 38.215 -1.075 38.475 0.235 ;
      RECT 37.765 -1.075 38.045 0.235 ;
      RECT 36.835 -1.075 37.095 0.235 ;
      RECT 36.405 -1.075 36.665 0.235 ;
      RECT 35.455 -1.075 35.735 0.235 ;
      RECT 34.105 -2.215 34.365 0.235 ;
      RECT 33.155 -1.075 33.435 0.235 ;
      RECT 24.975 -1.085 25.255 0.225 ;
      RECT 24.045 -1.085 24.305 0.225 ;
      RECT 23.595 -1.085 23.875 0.225 ;
      RECT 22.665 -1.085 22.925 0.225 ;
      RECT 22.235 -1.085 22.495 0.225 ;
      RECT 21.285 -1.085 21.565 0.225 ;
      RECT 19.935 -2.225 20.195 0.225 ;
      RECT 18.985 -1.085 19.265 0.225 ;
      RECT 10.81 -1.085 11.09 0.225 ;
      RECT 9.88 -1.085 10.14 0.225 ;
      RECT 9.43 -1.085 9.71 0.225 ;
      RECT 8.5 -1.085 8.76 0.225 ;
      RECT 8.07 -1.085 8.33 0.225 ;
      RECT 7.12 -1.085 7.4 0.225 ;
      RECT 5.77 -2.225 6.03 0.225 ;
      RECT 4.82 -1.085 5.1 0.225 ;
      RECT 73.425 -2.015 73.595 0.055 ;
      RECT 72.435 -2.015 72.605 0.055 ;
      RECT 69.69 -2.015 69.86 0.055 ;
      RECT 59.25 -2.015 59.42 0.055 ;
      RECT 58.26 -2.015 58.43 0.055 ;
      RECT 55.515 -2.015 55.685 0.055 ;
      RECT 45.075 -2.015 45.245 0.055 ;
      RECT 44.085 -2.015 44.255 0.055 ;
      RECT 41.34 -2.015 41.51 0.055 ;
      RECT 30.905 -2.025 31.075 0.045 ;
      RECT 29.915 -2.025 30.085 0.045 ;
      RECT 27.17 -2.025 27.34 0.045 ;
      RECT 16.74 -2.025 16.91 0.045 ;
      RECT 15.75 -2.025 15.92 0.045 ;
      RECT 13.005 -2.025 13.175 0.045 ;
      RECT 68.41 -1.285 74.395 -0.675 ;
      RECT 54.235 -1.285 60.22 -0.675 ;
      RECT 40.06 -1.285 46.045 -0.675 ;
      RECT 54.235 -1.075 61.335 -0.68 ;
      RECT 40.06 -1.075 47.16 -0.68 ;
      RECT 31.575 -1.075 32.985 -0.68 ;
      RECT 25.89 -1.075 32.985 -0.685 ;
      RECT 11.725 -1.295 17.71 -0.685 ;
      RECT 11.725 -1.085 18.815 -0.69 ;
      RECT 3.24 -1.085 4.65 -0.69 ;
      RECT 25.89 -1.075 74.395 -0.905 ;
      RECT 68.405 -1.285 74.395 -0.905 ;
      RECT 25.885 -1.295 31.875 -0.915 ;
      RECT 67.095 -1.925 67.265 -0.905 ;
      RECT 66.255 -1.585 66.425 -0.905 ;
      RECT 64.675 -2.215 65.005 -0.905 ;
      RECT 62.435 -2.215 62.765 -0.905 ;
      RECT 61.985 -2.215 62.215 -0.905 ;
      RECT 54.23 -1.285 61.315 -0.905 ;
      RECT 61.105 -2.215 61.315 -0.68 ;
      RECT 52.92 -1.925 53.09 -0.905 ;
      RECT 52.08 -1.585 52.25 -0.905 ;
      RECT 50.5 -2.215 50.83 -0.905 ;
      RECT 48.26 -2.215 48.59 -0.905 ;
      RECT 47.81 -2.215 48.04 -0.905 ;
      RECT 40.055 -1.285 47.14 -0.905 ;
      RECT 46.93 -2.215 47.14 -0.68 ;
      RECT 38.745 -1.925 38.915 -0.905 ;
      RECT 37.905 -1.585 38.075 -0.905 ;
      RECT 36.325 -2.215 36.655 -0.905 ;
      RECT 34.085 -2.215 34.415 -0.905 ;
      RECT 33.635 -2.215 33.865 -0.905 ;
      RECT 3.24 -1.085 32.965 -0.915 ;
      RECT 32.755 -2.215 32.965 -0.68 ;
      RECT 25.885 -1.29 32.965 -0.915 ;
      RECT 24.575 -1.935 24.745 -0.915 ;
      RECT 23.735 -1.595 23.905 -0.915 ;
      RECT 22.155 -2.225 22.485 -0.915 ;
      RECT 19.915 -2.225 20.245 -0.915 ;
      RECT 19.465 -2.225 19.695 -0.915 ;
      RECT 11.72 -1.295 18.795 -0.915 ;
      RECT 18.585 -2.225 18.795 -0.69 ;
      RECT 10.41 -1.935 10.58 -0.915 ;
      RECT 9.57 -1.595 9.74 -0.915 ;
      RECT 7.99 -2.225 8.32 -0.915 ;
      RECT 5.75 -2.225 6.08 -0.915 ;
      RECT 5.3 -2.225 5.53 -0.915 ;
      RECT 3.24 -1.3 4.63 -0.69 ;
      RECT 4.42 -2.225 4.63 -0.69 ;
      RECT 59.925 -1.29 61.315 -0.68 ;
      RECT 45.75 -1.29 47.14 -0.68 ;
      RECT 17.405 -1.3 18.795 -0.69 ;
      RECT 31.575 3.155 74.395 3.46 ;
      RECT 3.24 3.145 31.875 3.45 ;
      RECT 73.425 2.525 73.595 3.46 ;
      RECT 72.435 2.525 72.605 3.46 ;
      RECT 69.69 2.525 69.86 3.46 ;
      RECT 61.23 1.76 68.43 3.46 ;
      RECT 59.25 2.525 59.42 3.46 ;
      RECT 58.26 2.525 58.43 3.46 ;
      RECT 55.515 2.525 55.685 3.46 ;
      RECT 47.055 1.76 54.255 3.46 ;
      RECT 45.075 2.525 45.245 3.46 ;
      RECT 44.085 2.525 44.255 3.46 ;
      RECT 41.34 2.525 41.51 3.46 ;
      RECT 32.88 1.76 40.08 3.46 ;
      RECT 30.905 2.515 31.075 3.45 ;
      RECT 29.915 2.515 30.085 3.45 ;
      RECT 27.17 2.515 27.34 3.45 ;
      RECT 18.71 1.75 25.91 3.45 ;
      RECT 16.74 2.515 16.91 3.45 ;
      RECT 15.75 2.515 15.92 3.45 ;
      RECT 13.005 2.515 13.175 3.45 ;
      RECT 4.545 1.75 11.745 3.45 ;
      RECT 60.96 1.645 68.32 1.815 ;
      RECT 46.785 1.645 54.145 1.815 ;
      RECT 32.61 1.645 39.97 1.815 ;
      RECT 18.44 1.635 25.8 1.805 ;
      RECT 4.275 1.635 11.635 1.805 ;
      RECT 67.465 0.845 67.775 3.46 ;
      RECT 66.085 0.845 66.395 3.46 ;
      RECT 63.805 0.845 64.115 3.46 ;
      RECT 61.505 0.845 61.815 3.46 ;
      RECT 53.29 0.845 53.6 3.46 ;
      RECT 51.91 0.845 52.22 3.46 ;
      RECT 49.63 0.845 49.94 3.46 ;
      RECT 47.33 0.845 47.64 3.46 ;
      RECT 39.115 0.845 39.425 3.46 ;
      RECT 37.735 0.845 38.045 3.46 ;
      RECT 35.455 0.845 35.765 3.46 ;
      RECT 33.155 0.845 33.465 3.46 ;
      RECT 24.945 0.835 25.255 3.45 ;
      RECT 23.565 0.835 23.875 3.45 ;
      RECT 21.285 0.835 21.595 3.45 ;
      RECT 18.985 0.835 19.295 3.45 ;
      RECT 10.78 0.835 11.09 3.45 ;
      RECT 9.4 0.835 9.71 3.45 ;
      RECT 7.12 0.835 7.43 3.45 ;
      RECT 4.82 0.835 5.13 3.45 ;
      RECT 73.485 -3.68 73.655 -2.485 ;
      RECT 73.485 -3.68 73.95 -3.51 ;
      RECT 73.485 1.55 73.95 1.72 ;
      RECT 73.485 0.525 73.655 1.72 ;
      RECT 72.495 -3.68 72.665 -2.485 ;
      RECT 72.495 -3.68 72.96 -3.51 ;
      RECT 72.495 1.55 72.96 1.72 ;
      RECT 72.495 0.525 72.665 1.72 ;
      RECT 70.64 -2.785 70.81 -1.555 ;
      RECT 70.695 -4.565 70.865 -2.615 ;
      RECT 70.64 -4.845 70.81 -4.395 ;
      RECT 70.64 2.435 70.81 2.885 ;
      RECT 70.695 0.655 70.865 2.605 ;
      RECT 70.64 -0.405 70.81 0.825 ;
      RECT 70.12 -4.845 70.29 -1.555 ;
      RECT 70.12 -3.345 70.525 -3.015 ;
      RECT 70.12 -4.185 70.525 -3.855 ;
      RECT 70.12 -0.405 70.29 2.885 ;
      RECT 70.12 1.895 70.525 2.225 ;
      RECT 70.12 1.055 70.525 1.385 ;
      RECT 67.855 -1.925 68.235 -1.245 ;
      RECT 68.065 -3.055 68.235 -1.245 ;
      RECT 65.985 -3.055 66.215 -2.385 ;
      RECT 65.985 -3.055 68.235 -2.885 ;
      RECT 67.515 -3.375 67.685 -2.885 ;
      RECT 67.505 -2.265 67.675 -1.415 ;
      RECT 66.59 -2.265 67.895 -2.095 ;
      RECT 67.65 -2.715 67.895 -2.095 ;
      RECT 66.59 -2.635 66.76 -2.095 ;
      RECT 66.385 -2.635 66.76 -2.465 ;
      RECT 66.565 0.845 67.26 1.475 ;
      RECT 67.09 -0.735 67.26 1.475 ;
      RECT 66.995 -0.735 67.325 0.245 ;
      RECT 66.595 -1.925 66.925 -1.245 ;
      RECT 65.685 -1.925 66.085 -1.245 ;
      RECT 65.685 -1.925 66.925 -1.755 ;
      RECT 65.185 -2.345 65.505 -1.245 ;
      RECT 65.185 -2.345 65.635 -2.095 ;
      RECT 65.185 -2.345 65.815 -2.175 ;
      RECT 65.645 -3.395 65.815 -2.175 ;
      RECT 65.645 -3.395 66.6 -3.225 ;
      RECT 65.185 0.845 65.88 1.475 ;
      RECT 65.71 -0.735 65.88 1.475 ;
      RECT 65.615 -0.735 65.945 0.245 ;
      RECT 65.205 0.405 65.54 0.655 ;
      RECT 64.66 0.405 64.995 0.655 ;
      RECT 64.66 0.455 65.54 0.625 ;
      RECT 64.32 0.845 65.015 1.475 ;
      RECT 64.32 -0.735 64.49 1.475 ;
      RECT 64.255 -0.735 64.585 0.245 ;
      RECT 63.815 -2.215 64.145 -1.26 ;
      RECT 63.815 -2.215 64.495 -2.045 ;
      RECT 64.325 -3.455 64.495 -2.045 ;
      RECT 64.235 -3.455 64.565 -2.815 ;
      RECT 63.815 0.405 64.15 0.675 ;
      RECT 63.425 0.455 64.15 0.625 ;
      RECT 63.295 -2.215 63.625 -1.26 ;
      RECT 62.945 -2.215 63.625 -2.045 ;
      RECT 62.945 -3.455 63.115 -2.045 ;
      RECT 62.875 -3.455 63.205 -2.815 ;
      RECT 63.085 0.455 63.255 1.305 ;
      RECT 62.36 0.405 62.695 0.655 ;
      RECT 62.36 0.455 63.255 0.625 ;
      RECT 62.425 -2.635 62.775 -2.385 ;
      RECT 61.905 -2.635 62.235 -2.385 ;
      RECT 61.905 -2.605 62.775 -2.435 ;
      RECT 62.02 0.845 62.715 1.475 ;
      RECT 62.02 -0.735 62.19 1.475 ;
      RECT 61.955 -0.735 62.285 0.245 ;
      RECT 61.515 0.405 61.85 0.675 ;
      RECT 61.045 0.455 61.85 0.625 ;
      RECT 61.485 -2.225 61.815 -1.245 ;
      RECT 61.485 -3.455 61.735 -1.245 ;
      RECT 61.485 -3.455 61.815 -2.825 ;
      RECT 59.31 -3.68 59.48 -2.485 ;
      RECT 59.31 -3.68 59.775 -3.51 ;
      RECT 59.31 1.55 59.775 1.72 ;
      RECT 59.31 0.525 59.48 1.72 ;
      RECT 58.32 -3.68 58.49 -2.485 ;
      RECT 58.32 -3.68 58.785 -3.51 ;
      RECT 58.32 1.55 58.785 1.72 ;
      RECT 58.32 0.525 58.49 1.72 ;
      RECT 56.465 -2.785 56.635 -1.555 ;
      RECT 56.52 -4.565 56.69 -2.615 ;
      RECT 56.465 -4.845 56.635 -4.395 ;
      RECT 56.465 2.435 56.635 2.885 ;
      RECT 56.52 0.655 56.69 2.605 ;
      RECT 56.465 -0.405 56.635 0.825 ;
      RECT 55.945 -4.845 56.115 -1.555 ;
      RECT 55.945 -3.345 56.35 -3.015 ;
      RECT 55.945 -4.185 56.35 -3.855 ;
      RECT 55.945 -0.405 56.115 2.885 ;
      RECT 55.945 1.895 56.35 2.225 ;
      RECT 55.945 1.055 56.35 1.385 ;
      RECT 53.68 -1.925 54.06 -1.245 ;
      RECT 53.89 -3.055 54.06 -1.245 ;
      RECT 51.81 -3.055 52.04 -2.385 ;
      RECT 51.81 -3.055 54.06 -2.885 ;
      RECT 53.34 -3.375 53.51 -2.885 ;
      RECT 53.33 -2.265 53.5 -1.415 ;
      RECT 52.415 -2.265 53.72 -2.095 ;
      RECT 53.475 -2.715 53.72 -2.095 ;
      RECT 52.415 -2.635 52.585 -2.095 ;
      RECT 52.21 -2.635 52.585 -2.465 ;
      RECT 52.39 0.845 53.085 1.475 ;
      RECT 52.915 -0.735 53.085 1.475 ;
      RECT 52.82 -0.735 53.15 0.245 ;
      RECT 52.42 -1.925 52.75 -1.245 ;
      RECT 51.51 -1.925 51.91 -1.245 ;
      RECT 51.51 -1.925 52.75 -1.755 ;
      RECT 51.01 -2.345 51.33 -1.245 ;
      RECT 51.01 -2.345 51.46 -2.095 ;
      RECT 51.01 -2.345 51.64 -2.175 ;
      RECT 51.47 -3.395 51.64 -2.175 ;
      RECT 51.47 -3.395 52.425 -3.225 ;
      RECT 51.01 0.845 51.705 1.475 ;
      RECT 51.535 -0.735 51.705 1.475 ;
      RECT 51.44 -0.735 51.77 0.245 ;
      RECT 51.03 0.405 51.365 0.655 ;
      RECT 50.485 0.405 50.82 0.655 ;
      RECT 50.485 0.455 51.365 0.625 ;
      RECT 50.145 0.845 50.84 1.475 ;
      RECT 50.145 -0.735 50.315 1.475 ;
      RECT 50.08 -0.735 50.41 0.245 ;
      RECT 49.64 -2.215 49.97 -1.26 ;
      RECT 49.64 -2.215 50.32 -2.045 ;
      RECT 50.15 -3.455 50.32 -2.045 ;
      RECT 50.06 -3.455 50.39 -2.815 ;
      RECT 49.64 0.405 49.975 0.675 ;
      RECT 49.25 0.455 49.975 0.625 ;
      RECT 49.12 -2.215 49.45 -1.26 ;
      RECT 48.77 -2.215 49.45 -2.045 ;
      RECT 48.77 -3.455 48.94 -2.045 ;
      RECT 48.7 -3.455 49.03 -2.815 ;
      RECT 48.91 0.455 49.08 1.305 ;
      RECT 48.185 0.405 48.52 0.655 ;
      RECT 48.185 0.455 49.08 0.625 ;
      RECT 48.25 -2.635 48.6 -2.385 ;
      RECT 47.73 -2.635 48.06 -2.385 ;
      RECT 47.73 -2.605 48.6 -2.435 ;
      RECT 47.845 0.845 48.54 1.475 ;
      RECT 47.845 -0.735 48.015 1.475 ;
      RECT 47.78 -0.735 48.11 0.245 ;
      RECT 47.34 0.405 47.675 0.675 ;
      RECT 46.87 0.455 47.675 0.625 ;
      RECT 47.31 -2.225 47.64 -1.245 ;
      RECT 47.31 -3.455 47.56 -1.245 ;
      RECT 47.31 -3.455 47.64 -2.825 ;
      RECT 45.135 -3.68 45.305 -2.485 ;
      RECT 45.135 -3.68 45.6 -3.51 ;
      RECT 45.135 1.55 45.6 1.72 ;
      RECT 45.135 0.525 45.305 1.72 ;
      RECT 44.145 -3.68 44.315 -2.485 ;
      RECT 44.145 -3.68 44.61 -3.51 ;
      RECT 44.145 1.55 44.61 1.72 ;
      RECT 44.145 0.525 44.315 1.72 ;
      RECT 42.29 -2.785 42.46 -1.555 ;
      RECT 42.345 -4.565 42.515 -2.615 ;
      RECT 42.29 -4.845 42.46 -4.395 ;
      RECT 42.29 2.435 42.46 2.885 ;
      RECT 42.345 0.655 42.515 2.605 ;
      RECT 42.29 -0.405 42.46 0.825 ;
      RECT 41.77 -4.845 41.94 -1.555 ;
      RECT 41.77 -3.345 42.175 -3.015 ;
      RECT 41.77 -4.185 42.175 -3.855 ;
      RECT 41.77 -0.405 41.94 2.885 ;
      RECT 41.77 1.895 42.175 2.225 ;
      RECT 41.77 1.055 42.175 1.385 ;
      RECT 39.505 -1.925 39.885 -1.245 ;
      RECT 39.715 -3.055 39.885 -1.245 ;
      RECT 37.635 -3.055 37.865 -2.385 ;
      RECT 37.635 -3.055 39.885 -2.885 ;
      RECT 39.165 -3.375 39.335 -2.885 ;
      RECT 39.155 -2.265 39.325 -1.415 ;
      RECT 38.24 -2.265 39.545 -2.095 ;
      RECT 39.3 -2.715 39.545 -2.095 ;
      RECT 38.24 -2.635 38.41 -2.095 ;
      RECT 38.035 -2.635 38.41 -2.465 ;
      RECT 38.215 0.845 38.91 1.475 ;
      RECT 38.74 -0.735 38.91 1.475 ;
      RECT 38.645 -0.735 38.975 0.245 ;
      RECT 38.245 -1.925 38.575 -1.245 ;
      RECT 37.335 -1.925 37.735 -1.245 ;
      RECT 37.335 -1.925 38.575 -1.755 ;
      RECT 36.835 -2.345 37.155 -1.245 ;
      RECT 36.835 -2.345 37.285 -2.095 ;
      RECT 36.835 -2.345 37.465 -2.175 ;
      RECT 37.295 -3.395 37.465 -2.175 ;
      RECT 37.295 -3.395 38.25 -3.225 ;
      RECT 36.835 0.845 37.53 1.475 ;
      RECT 37.36 -0.735 37.53 1.475 ;
      RECT 37.265 -0.735 37.595 0.245 ;
      RECT 36.855 0.405 37.19 0.655 ;
      RECT 36.31 0.405 36.645 0.655 ;
      RECT 36.31 0.455 37.19 0.625 ;
      RECT 35.97 0.845 36.665 1.475 ;
      RECT 35.97 -0.735 36.14 1.475 ;
      RECT 35.905 -0.735 36.235 0.245 ;
      RECT 35.465 -2.215 35.795 -1.26 ;
      RECT 35.465 -2.215 36.145 -2.045 ;
      RECT 35.975 -3.455 36.145 -2.045 ;
      RECT 35.885 -3.455 36.215 -2.815 ;
      RECT 35.465 0.405 35.8 0.675 ;
      RECT 35.075 0.455 35.8 0.625 ;
      RECT 34.945 -2.215 35.275 -1.26 ;
      RECT 34.595 -2.215 35.275 -2.045 ;
      RECT 34.595 -3.455 34.765 -2.045 ;
      RECT 34.525 -3.455 34.855 -2.815 ;
      RECT 34.735 0.455 34.905 1.305 ;
      RECT 34.01 0.405 34.345 0.655 ;
      RECT 34.01 0.455 34.905 0.625 ;
      RECT 34.075 -2.635 34.425 -2.385 ;
      RECT 33.555 -2.635 33.885 -2.385 ;
      RECT 33.555 -2.605 34.425 -2.435 ;
      RECT 33.67 0.845 34.365 1.475 ;
      RECT 33.67 -0.735 33.84 1.475 ;
      RECT 33.605 -0.735 33.935 0.245 ;
      RECT 33.165 0.405 33.5 0.675 ;
      RECT 32.695 0.455 33.5 0.625 ;
      RECT 33.135 -2.225 33.465 -1.245 ;
      RECT 33.135 -3.455 33.385 -1.245 ;
      RECT 33.135 -3.455 33.465 -2.825 ;
      RECT 30.965 -3.69 31.135 -2.495 ;
      RECT 30.965 -3.69 31.43 -3.52 ;
      RECT 30.965 1.54 31.43 1.71 ;
      RECT 30.965 0.515 31.135 1.71 ;
      RECT 29.975 -3.69 30.145 -2.495 ;
      RECT 29.975 -3.69 30.44 -3.52 ;
      RECT 29.975 1.54 30.44 1.71 ;
      RECT 29.975 0.515 30.145 1.71 ;
      RECT 28.12 -2.795 28.29 -1.565 ;
      RECT 28.175 -4.575 28.345 -2.625 ;
      RECT 28.12 -4.855 28.29 -4.405 ;
      RECT 28.12 2.425 28.29 2.875 ;
      RECT 28.175 0.645 28.345 2.595 ;
      RECT 28.12 -0.415 28.29 0.815 ;
      RECT 27.6 -4.855 27.77 -1.565 ;
      RECT 27.6 -3.355 28.005 -3.025 ;
      RECT 27.6 -4.195 28.005 -3.865 ;
      RECT 27.6 -0.415 27.77 2.875 ;
      RECT 27.6 1.885 28.005 2.215 ;
      RECT 27.6 1.045 28.005 1.375 ;
      RECT 25.335 -1.935 25.715 -1.255 ;
      RECT 25.545 -3.065 25.715 -1.255 ;
      RECT 23.465 -3.065 23.695 -2.395 ;
      RECT 23.465 -3.065 25.715 -2.895 ;
      RECT 24.995 -3.385 25.165 -2.895 ;
      RECT 24.985 -2.275 25.155 -1.425 ;
      RECT 24.07 -2.275 25.375 -2.105 ;
      RECT 25.13 -2.725 25.375 -2.105 ;
      RECT 24.07 -2.645 24.24 -2.105 ;
      RECT 23.865 -2.645 24.24 -2.475 ;
      RECT 24.045 0.835 24.74 1.465 ;
      RECT 24.57 -0.745 24.74 1.465 ;
      RECT 24.475 -0.745 24.805 0.235 ;
      RECT 24.075 -1.935 24.405 -1.255 ;
      RECT 23.165 -1.935 23.565 -1.255 ;
      RECT 23.165 -1.935 24.405 -1.765 ;
      RECT 22.665 -2.355 22.985 -1.255 ;
      RECT 22.665 -2.355 23.115 -2.105 ;
      RECT 22.665 -2.355 23.295 -2.185 ;
      RECT 23.125 -3.405 23.295 -2.185 ;
      RECT 23.125 -3.405 24.08 -3.235 ;
      RECT 22.665 0.835 23.36 1.465 ;
      RECT 23.19 -0.745 23.36 1.465 ;
      RECT 23.095 -0.745 23.425 0.235 ;
      RECT 22.685 0.395 23.02 0.645 ;
      RECT 22.14 0.395 22.475 0.645 ;
      RECT 22.14 0.445 23.02 0.615 ;
      RECT 21.8 0.835 22.495 1.465 ;
      RECT 21.8 -0.745 21.97 1.465 ;
      RECT 21.735 -0.745 22.065 0.235 ;
      RECT 21.295 -2.225 21.625 -1.27 ;
      RECT 21.295 -2.225 21.975 -2.055 ;
      RECT 21.805 -3.465 21.975 -2.055 ;
      RECT 21.715 -3.465 22.045 -2.825 ;
      RECT 21.295 0.395 21.63 0.665 ;
      RECT 20.905 0.445 21.63 0.615 ;
      RECT 20.775 -2.225 21.105 -1.27 ;
      RECT 20.425 -2.225 21.105 -2.055 ;
      RECT 20.425 -3.465 20.595 -2.055 ;
      RECT 20.355 -3.465 20.685 -2.825 ;
      RECT 20.565 0.445 20.735 1.295 ;
      RECT 19.84 0.395 20.175 0.645 ;
      RECT 19.84 0.445 20.735 0.615 ;
      RECT 19.905 -2.645 20.255 -2.395 ;
      RECT 19.385 -2.645 19.715 -2.395 ;
      RECT 19.385 -2.615 20.255 -2.445 ;
      RECT 19.5 0.835 20.195 1.465 ;
      RECT 19.5 -0.745 19.67 1.465 ;
      RECT 19.435 -0.745 19.765 0.235 ;
      RECT 18.995 0.395 19.33 0.665 ;
      RECT 18.525 0.445 19.33 0.615 ;
      RECT 18.965 -2.235 19.295 -1.255 ;
      RECT 18.965 -3.465 19.215 -1.255 ;
      RECT 18.965 -3.465 19.295 -2.835 ;
      RECT 16.8 -3.69 16.97 -2.495 ;
      RECT 16.8 -3.69 17.265 -3.52 ;
      RECT 16.8 1.54 17.265 1.71 ;
      RECT 16.8 0.515 16.97 1.71 ;
      RECT 15.81 -3.69 15.98 -2.495 ;
      RECT 15.81 -3.69 16.275 -3.52 ;
      RECT 15.81 1.54 16.275 1.71 ;
      RECT 15.81 0.515 15.98 1.71 ;
      RECT 13.955 -2.795 14.125 -1.565 ;
      RECT 14.01 -4.575 14.18 -2.625 ;
      RECT 13.955 -4.855 14.125 -4.405 ;
      RECT 13.955 2.425 14.125 2.875 ;
      RECT 14.01 0.645 14.18 2.595 ;
      RECT 13.955 -0.415 14.125 0.815 ;
      RECT 13.435 -4.855 13.605 -1.565 ;
      RECT 13.435 -3.355 13.84 -3.025 ;
      RECT 13.435 -4.195 13.84 -3.865 ;
      RECT 13.435 -0.415 13.605 2.875 ;
      RECT 13.435 1.885 13.84 2.215 ;
      RECT 13.435 1.045 13.84 1.375 ;
      RECT 11.17 -1.935 11.55 -1.255 ;
      RECT 11.38 -3.065 11.55 -1.255 ;
      RECT 9.3 -3.065 9.53 -2.395 ;
      RECT 9.3 -3.065 11.55 -2.895 ;
      RECT 10.83 -3.385 11 -2.895 ;
      RECT 10.82 -2.275 10.99 -1.425 ;
      RECT 9.905 -2.275 11.21 -2.105 ;
      RECT 10.965 -2.725 11.21 -2.105 ;
      RECT 9.905 -2.645 10.075 -2.105 ;
      RECT 9.7 -2.645 10.075 -2.475 ;
      RECT 9.88 0.835 10.575 1.465 ;
      RECT 10.405 -0.745 10.575 1.465 ;
      RECT 10.31 -0.745 10.64 0.235 ;
      RECT 9.91 -1.935 10.24 -1.255 ;
      RECT 9 -1.935 9.4 -1.255 ;
      RECT 9 -1.935 10.24 -1.765 ;
      RECT 8.5 -2.355 8.82 -1.255 ;
      RECT 8.5 -2.355 8.95 -2.105 ;
      RECT 8.5 -2.355 9.13 -2.185 ;
      RECT 8.96 -3.405 9.13 -2.185 ;
      RECT 8.96 -3.405 9.915 -3.235 ;
      RECT 8.5 0.835 9.195 1.465 ;
      RECT 9.025 -0.745 9.195 1.465 ;
      RECT 8.93 -0.745 9.26 0.235 ;
      RECT 8.52 0.395 8.855 0.645 ;
      RECT 7.975 0.395 8.31 0.645 ;
      RECT 7.975 0.445 8.855 0.615 ;
      RECT 7.635 0.835 8.33 1.465 ;
      RECT 7.635 -0.745 7.805 1.465 ;
      RECT 7.57 -0.745 7.9 0.235 ;
      RECT 7.13 -2.225 7.46 -1.27 ;
      RECT 7.13 -2.225 7.81 -2.055 ;
      RECT 7.64 -3.465 7.81 -2.055 ;
      RECT 7.55 -3.465 7.88 -2.825 ;
      RECT 7.13 0.395 7.465 0.665 ;
      RECT 6.74 0.445 7.465 0.615 ;
      RECT 6.61 -2.225 6.94 -1.27 ;
      RECT 6.26 -2.225 6.94 -2.055 ;
      RECT 6.26 -3.465 6.43 -2.055 ;
      RECT 6.19 -3.465 6.52 -2.825 ;
      RECT 6.4 0.445 6.57 1.295 ;
      RECT 5.675 0.395 6.01 0.645 ;
      RECT 5.675 0.445 6.57 0.615 ;
      RECT 5.74 -2.645 6.09 -2.395 ;
      RECT 5.22 -2.645 5.55 -2.395 ;
      RECT 5.22 -2.615 6.09 -2.445 ;
      RECT 5.335 0.835 6.03 1.465 ;
      RECT 5.335 -0.745 5.505 1.465 ;
      RECT 5.27 -0.745 5.6 0.235 ;
      RECT 4.83 0.395 5.165 0.665 ;
      RECT 4.36 0.445 5.165 0.615 ;
      RECT 4.8 -2.235 5.13 -1.255 ;
      RECT 4.8 -3.465 5.05 -1.255 ;
      RECT 4.8 -3.465 5.13 -2.835 ;
      RECT 73.855 -4.845 74.025 -4.335 ;
      RECT 73.855 -3.025 74.025 -1.555 ;
      RECT 73.855 -0.405 74.025 1.065 ;
      RECT 73.855 2.375 74.025 2.885 ;
      RECT 72.865 -4.845 73.035 -4.335 ;
      RECT 72.865 -3.025 73.035 -1.555 ;
      RECT 72.865 -0.405 73.035 1.065 ;
      RECT 72.865 2.375 73.035 2.885 ;
      RECT 71.5 -4.845 71.67 -1.555 ;
      RECT 71.5 -0.405 71.67 2.885 ;
      RECT 71.07 -4.845 71.24 -4.335 ;
      RECT 71.07 -3.765 71.24 -1.555 ;
      RECT 71.07 -0.405 71.24 1.805 ;
      RECT 71.07 2.375 71.24 2.885 ;
      RECT 69.7 -3.76 69.87 -2.485 ;
      RECT 69.7 0.525 69.87 1.8 ;
      RECT 67.43 0.405 67.765 0.675 ;
      RECT 66.93 -2.635 67.48 -2.435 ;
      RECT 66.585 0.405 66.92 0.655 ;
      RECT 66.05 0.405 66.385 0.675 ;
      RECT 64.665 -2.635 65.015 -2.385 ;
      RECT 63.805 -2.635 64.155 -2.385 ;
      RECT 63.285 -2.635 63.635 -2.385 ;
      RECT 59.68 -4.845 59.85 -4.335 ;
      RECT 59.68 -3.025 59.85 -1.555 ;
      RECT 59.68 -0.405 59.85 1.065 ;
      RECT 59.68 2.375 59.85 2.885 ;
      RECT 58.69 -4.845 58.86 -4.335 ;
      RECT 58.69 -3.025 58.86 -1.555 ;
      RECT 58.69 -0.405 58.86 1.065 ;
      RECT 58.69 2.375 58.86 2.885 ;
      RECT 57.325 -4.845 57.495 -1.555 ;
      RECT 57.325 -0.405 57.495 2.885 ;
      RECT 56.895 -4.845 57.065 -4.335 ;
      RECT 56.895 -3.765 57.065 -1.555 ;
      RECT 56.895 -0.405 57.065 1.805 ;
      RECT 56.895 2.375 57.065 2.885 ;
      RECT 55.525 -3.76 55.695 -2.485 ;
      RECT 55.525 0.525 55.695 1.8 ;
      RECT 53.255 0.405 53.59 0.675 ;
      RECT 52.755 -2.635 53.305 -2.435 ;
      RECT 52.41 0.405 52.745 0.655 ;
      RECT 51.875 0.405 52.21 0.675 ;
      RECT 50.49 -2.635 50.84 -2.385 ;
      RECT 49.63 -2.635 49.98 -2.385 ;
      RECT 49.11 -2.635 49.46 -2.385 ;
      RECT 45.505 -4.845 45.675 -4.335 ;
      RECT 45.505 -3.025 45.675 -1.555 ;
      RECT 45.505 -0.405 45.675 1.065 ;
      RECT 45.505 2.375 45.675 2.885 ;
      RECT 44.515 -4.845 44.685 -4.335 ;
      RECT 44.515 -3.025 44.685 -1.555 ;
      RECT 44.515 -0.405 44.685 1.065 ;
      RECT 44.515 2.375 44.685 2.885 ;
      RECT 43.15 -4.845 43.32 -1.555 ;
      RECT 43.15 -0.405 43.32 2.885 ;
      RECT 42.72 -4.845 42.89 -4.335 ;
      RECT 42.72 -3.765 42.89 -1.555 ;
      RECT 42.72 -0.405 42.89 1.805 ;
      RECT 42.72 2.375 42.89 2.885 ;
      RECT 41.35 -3.76 41.52 -2.485 ;
      RECT 41.35 0.525 41.52 1.8 ;
      RECT 39.08 0.405 39.415 0.675 ;
      RECT 38.58 -2.635 39.13 -2.435 ;
      RECT 38.235 0.405 38.57 0.655 ;
      RECT 37.7 0.405 38.035 0.675 ;
      RECT 36.315 -2.635 36.665 -2.385 ;
      RECT 35.455 -2.635 35.805 -2.385 ;
      RECT 34.935 -2.635 35.285 -2.385 ;
      RECT 31.335 -4.855 31.505 -4.345 ;
      RECT 31.335 -3.035 31.505 -1.565 ;
      RECT 31.335 -0.415 31.505 1.055 ;
      RECT 31.335 2.365 31.505 2.875 ;
      RECT 30.345 -4.855 30.515 -4.345 ;
      RECT 30.345 -3.035 30.515 -1.565 ;
      RECT 30.345 -0.415 30.515 1.055 ;
      RECT 30.345 2.365 30.515 2.875 ;
      RECT 28.98 -4.855 29.15 -1.565 ;
      RECT 28.98 -0.415 29.15 2.875 ;
      RECT 28.55 -4.855 28.72 -4.345 ;
      RECT 28.55 -3.775 28.72 -1.565 ;
      RECT 28.55 -0.415 28.72 1.795 ;
      RECT 28.55 2.365 28.72 2.875 ;
      RECT 27.18 -3.77 27.35 -2.495 ;
      RECT 27.18 0.515 27.35 1.79 ;
      RECT 24.91 0.395 25.245 0.665 ;
      RECT 24.41 -2.645 24.96 -2.445 ;
      RECT 24.065 0.395 24.4 0.645 ;
      RECT 23.53 0.395 23.865 0.665 ;
      RECT 22.145 -2.645 22.495 -2.395 ;
      RECT 21.285 -2.645 21.635 -2.395 ;
      RECT 20.765 -2.645 21.115 -2.395 ;
      RECT 17.17 -4.855 17.34 -4.345 ;
      RECT 17.17 -3.035 17.34 -1.565 ;
      RECT 17.17 -0.415 17.34 1.055 ;
      RECT 17.17 2.365 17.34 2.875 ;
      RECT 16.18 -4.855 16.35 -4.345 ;
      RECT 16.18 -3.035 16.35 -1.565 ;
      RECT 16.18 -0.415 16.35 1.055 ;
      RECT 16.18 2.365 16.35 2.875 ;
      RECT 14.815 -4.855 14.985 -1.565 ;
      RECT 14.815 -0.415 14.985 2.875 ;
      RECT 14.385 -4.855 14.555 -4.345 ;
      RECT 14.385 -3.775 14.555 -1.565 ;
      RECT 14.385 -0.415 14.555 1.795 ;
      RECT 14.385 2.365 14.555 2.875 ;
      RECT 13.015 -3.77 13.185 -2.495 ;
      RECT 13.015 0.515 13.185 1.79 ;
      RECT 10.745 0.395 11.08 0.665 ;
      RECT 10.245 -2.645 10.795 -2.445 ;
      RECT 9.9 0.395 10.235 0.645 ;
      RECT 9.365 0.395 9.7 0.665 ;
      RECT 7.98 -2.645 8.33 -2.395 ;
      RECT 7.12 -2.645 7.47 -2.395 ;
      RECT 6.6 -2.645 6.95 -2.395 ;
  END
END sky130_osu_ring_oscillator_mpr2ct_8

MACRO sky130_osu_ring_oscillator_mpr2ea_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ea_8 0 0 ;
  SIZE 81.625 BY 8.88 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT 70.91 3.535 71.24 3.865 ;
      RECT 69.705 3.55 71.24 3.85 ;
      RECT 69.705 2.43 70.005 3.85 ;
      RECT 69.45 2.415 69.78 2.745 ;
      RECT 54.585 3.535 54.915 3.865 ;
      RECT 53.38 3.55 54.915 3.85 ;
      RECT 53.38 2.43 53.68 3.85 ;
      RECT 53.125 2.415 53.455 2.745 ;
      RECT 38.265 3.535 38.595 3.865 ;
      RECT 37.06 3.55 38.595 3.85 ;
      RECT 37.06 2.43 37.36 3.85 ;
      RECT 36.805 2.415 37.135 2.745 ;
      RECT 21.94 3.535 22.27 3.865 ;
      RECT 20.735 3.55 22.27 3.85 ;
      RECT 20.735 2.43 21.035 3.85 ;
      RECT 20.48 2.415 20.81 2.745 ;
      RECT 5.62 3.535 5.95 3.865 ;
      RECT 4.415 3.55 5.95 3.85 ;
      RECT 4.415 2.43 4.715 3.85 ;
      RECT 4.16 2.415 4.49 2.745 ;
      RECT 74.93 2.975 75.26 3.705 ;
      RECT 74.45 1.85 74.78 2.58 ;
      RECT 72.85 2.575 73.18 3.305 ;
      RECT 71.29 2.015 71.62 2.745 ;
      RECT 70.41 2.015 70.74 2.745 ;
      RECT 68.73 2.415 69.06 3.145 ;
      RECT 67.73 1.855 68.06 2.585 ;
      RECT 66.29 2.575 66.62 3.305 ;
      RECT 58.605 2.975 58.935 3.705 ;
      RECT 58.125 1.85 58.455 2.58 ;
      RECT 56.525 2.575 56.855 3.305 ;
      RECT 54.965 2.015 55.295 2.745 ;
      RECT 54.085 2.015 54.415 2.745 ;
      RECT 52.405 2.415 52.735 3.145 ;
      RECT 51.405 1.855 51.735 2.585 ;
      RECT 49.965 2.575 50.295 3.305 ;
      RECT 42.285 2.975 42.615 3.705 ;
      RECT 41.805 1.85 42.135 2.58 ;
      RECT 40.205 2.575 40.535 3.305 ;
      RECT 38.645 2.015 38.975 2.745 ;
      RECT 37.765 2.015 38.095 2.745 ;
      RECT 36.085 2.415 36.415 3.145 ;
      RECT 35.085 1.855 35.415 2.585 ;
      RECT 33.645 2.575 33.975 3.305 ;
      RECT 25.96 2.975 26.29 3.705 ;
      RECT 25.48 1.85 25.81 2.58 ;
      RECT 23.88 2.575 24.21 3.305 ;
      RECT 22.32 2.015 22.65 2.745 ;
      RECT 21.44 2.015 21.77 2.745 ;
      RECT 19.76 2.415 20.09 3.145 ;
      RECT 18.76 1.855 19.09 2.585 ;
      RECT 17.32 2.575 17.65 3.305 ;
      RECT 9.64 2.975 9.97 3.705 ;
      RECT 9.16 1.85 9.49 2.58 ;
      RECT 7.56 2.575 7.89 3.305 ;
      RECT 6 2.015 6.33 2.745 ;
      RECT 5.12 2.015 5.45 2.745 ;
      RECT 3.44 2.415 3.77 3.145 ;
      RECT 2.44 1.855 2.77 2.585 ;
      RECT 1 2.575 1.33 3.305 ;
    LAYER via2 ;
      RECT 74.995 3.04 75.195 3.24 ;
      RECT 74.515 2.315 74.715 2.515 ;
      RECT 72.915 3.04 73.115 3.24 ;
      RECT 71.355 2.48 71.555 2.68 ;
      RECT 70.975 3.6 71.175 3.8 ;
      RECT 70.475 2.48 70.675 2.68 ;
      RECT 69.515 2.48 69.715 2.68 ;
      RECT 68.795 2.48 68.995 2.68 ;
      RECT 67.795 1.92 67.995 2.12 ;
      RECT 66.355 3.04 66.555 3.24 ;
      RECT 58.67 3.04 58.87 3.24 ;
      RECT 58.19 2.315 58.39 2.515 ;
      RECT 56.59 3.04 56.79 3.24 ;
      RECT 55.03 2.48 55.23 2.68 ;
      RECT 54.65 3.6 54.85 3.8 ;
      RECT 54.15 2.48 54.35 2.68 ;
      RECT 53.19 2.48 53.39 2.68 ;
      RECT 52.47 2.48 52.67 2.68 ;
      RECT 51.47 1.92 51.67 2.12 ;
      RECT 50.03 3.04 50.23 3.24 ;
      RECT 42.35 3.04 42.55 3.24 ;
      RECT 41.87 2.315 42.07 2.515 ;
      RECT 40.27 3.04 40.47 3.24 ;
      RECT 38.71 2.48 38.91 2.68 ;
      RECT 38.33 3.6 38.53 3.8 ;
      RECT 37.83 2.48 38.03 2.68 ;
      RECT 36.87 2.48 37.07 2.68 ;
      RECT 36.15 2.48 36.35 2.68 ;
      RECT 35.15 1.92 35.35 2.12 ;
      RECT 33.71 3.04 33.91 3.24 ;
      RECT 26.025 3.04 26.225 3.24 ;
      RECT 25.545 2.315 25.745 2.515 ;
      RECT 23.945 3.04 24.145 3.24 ;
      RECT 22.385 2.48 22.585 2.68 ;
      RECT 22.005 3.6 22.205 3.8 ;
      RECT 21.505 2.48 21.705 2.68 ;
      RECT 20.545 2.48 20.745 2.68 ;
      RECT 19.825 2.48 20.025 2.68 ;
      RECT 18.825 1.92 19.025 2.12 ;
      RECT 17.385 3.04 17.585 3.24 ;
      RECT 9.705 3.04 9.905 3.24 ;
      RECT 9.225 2.315 9.425 2.515 ;
      RECT 7.625 3.04 7.825 3.24 ;
      RECT 6.065 2.48 6.265 2.68 ;
      RECT 5.685 3.6 5.885 3.8 ;
      RECT 5.185 2.48 5.385 2.68 ;
      RECT 4.225 2.48 4.425 2.68 ;
      RECT 3.505 2.48 3.705 2.68 ;
      RECT 2.505 1.92 2.705 2.12 ;
      RECT 1.065 3.04 1.265 3.24 ;
    LAYER met2 ;
      RECT 12.605 6.28 12.925 6.605 ;
      RECT 12.635 5.695 12.805 6.605 ;
      RECT 12.635 5.695 12.81 6.045 ;
      RECT 12.635 5.695 13.61 5.87 ;
      RECT 13.435 1.965 13.61 5.87 ;
      RECT 9.665 2.955 9.945 3.325 ;
      RECT 9.665 3.01 10.555 3.175 ;
      RECT 10.39 2.025 10.555 3.175 ;
      RECT 9.675 2.7 9.935 3.325 ;
      RECT 13.38 1.965 13.73 2.315 ;
      RECT 10.39 2.04 13.73 2.195 ;
      RECT 11.335 2.025 13.73 2.195 ;
      RECT 10.39 2.025 10.97 2.195 ;
      RECT 11.63 0.305 11.815 2.195 ;
      RECT 81.055 1.095 81.395 1.445 ;
      RECT 81.085 0.305 81.27 1.445 ;
      RECT 11.63 0.305 81.27 0.49 ;
      RECT 77.895 6.28 78.215 6.605 ;
      RECT 77.925 5.695 78.095 6.605 ;
      RECT 77.925 5.695 78.1 6.045 ;
      RECT 77.925 5.695 78.9 5.87 ;
      RECT 78.725 1.965 78.9 5.87 ;
      RECT 74.955 2.955 75.235 3.325 ;
      RECT 74.955 3.01 75.845 3.175 ;
      RECT 75.68 2.025 75.845 3.175 ;
      RECT 74.965 2.7 75.225 3.325 ;
      RECT 78.67 1.965 79.02 2.315 ;
      RECT 75.68 2.04 79.02 2.195 ;
      RECT 76.625 2.025 79.02 2.195 ;
      RECT 75.68 2.025 76.26 2.195 ;
      RECT 76.91 0.81 77.095 2.195 ;
      RECT 64.73 1.095 65.07 1.445 ;
      RECT 64.73 1.125 65.54 1.31 ;
      RECT 65.355 0.81 65.54 1.31 ;
      RECT 65.355 0.81 77.095 0.995 ;
      RECT 78.695 6.655 79.02 6.98 ;
      RECT 77.58 6.745 79.02 6.915 ;
      RECT 77.58 2.395 77.74 6.915 ;
      RECT 77.895 2.365 78.215 2.685 ;
      RECT 77.58 2.395 78.215 2.565 ;
      RECT 76.845 5.84 77.185 6.19 ;
      RECT 76.93 2.705 77.1 6.19 ;
      RECT 76.855 2.705 77.195 3.055 ;
      RECT 66.315 2.955 66.595 3.325 ;
      RECT 66.325 1.29 66.495 3.325 ;
      RECT 76.365 1.29 76.535 1.815 ;
      RECT 76.275 1.46 76.615 1.81 ;
      RECT 66.325 1.29 76.535 1.46 ;
      RECT 72.995 2.395 73.275 2.765 ;
      RECT 71.925 2.42 72.185 2.74 ;
      RECT 74.475 2.23 74.755 2.6 ;
      RECT 75.085 2.14 75.345 2.46 ;
      RECT 71.985 1.58 72.125 2.74 ;
      RECT 73.065 1.58 73.205 2.765 ;
      RECT 74.185 2.23 75.345 2.37 ;
      RECT 74.185 1.58 74.325 2.37 ;
      RECT 71.985 1.58 74.325 1.72 ;
      RECT 72.015 3.72 74.19 3.885 ;
      RECT 74.045 2.6 74.19 3.885 ;
      RECT 70.935 3.515 71.215 3.885 ;
      RECT 70.935 3.63 72.155 3.77 ;
      RECT 73.765 2.6 74.19 2.74 ;
      RECT 73.765 2.42 74.025 2.74 ;
      RECT 67.105 4 70.765 4.14 ;
      RECT 70.625 3.185 70.765 4.14 ;
      RECT 67.105 3.07 67.245 4.14 ;
      RECT 73.645 3.26 73.905 3.58 ;
      RECT 70.625 3.185 73.155 3.325 ;
      RECT 72.875 2.955 73.155 3.325 ;
      RECT 67.105 3.07 67.555 3.325 ;
      RECT 67.275 2.955 67.555 3.325 ;
      RECT 73.645 3.07 73.845 3.58 ;
      RECT 72.875 3.07 73.845 3.21 ;
      RECT 73.445 1.86 73.585 3.21 ;
      RECT 73.385 1.86 73.645 2.18 ;
      RECT 67.285 2.42 67.545 2.74 ;
      RECT 67.285 2.51 68.325 2.65 ;
      RECT 68.185 1.72 68.325 2.65 ;
      RECT 70.945 1.86 71.205 2.18 ;
      RECT 68.185 1.72 71.145 1.86 ;
      RECT 70.325 2.7 70.585 3.02 ;
      RECT 70.325 2.7 70.645 2.93 ;
      RECT 70.435 2.395 70.715 2.765 ;
      RECT 70.025 3.26 70.345 3.58 ;
      RECT 70.025 2.14 70.165 3.58 ;
      RECT 69.965 2.14 70.225 2.46 ;
      RECT 67.525 3.54 67.785 3.86 ;
      RECT 67.525 3.63 69.205 3.77 ;
      RECT 69.065 3.35 69.205 3.77 ;
      RECT 69.065 3.35 69.505 3.58 ;
      RECT 69.245 3.26 69.505 3.58 ;
      RECT 68.565 2.42 68.965 2.93 ;
      RECT 68.755 2.395 69.035 2.765 ;
      RECT 68.505 2.42 69.035 2.74 ;
      RECT 61.57 6.28 61.89 6.605 ;
      RECT 61.6 5.695 61.77 6.605 ;
      RECT 61.6 5.695 61.775 6.045 ;
      RECT 61.6 5.695 62.575 5.87 ;
      RECT 62.4 1.965 62.575 5.87 ;
      RECT 58.63 2.955 58.91 3.325 ;
      RECT 58.63 3.01 59.52 3.175 ;
      RECT 59.355 2.025 59.52 3.175 ;
      RECT 58.64 2.7 58.9 3.325 ;
      RECT 62.345 1.965 62.695 2.315 ;
      RECT 59.355 2.04 62.695 2.195 ;
      RECT 60.3 2.025 62.695 2.195 ;
      RECT 59.355 2.025 59.935 2.195 ;
      RECT 60.585 0.73 60.77 2.195 ;
      RECT 48.41 1.09 48.75 1.44 ;
      RECT 48.41 1.12 49.22 1.305 ;
      RECT 49.035 0.73 49.22 1.305 ;
      RECT 49.035 0.73 60.77 0.915 ;
      RECT 62.37 6.655 62.695 6.98 ;
      RECT 61.255 6.745 62.695 6.915 ;
      RECT 61.255 2.395 61.415 6.915 ;
      RECT 61.57 2.365 61.89 2.685 ;
      RECT 61.255 2.395 61.89 2.565 ;
      RECT 60.52 5.84 60.86 6.19 ;
      RECT 60.605 2.705 60.775 6.19 ;
      RECT 60.53 2.705 60.87 3.055 ;
      RECT 49.99 2.955 50.27 3.325 ;
      RECT 50 1.29 50.17 3.325 ;
      RECT 60.04 1.29 60.21 1.815 ;
      RECT 59.95 1.46 60.29 1.81 ;
      RECT 50 1.29 60.21 1.46 ;
      RECT 56.67 2.395 56.95 2.765 ;
      RECT 55.6 2.42 55.86 2.74 ;
      RECT 58.15 2.23 58.43 2.6 ;
      RECT 58.76 2.14 59.02 2.46 ;
      RECT 55.66 1.58 55.8 2.74 ;
      RECT 56.74 1.58 56.88 2.765 ;
      RECT 57.86 2.23 59.02 2.37 ;
      RECT 57.86 1.58 58 2.37 ;
      RECT 55.66 1.58 58 1.72 ;
      RECT 55.69 3.72 57.865 3.885 ;
      RECT 57.72 2.6 57.865 3.885 ;
      RECT 54.61 3.515 54.89 3.885 ;
      RECT 54.61 3.63 55.83 3.77 ;
      RECT 57.44 2.6 57.865 2.74 ;
      RECT 57.44 2.42 57.7 2.74 ;
      RECT 50.78 4 54.44 4.14 ;
      RECT 54.3 3.185 54.44 4.14 ;
      RECT 50.78 3.07 50.92 4.14 ;
      RECT 57.32 3.26 57.58 3.58 ;
      RECT 54.3 3.185 56.83 3.325 ;
      RECT 56.55 2.955 56.83 3.325 ;
      RECT 50.78 3.07 51.23 3.325 ;
      RECT 50.95 2.955 51.23 3.325 ;
      RECT 57.32 3.07 57.52 3.58 ;
      RECT 56.55 3.07 57.52 3.21 ;
      RECT 57.12 1.86 57.26 3.21 ;
      RECT 57.06 1.86 57.32 2.18 ;
      RECT 50.96 2.42 51.22 2.74 ;
      RECT 50.96 2.51 52 2.65 ;
      RECT 51.86 1.72 52 2.65 ;
      RECT 54.62 1.86 54.88 2.18 ;
      RECT 51.86 1.72 54.82 1.86 ;
      RECT 54 2.7 54.26 3.02 ;
      RECT 54 2.7 54.32 2.93 ;
      RECT 54.11 2.395 54.39 2.765 ;
      RECT 53.7 3.26 54.02 3.58 ;
      RECT 53.7 2.14 53.84 3.58 ;
      RECT 53.64 2.14 53.9 2.46 ;
      RECT 51.2 3.54 51.46 3.86 ;
      RECT 51.2 3.63 52.88 3.77 ;
      RECT 52.74 3.35 52.88 3.77 ;
      RECT 52.74 3.35 53.18 3.58 ;
      RECT 52.92 3.26 53.18 3.58 ;
      RECT 52.24 2.42 52.64 2.93 ;
      RECT 52.43 2.395 52.71 2.765 ;
      RECT 52.18 2.42 52.71 2.74 ;
      RECT 45.25 6.28 45.57 6.605 ;
      RECT 45.28 5.695 45.45 6.605 ;
      RECT 45.28 5.695 45.455 6.045 ;
      RECT 45.28 5.695 46.255 5.87 ;
      RECT 46.08 1.965 46.255 5.87 ;
      RECT 42.31 2.955 42.59 3.325 ;
      RECT 42.31 3.01 43.2 3.175 ;
      RECT 43.035 2.025 43.2 3.175 ;
      RECT 42.32 2.7 42.58 3.325 ;
      RECT 46.025 1.965 46.375 2.315 ;
      RECT 43.035 2.04 46.375 2.195 ;
      RECT 43.98 2.025 46.375 2.195 ;
      RECT 43.035 2.025 43.615 2.195 ;
      RECT 44.26 0.93 44.445 2.195 ;
      RECT 32.09 1.1 32.43 1.45 ;
      RECT 32.09 1.13 32.9 1.315 ;
      RECT 32.715 0.93 32.9 1.315 ;
      RECT 32.715 0.93 44.445 1.115 ;
      RECT 46.05 6.655 46.375 6.98 ;
      RECT 44.935 6.745 46.375 6.915 ;
      RECT 44.935 2.395 45.095 6.915 ;
      RECT 45.25 2.365 45.57 2.685 ;
      RECT 44.935 2.395 45.57 2.565 ;
      RECT 44.2 5.84 44.54 6.19 ;
      RECT 44.285 2.705 44.455 6.19 ;
      RECT 44.21 2.705 44.55 3.055 ;
      RECT 33.67 2.955 33.95 3.325 ;
      RECT 33.68 1.29 33.85 3.325 ;
      RECT 43.72 1.29 43.89 1.815 ;
      RECT 43.63 1.46 43.97 1.81 ;
      RECT 33.68 1.29 43.89 1.46 ;
      RECT 40.35 2.395 40.63 2.765 ;
      RECT 39.28 2.42 39.54 2.74 ;
      RECT 41.83 2.23 42.11 2.6 ;
      RECT 42.44 2.14 42.7 2.46 ;
      RECT 39.34 1.58 39.48 2.74 ;
      RECT 40.42 1.58 40.56 2.765 ;
      RECT 41.54 2.23 42.7 2.37 ;
      RECT 41.54 1.58 41.68 2.37 ;
      RECT 39.34 1.58 41.68 1.72 ;
      RECT 39.37 3.72 41.545 3.885 ;
      RECT 41.4 2.6 41.545 3.885 ;
      RECT 38.29 3.515 38.57 3.885 ;
      RECT 38.29 3.63 39.51 3.77 ;
      RECT 41.12 2.6 41.545 2.74 ;
      RECT 41.12 2.42 41.38 2.74 ;
      RECT 34.46 4 38.12 4.14 ;
      RECT 37.98 3.185 38.12 4.14 ;
      RECT 34.46 3.07 34.6 4.14 ;
      RECT 41 3.26 41.26 3.58 ;
      RECT 37.98 3.185 40.51 3.325 ;
      RECT 40.23 2.955 40.51 3.325 ;
      RECT 34.46 3.07 34.91 3.325 ;
      RECT 34.63 2.955 34.91 3.325 ;
      RECT 41 3.07 41.2 3.58 ;
      RECT 40.23 3.07 41.2 3.21 ;
      RECT 40.8 1.86 40.94 3.21 ;
      RECT 40.74 1.86 41 2.18 ;
      RECT 34.64 2.42 34.9 2.74 ;
      RECT 34.64 2.51 35.68 2.65 ;
      RECT 35.54 1.72 35.68 2.65 ;
      RECT 38.3 1.86 38.56 2.18 ;
      RECT 35.54 1.72 38.5 1.86 ;
      RECT 37.68 2.7 37.94 3.02 ;
      RECT 37.68 2.7 38 2.93 ;
      RECT 37.79 2.395 38.07 2.765 ;
      RECT 37.38 3.26 37.7 3.58 ;
      RECT 37.38 2.14 37.52 3.58 ;
      RECT 37.32 2.14 37.58 2.46 ;
      RECT 34.88 3.54 35.14 3.86 ;
      RECT 34.88 3.63 36.56 3.77 ;
      RECT 36.42 3.35 36.56 3.77 ;
      RECT 36.42 3.35 36.86 3.58 ;
      RECT 36.6 3.26 36.86 3.58 ;
      RECT 35.92 2.42 36.32 2.93 ;
      RECT 36.11 2.395 36.39 2.765 ;
      RECT 35.86 2.42 36.39 2.74 ;
      RECT 28.925 6.28 29.245 6.605 ;
      RECT 28.955 5.695 29.125 6.605 ;
      RECT 28.955 5.695 29.13 6.045 ;
      RECT 28.955 5.695 29.93 5.87 ;
      RECT 29.755 1.965 29.93 5.87 ;
      RECT 25.985 2.955 26.265 3.325 ;
      RECT 25.985 3.01 26.875 3.175 ;
      RECT 26.71 2.025 26.875 3.175 ;
      RECT 25.995 2.7 26.255 3.325 ;
      RECT 29.7 1.965 30.05 2.315 ;
      RECT 26.71 2.04 30.05 2.195 ;
      RECT 27.655 2.025 30.05 2.195 ;
      RECT 26.71 2.025 27.29 2.195 ;
      RECT 27.935 0.815 28.12 2.195 ;
      RECT 15.77 1.1 16.11 1.45 ;
      RECT 15.77 1.13 16.58 1.315 ;
      RECT 16.395 0.815 16.58 1.315 ;
      RECT 16.395 0.815 28.12 1 ;
      RECT 29.725 6.655 30.05 6.98 ;
      RECT 28.61 6.745 30.05 6.915 ;
      RECT 28.61 2.395 28.77 6.915 ;
      RECT 28.925 2.365 29.245 2.685 ;
      RECT 28.61 2.395 29.245 2.565 ;
      RECT 27.875 5.84 28.215 6.19 ;
      RECT 27.96 2.705 28.13 6.19 ;
      RECT 27.885 2.705 28.225 3.055 ;
      RECT 17.345 2.955 17.625 3.325 ;
      RECT 17.355 1.29 17.525 3.325 ;
      RECT 27.395 1.29 27.565 1.815 ;
      RECT 27.305 1.46 27.645 1.81 ;
      RECT 17.355 1.29 27.565 1.46 ;
      RECT 24.025 2.395 24.305 2.765 ;
      RECT 22.955 2.42 23.215 2.74 ;
      RECT 25.505 2.23 25.785 2.6 ;
      RECT 26.115 2.14 26.375 2.46 ;
      RECT 23.015 1.58 23.155 2.74 ;
      RECT 24.095 1.58 24.235 2.765 ;
      RECT 25.215 2.23 26.375 2.37 ;
      RECT 25.215 1.58 25.355 2.37 ;
      RECT 23.015 1.58 25.355 1.72 ;
      RECT 23.045 3.72 25.22 3.885 ;
      RECT 25.075 2.6 25.22 3.885 ;
      RECT 21.965 3.515 22.245 3.885 ;
      RECT 21.965 3.63 23.185 3.77 ;
      RECT 24.795 2.6 25.22 2.74 ;
      RECT 24.795 2.42 25.055 2.74 ;
      RECT 18.135 4 21.795 4.14 ;
      RECT 21.655 3.185 21.795 4.14 ;
      RECT 18.135 3.07 18.275 4.14 ;
      RECT 24.675 3.26 24.935 3.58 ;
      RECT 21.655 3.185 24.185 3.325 ;
      RECT 23.905 2.955 24.185 3.325 ;
      RECT 18.135 3.07 18.585 3.325 ;
      RECT 18.305 2.955 18.585 3.325 ;
      RECT 24.675 3.07 24.875 3.58 ;
      RECT 23.905 3.07 24.875 3.21 ;
      RECT 24.475 1.86 24.615 3.21 ;
      RECT 24.415 1.86 24.675 2.18 ;
      RECT 18.315 2.42 18.575 2.74 ;
      RECT 18.315 2.51 19.355 2.65 ;
      RECT 19.215 1.72 19.355 2.65 ;
      RECT 21.975 1.86 22.235 2.18 ;
      RECT 19.215 1.72 22.175 1.86 ;
      RECT 21.355 2.7 21.615 3.02 ;
      RECT 21.355 2.7 21.675 2.93 ;
      RECT 21.465 2.395 21.745 2.765 ;
      RECT 21.055 3.26 21.375 3.58 ;
      RECT 21.055 2.14 21.195 3.58 ;
      RECT 20.995 2.14 21.255 2.46 ;
      RECT 18.555 3.54 18.815 3.86 ;
      RECT 18.555 3.63 20.235 3.77 ;
      RECT 20.095 3.35 20.235 3.77 ;
      RECT 20.095 3.35 20.535 3.58 ;
      RECT 20.275 3.26 20.535 3.58 ;
      RECT 19.595 2.42 19.995 2.93 ;
      RECT 19.785 2.395 20.065 2.765 ;
      RECT 19.535 2.42 20.065 2.74 ;
      RECT 13.405 6.655 13.73 6.98 ;
      RECT 12.29 6.745 13.73 6.915 ;
      RECT 12.29 2.395 12.45 6.915 ;
      RECT 12.605 2.365 12.925 2.685 ;
      RECT 12.29 2.395 12.925 2.565 ;
      RECT 11.555 5.84 11.895 6.19 ;
      RECT 11.64 2.705 11.81 6.19 ;
      RECT 11.565 2.705 11.905 3.055 ;
      RECT 1.025 2.955 1.305 3.325 ;
      RECT 1.035 1.29 1.205 3.325 ;
      RECT 11.075 1.29 11.245 1.815 ;
      RECT 10.985 1.46 11.325 1.81 ;
      RECT 1.035 1.29 11.245 1.46 ;
      RECT 7.705 2.395 7.985 2.765 ;
      RECT 6.635 2.42 6.895 2.74 ;
      RECT 9.185 2.23 9.465 2.6 ;
      RECT 9.795 2.14 10.055 2.46 ;
      RECT 6.695 1.58 6.835 2.74 ;
      RECT 7.775 1.58 7.915 2.765 ;
      RECT 8.895 2.23 10.055 2.37 ;
      RECT 8.895 1.58 9.035 2.37 ;
      RECT 6.695 1.58 9.035 1.72 ;
      RECT 6.725 3.72 8.9 3.885 ;
      RECT 8.755 2.6 8.9 3.885 ;
      RECT 5.645 3.515 5.925 3.885 ;
      RECT 5.645 3.63 6.865 3.77 ;
      RECT 8.475 2.6 8.9 2.74 ;
      RECT 8.475 2.42 8.735 2.74 ;
      RECT 1.815 4 5.475 4.14 ;
      RECT 5.335 3.185 5.475 4.14 ;
      RECT 1.815 3.07 1.955 4.14 ;
      RECT 8.355 3.26 8.615 3.58 ;
      RECT 5.335 3.185 7.865 3.325 ;
      RECT 7.585 2.955 7.865 3.325 ;
      RECT 1.815 3.07 2.265 3.325 ;
      RECT 1.985 2.955 2.265 3.325 ;
      RECT 8.355 3.07 8.555 3.58 ;
      RECT 7.585 3.07 8.555 3.21 ;
      RECT 8.155 1.86 8.295 3.21 ;
      RECT 8.095 1.86 8.355 2.18 ;
      RECT 1.995 2.42 2.255 2.74 ;
      RECT 1.995 2.51 3.035 2.65 ;
      RECT 2.895 1.72 3.035 2.65 ;
      RECT 5.655 1.86 5.915 2.18 ;
      RECT 2.895 1.72 5.855 1.86 ;
      RECT 5.035 2.7 5.295 3.02 ;
      RECT 5.035 2.7 5.355 2.93 ;
      RECT 5.145 2.395 5.425 2.765 ;
      RECT 4.735 3.26 5.055 3.58 ;
      RECT 4.735 2.14 4.875 3.58 ;
      RECT 4.675 2.14 4.935 2.46 ;
      RECT 2.235 3.54 2.495 3.86 ;
      RECT 2.235 3.63 3.915 3.77 ;
      RECT 3.775 3.35 3.915 3.77 ;
      RECT 3.775 3.35 4.215 3.58 ;
      RECT 3.955 3.26 4.215 3.58 ;
      RECT 3.275 2.42 3.675 2.93 ;
      RECT 3.465 2.395 3.745 2.765 ;
      RECT 3.215 2.42 3.745 2.74 ;
      RECT 71.315 2.395 71.595 2.765 ;
      RECT 69.475 2.395 69.755 2.765 ;
      RECT 67.755 1.835 68.035 2.205 ;
      RECT 54.99 2.395 55.27 2.765 ;
      RECT 53.15 2.395 53.43 2.765 ;
      RECT 51.43 1.835 51.71 2.205 ;
      RECT 38.67 2.395 38.95 2.765 ;
      RECT 36.83 2.395 37.11 2.765 ;
      RECT 35.11 1.835 35.39 2.205 ;
      RECT 22.345 2.395 22.625 2.765 ;
      RECT 20.505 2.395 20.785 2.765 ;
      RECT 18.785 1.835 19.065 2.205 ;
      RECT 6.025 2.395 6.305 2.765 ;
      RECT 4.185 2.395 4.465 2.765 ;
      RECT 2.465 1.835 2.745 2.205 ;
    LAYER via1 ;
      RECT 81.155 1.195 81.305 1.345 ;
      RECT 78.785 6.74 78.935 6.89 ;
      RECT 78.77 2.065 78.92 2.215 ;
      RECT 77.98 2.45 78.13 2.6 ;
      RECT 77.98 6.37 78.13 6.52 ;
      RECT 76.955 2.805 77.105 2.955 ;
      RECT 76.945 5.94 77.095 6.09 ;
      RECT 76.375 1.56 76.525 1.71 ;
      RECT 75.14 2.225 75.29 2.375 ;
      RECT 75.02 2.785 75.17 2.935 ;
      RECT 73.82 2.505 73.97 2.655 ;
      RECT 73.7 3.345 73.85 3.495 ;
      RECT 73.44 1.945 73.59 2.095 ;
      RECT 71.98 2.505 72.13 2.655 ;
      RECT 71.38 2.505 71.53 2.655 ;
      RECT 71 1.945 71.15 2.095 ;
      RECT 70.38 2.785 70.53 2.935 ;
      RECT 70.14 3.345 70.29 3.495 ;
      RECT 70.02 2.225 70.17 2.375 ;
      RECT 69.54 2.505 69.69 2.655 ;
      RECT 69.3 3.345 69.45 3.495 ;
      RECT 68.56 2.505 68.71 2.655 ;
      RECT 67.82 1.945 67.97 2.095 ;
      RECT 67.58 3.625 67.73 3.775 ;
      RECT 67.34 2.505 67.49 2.655 ;
      RECT 67.34 3.065 67.49 3.215 ;
      RECT 66.38 3.065 66.53 3.215 ;
      RECT 64.83 1.195 64.98 1.345 ;
      RECT 62.46 6.74 62.61 6.89 ;
      RECT 62.445 2.065 62.595 2.215 ;
      RECT 61.655 2.45 61.805 2.6 ;
      RECT 61.655 6.37 61.805 6.52 ;
      RECT 60.63 2.805 60.78 2.955 ;
      RECT 60.62 5.94 60.77 6.09 ;
      RECT 60.05 1.56 60.2 1.71 ;
      RECT 58.815 2.225 58.965 2.375 ;
      RECT 58.695 2.785 58.845 2.935 ;
      RECT 57.495 2.505 57.645 2.655 ;
      RECT 57.375 3.345 57.525 3.495 ;
      RECT 57.115 1.945 57.265 2.095 ;
      RECT 55.655 2.505 55.805 2.655 ;
      RECT 55.055 2.505 55.205 2.655 ;
      RECT 54.675 1.945 54.825 2.095 ;
      RECT 54.055 2.785 54.205 2.935 ;
      RECT 53.815 3.345 53.965 3.495 ;
      RECT 53.695 2.225 53.845 2.375 ;
      RECT 53.215 2.505 53.365 2.655 ;
      RECT 52.975 3.345 53.125 3.495 ;
      RECT 52.235 2.505 52.385 2.655 ;
      RECT 51.495 1.945 51.645 2.095 ;
      RECT 51.255 3.625 51.405 3.775 ;
      RECT 51.015 2.505 51.165 2.655 ;
      RECT 51.015 3.065 51.165 3.215 ;
      RECT 50.055 3.065 50.205 3.215 ;
      RECT 48.51 1.19 48.66 1.34 ;
      RECT 46.14 6.74 46.29 6.89 ;
      RECT 46.125 2.065 46.275 2.215 ;
      RECT 45.335 2.45 45.485 2.6 ;
      RECT 45.335 6.37 45.485 6.52 ;
      RECT 44.31 2.805 44.46 2.955 ;
      RECT 44.3 5.94 44.45 6.09 ;
      RECT 43.73 1.56 43.88 1.71 ;
      RECT 42.495 2.225 42.645 2.375 ;
      RECT 42.375 2.785 42.525 2.935 ;
      RECT 41.175 2.505 41.325 2.655 ;
      RECT 41.055 3.345 41.205 3.495 ;
      RECT 40.795 1.945 40.945 2.095 ;
      RECT 39.335 2.505 39.485 2.655 ;
      RECT 38.735 2.505 38.885 2.655 ;
      RECT 38.355 1.945 38.505 2.095 ;
      RECT 37.735 2.785 37.885 2.935 ;
      RECT 37.495 3.345 37.645 3.495 ;
      RECT 37.375 2.225 37.525 2.375 ;
      RECT 36.895 2.505 37.045 2.655 ;
      RECT 36.655 3.345 36.805 3.495 ;
      RECT 35.915 2.505 36.065 2.655 ;
      RECT 35.175 1.945 35.325 2.095 ;
      RECT 34.935 3.625 35.085 3.775 ;
      RECT 34.695 2.505 34.845 2.655 ;
      RECT 34.695 3.065 34.845 3.215 ;
      RECT 33.735 3.065 33.885 3.215 ;
      RECT 32.19 1.2 32.34 1.35 ;
      RECT 29.815 6.74 29.965 6.89 ;
      RECT 29.8 2.065 29.95 2.215 ;
      RECT 29.01 2.45 29.16 2.6 ;
      RECT 29.01 6.37 29.16 6.52 ;
      RECT 27.985 2.805 28.135 2.955 ;
      RECT 27.975 5.94 28.125 6.09 ;
      RECT 27.405 1.56 27.555 1.71 ;
      RECT 26.17 2.225 26.32 2.375 ;
      RECT 26.05 2.785 26.2 2.935 ;
      RECT 24.85 2.505 25 2.655 ;
      RECT 24.73 3.345 24.88 3.495 ;
      RECT 24.47 1.945 24.62 2.095 ;
      RECT 23.01 2.505 23.16 2.655 ;
      RECT 22.41 2.505 22.56 2.655 ;
      RECT 22.03 1.945 22.18 2.095 ;
      RECT 21.41 2.785 21.56 2.935 ;
      RECT 21.17 3.345 21.32 3.495 ;
      RECT 21.05 2.225 21.2 2.375 ;
      RECT 20.57 2.505 20.72 2.655 ;
      RECT 20.33 3.345 20.48 3.495 ;
      RECT 19.59 2.505 19.74 2.655 ;
      RECT 18.85 1.945 19 2.095 ;
      RECT 18.61 3.625 18.76 3.775 ;
      RECT 18.37 2.505 18.52 2.655 ;
      RECT 18.37 3.065 18.52 3.215 ;
      RECT 17.41 3.065 17.56 3.215 ;
      RECT 15.87 1.2 16.02 1.35 ;
      RECT 13.495 6.74 13.645 6.89 ;
      RECT 13.48 2.065 13.63 2.215 ;
      RECT 12.69 2.45 12.84 2.6 ;
      RECT 12.69 6.37 12.84 6.52 ;
      RECT 11.665 2.805 11.815 2.955 ;
      RECT 11.655 5.94 11.805 6.09 ;
      RECT 11.085 1.56 11.235 1.71 ;
      RECT 9.85 2.225 10 2.375 ;
      RECT 9.73 2.785 9.88 2.935 ;
      RECT 8.53 2.505 8.68 2.655 ;
      RECT 8.41 3.345 8.56 3.495 ;
      RECT 8.15 1.945 8.3 2.095 ;
      RECT 6.69 2.505 6.84 2.655 ;
      RECT 6.09 2.505 6.24 2.655 ;
      RECT 5.71 1.945 5.86 2.095 ;
      RECT 5.09 2.785 5.24 2.935 ;
      RECT 4.85 3.345 5 3.495 ;
      RECT 4.73 2.225 4.88 2.375 ;
      RECT 4.25 2.505 4.4 2.655 ;
      RECT 4.01 3.345 4.16 3.495 ;
      RECT 3.27 2.505 3.42 2.655 ;
      RECT 2.53 1.945 2.68 2.095 ;
      RECT 2.29 3.625 2.44 3.775 ;
      RECT 2.05 2.505 2.2 2.655 ;
      RECT 2.05 3.065 2.2 3.215 ;
      RECT 1.09 3.065 1.24 3.215 ;
    LAYER met1 ;
      RECT 66.04 0 75.7 1.74 ;
      RECT 49.715 0 59.375 1.74 ;
      RECT 33.395 0 43.055 1.74 ;
      RECT 17.07 0 26.73 1.74 ;
      RECT 0.75 0 10.41 1.74 ;
      RECT 66.04 0 75.855 1.585 ;
      RECT 49.715 0 59.53 1.585 ;
      RECT 33.395 0 43.21 1.585 ;
      RECT 17.07 0 26.885 1.585 ;
      RECT 0.75 0 10.565 1.585 ;
      RECT 0.005 0 81.625 0.305 ;
      RECT 0.005 4.135 81.625 4.745 ;
      RECT 66.04 3.98 75.7 4.745 ;
      RECT 49.715 3.98 59.375 4.745 ;
      RECT 33.395 3.98 43.055 4.745 ;
      RECT 17.07 3.98 26.73 4.745 ;
      RECT 0.75 3.98 10.41 4.745 ;
      RECT 81.025 2.365 81.315 2.595 ;
      RECT 81.085 0.885 81.255 2.595 ;
      RECT 81.055 1.095 81.395 1.445 ;
      RECT 81.025 0.885 81.315 1.115 ;
      RECT 81.025 7.765 81.315 7.995 ;
      RECT 81.085 6.285 81.255 7.995 ;
      RECT 81.025 6.285 81.315 6.515 ;
      RECT 80.615 2.735 80.945 2.965 ;
      RECT 80.615 2.765 81.115 2.935 ;
      RECT 80.615 2.395 80.805 2.965 ;
      RECT 80.035 2.365 80.325 2.595 ;
      RECT 80.035 2.395 80.805 2.565 ;
      RECT 80.095 0.885 80.265 2.595 ;
      RECT 80.035 0.885 80.325 1.115 ;
      RECT 80.035 7.765 80.325 7.995 ;
      RECT 80.095 6.285 80.265 7.995 ;
      RECT 80.035 6.285 80.325 6.515 ;
      RECT 80.035 6.325 80.885 6.485 ;
      RECT 80.715 5.915 80.885 6.485 ;
      RECT 80.035 6.32 80.425 6.485 ;
      RECT 80.655 5.915 80.945 6.145 ;
      RECT 80.655 5.945 81.115 6.115 ;
      RECT 79.665 2.735 79.955 2.965 ;
      RECT 79.665 2.765 80.125 2.935 ;
      RECT 79.725 1.655 79.89 2.965 ;
      RECT 78.24 1.625 78.53 1.855 ;
      RECT 78.24 1.655 79.89 1.825 ;
      RECT 78.3 0.885 78.47 1.855 ;
      RECT 78.24 0.885 78.53 1.115 ;
      RECT 78.24 7.765 78.53 7.995 ;
      RECT 78.3 7.025 78.47 7.995 ;
      RECT 78.3 7.12 79.89 7.29 ;
      RECT 79.72 5.915 79.89 7.29 ;
      RECT 78.24 7.025 78.53 7.255 ;
      RECT 79.665 5.915 79.955 6.145 ;
      RECT 79.665 5.945 80.125 6.115 ;
      RECT 78.67 1.965 79.02 2.315 ;
      RECT 78.5 2.025 79.02 2.195 ;
      RECT 78.695 6.655 79.02 6.98 ;
      RECT 78.67 6.655 79.02 6.885 ;
      RECT 78.5 6.685 79.02 6.855 ;
      RECT 77.895 2.365 78.215 2.685 ;
      RECT 77.865 2.365 78.215 2.595 ;
      RECT 76.365 2.395 78.215 2.565 ;
      RECT 76.365 1.46 76.535 2.565 ;
      RECT 76.275 1.46 76.615 1.81 ;
      RECT 77.895 6.28 78.215 6.605 ;
      RECT 77.865 6.285 78.215 6.515 ;
      RECT 77.695 6.315 78.215 6.485 ;
      RECT 76.855 2.705 77.195 3.055 ;
      RECT 76.855 2.765 77.33 2.935 ;
      RECT 76.845 5.84 77.185 6.19 ;
      RECT 76.845 5.945 77.33 6.115 ;
      RECT 74.35 2.465 74.64 2.695 ;
      RECT 74.35 2.465 74.805 2.65 ;
      RECT 74.665 2.37 75.285 2.51 ;
      RECT 75.055 2.17 75.375 2.43 ;
      RECT 73.445 2.93 75.045 3.07 ;
      RECT 73.445 2.93 75.21 3.055 ;
      RECT 74.935 2.73 75.255 2.99 ;
      RECT 74.89 2.745 75.36 2.975 ;
      RECT 73.11 2.79 73.585 2.975 ;
      RECT 73.11 2.745 73.4 2.975 ;
      RECT 74.89 2.735 75.255 2.99 ;
      RECT 73.735 2.45 74.055 2.71 ;
      RECT 73.735 2.45 74.2 2.695 ;
      RECT 74.06 2.07 74.2 2.695 ;
      RECT 74.06 2.07 74.325 2.21 ;
      RECT 74.59 1.905 74.88 2.135 ;
      RECT 74.185 1.95 74.88 2.09 ;
      RECT 73.63 3.29 73.92 3.815 ;
      RECT 73.615 3.29 73.935 3.55 ;
      RECT 73.355 1.89 73.675 2.15 ;
      RECT 73.355 1.905 73.92 2.135 ;
      RECT 72.63 3.585 72.92 3.815 ;
      RECT 72.825 2.23 72.965 3.77 ;
      RECT 72.87 2.185 73.16 2.415 ;
      RECT 72.465 2.23 73.16 2.37 ;
      RECT 72.465 2.07 72.605 2.37 ;
      RECT 71.005 2.07 72.605 2.21 ;
      RECT 70.915 1.89 71.235 2.15 ;
      RECT 70.915 1.905 71.48 2.15 ;
      RECT 70.025 2.93 72.605 3.07 ;
      RECT 72.39 2.745 72.68 2.975 ;
      RECT 69.95 2.745 70.615 2.975 ;
      RECT 70.295 2.73 70.615 3.07 ;
      RECT 71.295 2.45 71.615 2.71 ;
      RECT 71.295 2.465 71.72 2.695 ;
      RECT 69.935 2.17 70.255 2.43 ;
      RECT 70.43 2.185 70.72 2.415 ;
      RECT 69.935 2.23 70.72 2.37 ;
      RECT 70.055 3.29 70.375 3.55 ;
      RECT 69.215 3.29 69.535 3.55 ;
      RECT 70.055 3.305 70.48 3.535 ;
      RECT 69.215 3.35 70.48 3.49 ;
      RECT 68.75 3.025 69.04 3.255 ;
      RECT 68.825 1.95 68.965 3.255 ;
      RECT 68.475 2.45 68.965 2.71 ;
      RECT 68.23 2.465 68.965 2.695 ;
      RECT 69.23 1.905 69.52 2.135 ;
      RECT 68.825 1.95 69.52 2.09 ;
      RECT 67.99 3.305 68.28 3.535 ;
      RECT 67.99 3.305 68.445 3.49 ;
      RECT 68.305 2.93 68.445 3.49 ;
      RECT 67.945 2.93 68.445 3.07 ;
      RECT 67.945 1.95 68.085 3.07 ;
      RECT 67.735 1.89 68.055 2.15 ;
      RECT 67.495 3.57 67.815 3.83 ;
      RECT 66.79 3.585 67.08 3.815 ;
      RECT 66.79 3.63 67.815 3.77 ;
      RECT 66.865 3.58 67.125 3.77 ;
      RECT 67.255 2.45 67.575 2.71 ;
      RECT 67.255 2.465 67.8 2.695 ;
      RECT 67.255 3.01 67.575 3.27 ;
      RECT 67.255 3.025 67.8 3.255 ;
      RECT 66.295 3.01 66.615 3.27 ;
      RECT 66.385 1.95 66.525 3.27 ;
      RECT 66.79 1.905 67.08 2.135 ;
      RECT 66.385 1.95 67.08 2.09 ;
      RECT 64.7 2.365 64.99 2.595 ;
      RECT 64.76 0.885 64.93 2.595 ;
      RECT 64.73 1.095 65.07 1.445 ;
      RECT 64.7 0.885 64.99 1.115 ;
      RECT 64.7 7.765 64.99 7.995 ;
      RECT 64.76 6.285 64.93 7.995 ;
      RECT 64.7 6.285 64.99 6.515 ;
      RECT 64.29 2.735 64.62 2.965 ;
      RECT 64.29 2.765 64.79 2.935 ;
      RECT 64.29 2.395 64.48 2.965 ;
      RECT 63.71 2.365 64 2.595 ;
      RECT 63.71 2.395 64.48 2.565 ;
      RECT 63.77 0.885 63.94 2.595 ;
      RECT 63.71 0.885 64 1.115 ;
      RECT 63.71 7.765 64 7.995 ;
      RECT 63.77 6.285 63.94 7.995 ;
      RECT 63.71 6.285 64 6.515 ;
      RECT 63.71 6.325 64.56 6.485 ;
      RECT 64.39 5.915 64.56 6.485 ;
      RECT 63.71 6.32 64.1 6.485 ;
      RECT 64.33 5.915 64.62 6.145 ;
      RECT 64.33 5.945 64.79 6.115 ;
      RECT 63.34 2.735 63.63 2.965 ;
      RECT 63.34 2.765 63.8 2.935 ;
      RECT 63.4 1.655 63.565 2.965 ;
      RECT 61.915 1.625 62.205 1.855 ;
      RECT 61.915 1.655 63.565 1.825 ;
      RECT 61.975 0.885 62.145 1.855 ;
      RECT 61.915 0.885 62.205 1.115 ;
      RECT 61.915 7.765 62.205 7.995 ;
      RECT 61.975 7.025 62.145 7.995 ;
      RECT 61.975 7.12 63.565 7.29 ;
      RECT 63.395 5.915 63.565 7.29 ;
      RECT 61.915 7.025 62.205 7.255 ;
      RECT 63.34 5.915 63.63 6.145 ;
      RECT 63.34 5.945 63.8 6.115 ;
      RECT 62.345 1.965 62.695 2.315 ;
      RECT 62.175 2.025 62.695 2.195 ;
      RECT 62.37 6.655 62.695 6.98 ;
      RECT 62.345 6.655 62.695 6.885 ;
      RECT 62.175 6.685 62.695 6.855 ;
      RECT 61.57 2.365 61.89 2.685 ;
      RECT 61.54 2.365 61.89 2.595 ;
      RECT 60.04 2.395 61.89 2.565 ;
      RECT 60.04 1.46 60.21 2.565 ;
      RECT 59.95 1.46 60.29 1.81 ;
      RECT 61.57 6.28 61.89 6.605 ;
      RECT 61.54 6.285 61.89 6.515 ;
      RECT 61.37 6.315 61.89 6.485 ;
      RECT 60.53 2.705 60.87 3.055 ;
      RECT 60.53 2.765 61.005 2.935 ;
      RECT 60.52 5.84 60.86 6.19 ;
      RECT 60.52 5.945 61.005 6.115 ;
      RECT 58.025 2.465 58.315 2.695 ;
      RECT 58.025 2.465 58.48 2.65 ;
      RECT 58.34 2.37 58.96 2.51 ;
      RECT 58.73 2.17 59.05 2.43 ;
      RECT 57.12 2.93 58.72 3.07 ;
      RECT 57.12 2.93 58.885 3.055 ;
      RECT 58.61 2.73 58.93 2.99 ;
      RECT 58.565 2.745 59.035 2.975 ;
      RECT 56.785 2.79 57.26 2.975 ;
      RECT 56.785 2.745 57.075 2.975 ;
      RECT 58.565 2.735 58.93 2.99 ;
      RECT 57.41 2.45 57.73 2.71 ;
      RECT 57.41 2.45 57.875 2.695 ;
      RECT 57.735 2.07 57.875 2.695 ;
      RECT 57.735 2.07 58 2.21 ;
      RECT 58.265 1.905 58.555 2.135 ;
      RECT 57.86 1.95 58.555 2.09 ;
      RECT 57.305 3.29 57.595 3.815 ;
      RECT 57.29 3.29 57.61 3.55 ;
      RECT 57.03 1.89 57.35 2.15 ;
      RECT 57.03 1.905 57.595 2.135 ;
      RECT 56.305 3.585 56.595 3.815 ;
      RECT 56.5 2.23 56.64 3.77 ;
      RECT 56.545 2.185 56.835 2.415 ;
      RECT 56.14 2.23 56.835 2.37 ;
      RECT 56.14 2.07 56.28 2.37 ;
      RECT 54.68 2.07 56.28 2.21 ;
      RECT 54.59 1.89 54.91 2.15 ;
      RECT 54.59 1.905 55.155 2.15 ;
      RECT 53.7 2.93 56.28 3.07 ;
      RECT 56.065 2.745 56.355 2.975 ;
      RECT 53.625 2.745 54.29 2.975 ;
      RECT 53.97 2.73 54.29 3.07 ;
      RECT 54.97 2.45 55.29 2.71 ;
      RECT 54.97 2.465 55.395 2.695 ;
      RECT 53.61 2.17 53.93 2.43 ;
      RECT 54.105 2.185 54.395 2.415 ;
      RECT 53.61 2.23 54.395 2.37 ;
      RECT 53.73 3.29 54.05 3.55 ;
      RECT 52.89 3.29 53.21 3.55 ;
      RECT 53.73 3.305 54.155 3.535 ;
      RECT 52.89 3.35 54.155 3.49 ;
      RECT 52.425 3.025 52.715 3.255 ;
      RECT 52.5 1.95 52.64 3.255 ;
      RECT 52.15 2.45 52.64 2.71 ;
      RECT 51.905 2.465 52.64 2.695 ;
      RECT 52.905 1.905 53.195 2.135 ;
      RECT 52.5 1.95 53.195 2.09 ;
      RECT 51.665 3.305 51.955 3.535 ;
      RECT 51.665 3.305 52.12 3.49 ;
      RECT 51.98 2.93 52.12 3.49 ;
      RECT 51.62 2.93 52.12 3.07 ;
      RECT 51.62 1.95 51.76 3.07 ;
      RECT 51.41 1.89 51.73 2.15 ;
      RECT 51.17 3.57 51.49 3.83 ;
      RECT 50.465 3.585 50.755 3.815 ;
      RECT 50.465 3.63 51.49 3.77 ;
      RECT 50.54 3.58 50.8 3.77 ;
      RECT 50.93 2.45 51.25 2.71 ;
      RECT 50.93 2.465 51.475 2.695 ;
      RECT 50.93 3.01 51.25 3.27 ;
      RECT 50.93 3.025 51.475 3.255 ;
      RECT 49.97 3.01 50.29 3.27 ;
      RECT 50.06 1.95 50.2 3.27 ;
      RECT 50.465 1.905 50.755 2.135 ;
      RECT 50.06 1.95 50.755 2.09 ;
      RECT 48.38 2.365 48.67 2.595 ;
      RECT 48.44 0.885 48.61 2.595 ;
      RECT 48.41 1.09 48.75 1.44 ;
      RECT 48.38 0.885 48.67 1.115 ;
      RECT 48.38 7.765 48.67 7.995 ;
      RECT 48.44 6.285 48.61 7.995 ;
      RECT 48.38 6.285 48.67 6.515 ;
      RECT 47.97 2.735 48.3 2.965 ;
      RECT 47.97 2.765 48.47 2.935 ;
      RECT 47.97 2.395 48.16 2.965 ;
      RECT 47.39 2.365 47.68 2.595 ;
      RECT 47.39 2.395 48.16 2.565 ;
      RECT 47.45 0.885 47.62 2.595 ;
      RECT 47.39 0.885 47.68 1.115 ;
      RECT 47.39 7.765 47.68 7.995 ;
      RECT 47.45 6.285 47.62 7.995 ;
      RECT 47.39 6.285 47.68 6.515 ;
      RECT 47.39 6.325 48.24 6.485 ;
      RECT 48.07 5.915 48.24 6.485 ;
      RECT 47.39 6.32 47.78 6.485 ;
      RECT 48.01 5.915 48.3 6.145 ;
      RECT 48.01 5.945 48.47 6.115 ;
      RECT 47.02 2.735 47.31 2.965 ;
      RECT 47.02 2.765 47.48 2.935 ;
      RECT 47.08 1.655 47.245 2.965 ;
      RECT 45.595 1.625 45.885 1.855 ;
      RECT 45.595 1.655 47.245 1.825 ;
      RECT 45.655 0.885 45.825 1.855 ;
      RECT 45.595 0.885 45.885 1.115 ;
      RECT 45.595 7.765 45.885 7.995 ;
      RECT 45.655 7.025 45.825 7.995 ;
      RECT 45.655 7.12 47.245 7.29 ;
      RECT 47.075 5.915 47.245 7.29 ;
      RECT 45.595 7.025 45.885 7.255 ;
      RECT 47.02 5.915 47.31 6.145 ;
      RECT 47.02 5.945 47.48 6.115 ;
      RECT 46.025 1.965 46.375 2.315 ;
      RECT 45.855 2.025 46.375 2.195 ;
      RECT 46.05 6.655 46.375 6.98 ;
      RECT 46.025 6.655 46.375 6.885 ;
      RECT 45.855 6.685 46.375 6.855 ;
      RECT 45.25 2.365 45.57 2.685 ;
      RECT 45.22 2.365 45.57 2.595 ;
      RECT 43.72 2.395 45.57 2.565 ;
      RECT 43.72 1.46 43.89 2.565 ;
      RECT 43.63 1.46 43.97 1.81 ;
      RECT 45.25 6.28 45.57 6.605 ;
      RECT 45.22 6.285 45.57 6.515 ;
      RECT 45.05 6.315 45.57 6.485 ;
      RECT 44.21 2.705 44.55 3.055 ;
      RECT 44.21 2.765 44.685 2.935 ;
      RECT 44.2 5.84 44.54 6.19 ;
      RECT 44.2 5.945 44.685 6.115 ;
      RECT 41.705 2.465 41.995 2.695 ;
      RECT 41.705 2.465 42.16 2.65 ;
      RECT 42.02 2.37 42.64 2.51 ;
      RECT 42.41 2.17 42.73 2.43 ;
      RECT 40.8 2.93 42.4 3.07 ;
      RECT 40.8 2.93 42.565 3.055 ;
      RECT 42.29 2.73 42.61 2.99 ;
      RECT 42.245 2.745 42.715 2.975 ;
      RECT 40.465 2.79 40.94 2.975 ;
      RECT 40.465 2.745 40.755 2.975 ;
      RECT 42.245 2.735 42.61 2.99 ;
      RECT 41.09 2.45 41.41 2.71 ;
      RECT 41.09 2.45 41.555 2.695 ;
      RECT 41.415 2.07 41.555 2.695 ;
      RECT 41.415 2.07 41.68 2.21 ;
      RECT 41.945 1.905 42.235 2.135 ;
      RECT 41.54 1.95 42.235 2.09 ;
      RECT 40.985 3.29 41.275 3.815 ;
      RECT 40.97 3.29 41.29 3.55 ;
      RECT 40.71 1.89 41.03 2.15 ;
      RECT 40.71 1.905 41.275 2.135 ;
      RECT 39.985 3.585 40.275 3.815 ;
      RECT 40.18 2.23 40.32 3.77 ;
      RECT 40.225 2.185 40.515 2.415 ;
      RECT 39.82 2.23 40.515 2.37 ;
      RECT 39.82 2.07 39.96 2.37 ;
      RECT 38.36 2.07 39.96 2.21 ;
      RECT 38.27 1.89 38.59 2.15 ;
      RECT 38.27 1.905 38.835 2.15 ;
      RECT 37.38 2.93 39.96 3.07 ;
      RECT 39.745 2.745 40.035 2.975 ;
      RECT 37.305 2.745 37.97 2.975 ;
      RECT 37.65 2.73 37.97 3.07 ;
      RECT 38.65 2.45 38.97 2.71 ;
      RECT 38.65 2.465 39.075 2.695 ;
      RECT 37.29 2.17 37.61 2.43 ;
      RECT 37.785 2.185 38.075 2.415 ;
      RECT 37.29 2.23 38.075 2.37 ;
      RECT 37.41 3.29 37.73 3.55 ;
      RECT 36.57 3.29 36.89 3.55 ;
      RECT 37.41 3.305 37.835 3.535 ;
      RECT 36.57 3.35 37.835 3.49 ;
      RECT 36.105 3.025 36.395 3.255 ;
      RECT 36.18 1.95 36.32 3.255 ;
      RECT 35.83 2.45 36.32 2.71 ;
      RECT 35.585 2.465 36.32 2.695 ;
      RECT 36.585 1.905 36.875 2.135 ;
      RECT 36.18 1.95 36.875 2.09 ;
      RECT 35.345 3.305 35.635 3.535 ;
      RECT 35.345 3.305 35.8 3.49 ;
      RECT 35.66 2.93 35.8 3.49 ;
      RECT 35.3 2.93 35.8 3.07 ;
      RECT 35.3 1.95 35.44 3.07 ;
      RECT 35.09 1.89 35.41 2.15 ;
      RECT 34.85 3.57 35.17 3.83 ;
      RECT 34.145 3.585 34.435 3.815 ;
      RECT 34.145 3.63 35.17 3.77 ;
      RECT 34.22 3.58 34.48 3.77 ;
      RECT 34.61 2.45 34.93 2.71 ;
      RECT 34.61 2.465 35.155 2.695 ;
      RECT 34.61 3.01 34.93 3.27 ;
      RECT 34.61 3.025 35.155 3.255 ;
      RECT 33.65 3.01 33.97 3.27 ;
      RECT 33.74 1.95 33.88 3.27 ;
      RECT 34.145 1.905 34.435 2.135 ;
      RECT 33.74 1.95 34.435 2.09 ;
      RECT 32.055 2.365 32.345 2.595 ;
      RECT 32.115 0.885 32.285 2.595 ;
      RECT 32.09 1.1 32.43 1.45 ;
      RECT 32.055 0.885 32.345 1.115 ;
      RECT 32.055 7.765 32.345 7.995 ;
      RECT 32.115 6.285 32.285 7.995 ;
      RECT 32.055 6.285 32.345 6.515 ;
      RECT 31.645 2.735 31.975 2.965 ;
      RECT 31.645 2.765 32.145 2.935 ;
      RECT 31.645 2.395 31.835 2.965 ;
      RECT 31.065 2.365 31.355 2.595 ;
      RECT 31.065 2.395 31.835 2.565 ;
      RECT 31.125 0.885 31.295 2.595 ;
      RECT 31.065 0.885 31.355 1.115 ;
      RECT 31.065 7.765 31.355 7.995 ;
      RECT 31.125 6.285 31.295 7.995 ;
      RECT 31.065 6.285 31.355 6.515 ;
      RECT 31.065 6.325 31.915 6.485 ;
      RECT 31.745 5.915 31.915 6.485 ;
      RECT 31.065 6.32 31.455 6.485 ;
      RECT 31.685 5.915 31.975 6.145 ;
      RECT 31.685 5.945 32.145 6.115 ;
      RECT 30.695 2.735 30.985 2.965 ;
      RECT 30.695 2.765 31.155 2.935 ;
      RECT 30.755 1.655 30.92 2.965 ;
      RECT 29.27 1.625 29.56 1.855 ;
      RECT 29.27 1.655 30.92 1.825 ;
      RECT 29.33 0.885 29.5 1.855 ;
      RECT 29.27 0.885 29.56 1.115 ;
      RECT 29.27 7.765 29.56 7.995 ;
      RECT 29.33 7.025 29.5 7.995 ;
      RECT 29.33 7.12 30.92 7.29 ;
      RECT 30.75 5.915 30.92 7.29 ;
      RECT 29.27 7.025 29.56 7.255 ;
      RECT 30.695 5.915 30.985 6.145 ;
      RECT 30.695 5.945 31.155 6.115 ;
      RECT 29.7 1.965 30.05 2.315 ;
      RECT 29.53 2.025 30.05 2.195 ;
      RECT 29.725 6.655 30.05 6.98 ;
      RECT 29.7 6.655 30.05 6.885 ;
      RECT 29.53 6.685 30.05 6.855 ;
      RECT 28.925 2.365 29.245 2.685 ;
      RECT 28.895 2.365 29.245 2.595 ;
      RECT 27.395 2.395 29.245 2.565 ;
      RECT 27.395 1.46 27.565 2.565 ;
      RECT 27.305 1.46 27.645 1.81 ;
      RECT 28.925 6.28 29.245 6.605 ;
      RECT 28.895 6.285 29.245 6.515 ;
      RECT 28.725 6.315 29.245 6.485 ;
      RECT 27.885 2.705 28.225 3.055 ;
      RECT 27.885 2.765 28.36 2.935 ;
      RECT 27.875 5.84 28.215 6.19 ;
      RECT 27.875 5.945 28.36 6.115 ;
      RECT 25.38 2.465 25.67 2.695 ;
      RECT 25.38 2.465 25.835 2.65 ;
      RECT 25.695 2.37 26.315 2.51 ;
      RECT 26.085 2.17 26.405 2.43 ;
      RECT 24.475 2.93 26.075 3.07 ;
      RECT 24.475 2.93 26.24 3.055 ;
      RECT 25.965 2.73 26.285 2.99 ;
      RECT 25.92 2.745 26.39 2.975 ;
      RECT 24.14 2.79 24.615 2.975 ;
      RECT 24.14 2.745 24.43 2.975 ;
      RECT 25.92 2.735 26.285 2.99 ;
      RECT 24.765 2.45 25.085 2.71 ;
      RECT 24.765 2.45 25.23 2.695 ;
      RECT 25.09 2.07 25.23 2.695 ;
      RECT 25.09 2.07 25.355 2.21 ;
      RECT 25.62 1.905 25.91 2.135 ;
      RECT 25.215 1.95 25.91 2.09 ;
      RECT 24.66 3.29 24.95 3.815 ;
      RECT 24.645 3.29 24.965 3.55 ;
      RECT 24.385 1.89 24.705 2.15 ;
      RECT 24.385 1.905 24.95 2.135 ;
      RECT 23.66 3.585 23.95 3.815 ;
      RECT 23.855 2.23 23.995 3.77 ;
      RECT 23.9 2.185 24.19 2.415 ;
      RECT 23.495 2.23 24.19 2.37 ;
      RECT 23.495 2.07 23.635 2.37 ;
      RECT 22.035 2.07 23.635 2.21 ;
      RECT 21.945 1.89 22.265 2.15 ;
      RECT 21.945 1.905 22.51 2.15 ;
      RECT 21.055 2.93 23.635 3.07 ;
      RECT 23.42 2.745 23.71 2.975 ;
      RECT 20.98 2.745 21.645 2.975 ;
      RECT 21.325 2.73 21.645 3.07 ;
      RECT 22.325 2.45 22.645 2.71 ;
      RECT 22.325 2.465 22.75 2.695 ;
      RECT 20.965 2.17 21.285 2.43 ;
      RECT 21.46 2.185 21.75 2.415 ;
      RECT 20.965 2.23 21.75 2.37 ;
      RECT 21.085 3.29 21.405 3.55 ;
      RECT 20.245 3.29 20.565 3.55 ;
      RECT 21.085 3.305 21.51 3.535 ;
      RECT 20.245 3.35 21.51 3.49 ;
      RECT 19.78 3.025 20.07 3.255 ;
      RECT 19.855 1.95 19.995 3.255 ;
      RECT 19.505 2.45 19.995 2.71 ;
      RECT 19.26 2.465 19.995 2.695 ;
      RECT 20.26 1.905 20.55 2.135 ;
      RECT 19.855 1.95 20.55 2.09 ;
      RECT 19.02 3.305 19.31 3.535 ;
      RECT 19.02 3.305 19.475 3.49 ;
      RECT 19.335 2.93 19.475 3.49 ;
      RECT 18.975 2.93 19.475 3.07 ;
      RECT 18.975 1.95 19.115 3.07 ;
      RECT 18.765 1.89 19.085 2.15 ;
      RECT 18.525 3.57 18.845 3.83 ;
      RECT 17.82 3.585 18.11 3.815 ;
      RECT 17.82 3.63 18.845 3.77 ;
      RECT 17.895 3.58 18.155 3.77 ;
      RECT 18.285 2.45 18.605 2.71 ;
      RECT 18.285 2.465 18.83 2.695 ;
      RECT 18.285 3.01 18.605 3.27 ;
      RECT 18.285 3.025 18.83 3.255 ;
      RECT 17.325 3.01 17.645 3.27 ;
      RECT 17.415 1.95 17.555 3.27 ;
      RECT 17.82 1.905 18.11 2.135 ;
      RECT 17.415 1.95 18.11 2.09 ;
      RECT 15.735 2.365 16.025 2.595 ;
      RECT 15.795 0.885 15.965 2.595 ;
      RECT 15.77 1.1 16.11 1.45 ;
      RECT 15.735 0.885 16.025 1.115 ;
      RECT 15.735 7.765 16.025 7.995 ;
      RECT 15.795 6.285 15.965 7.995 ;
      RECT 15.735 6.285 16.025 6.515 ;
      RECT 15.325 2.735 15.655 2.965 ;
      RECT 15.325 2.765 15.825 2.935 ;
      RECT 15.325 2.395 15.515 2.965 ;
      RECT 14.745 2.365 15.035 2.595 ;
      RECT 14.745 2.395 15.515 2.565 ;
      RECT 14.805 0.885 14.975 2.595 ;
      RECT 14.745 0.885 15.035 1.115 ;
      RECT 14.745 7.765 15.035 7.995 ;
      RECT 14.805 6.285 14.975 7.995 ;
      RECT 14.745 6.285 15.035 6.515 ;
      RECT 14.745 6.325 15.595 6.485 ;
      RECT 15.425 5.915 15.595 6.485 ;
      RECT 14.745 6.32 15.135 6.485 ;
      RECT 15.365 5.915 15.655 6.145 ;
      RECT 15.365 5.945 15.825 6.115 ;
      RECT 14.375 2.735 14.665 2.965 ;
      RECT 14.375 2.765 14.835 2.935 ;
      RECT 14.435 1.655 14.6 2.965 ;
      RECT 12.95 1.625 13.24 1.855 ;
      RECT 12.95 1.655 14.6 1.825 ;
      RECT 13.01 0.885 13.18 1.855 ;
      RECT 12.95 0.885 13.24 1.115 ;
      RECT 12.95 7.765 13.24 7.995 ;
      RECT 13.01 7.025 13.18 7.995 ;
      RECT 13.01 7.12 14.6 7.29 ;
      RECT 14.43 5.915 14.6 7.29 ;
      RECT 12.95 7.025 13.24 7.255 ;
      RECT 14.375 5.915 14.665 6.145 ;
      RECT 14.375 5.945 14.835 6.115 ;
      RECT 13.38 1.965 13.73 2.315 ;
      RECT 13.21 2.025 13.73 2.195 ;
      RECT 13.405 6.655 13.73 6.98 ;
      RECT 13.38 6.655 13.73 6.885 ;
      RECT 13.21 6.685 13.73 6.855 ;
      RECT 12.605 2.365 12.925 2.685 ;
      RECT 12.575 2.365 12.925 2.595 ;
      RECT 11.075 2.395 12.925 2.565 ;
      RECT 11.075 1.46 11.245 2.565 ;
      RECT 10.985 1.46 11.325 1.81 ;
      RECT 12.605 6.28 12.925 6.605 ;
      RECT 12.575 6.285 12.925 6.515 ;
      RECT 12.405 6.315 12.925 6.485 ;
      RECT 11.565 2.705 11.905 3.055 ;
      RECT 11.565 2.765 12.04 2.935 ;
      RECT 11.555 5.84 11.895 6.19 ;
      RECT 11.555 5.945 12.04 6.115 ;
      RECT 9.06 2.465 9.35 2.695 ;
      RECT 9.06 2.465 9.515 2.65 ;
      RECT 9.375 2.37 9.995 2.51 ;
      RECT 9.765 2.17 10.085 2.43 ;
      RECT 8.155 2.93 9.755 3.07 ;
      RECT 8.155 2.93 9.92 3.055 ;
      RECT 9.645 2.73 9.965 2.99 ;
      RECT 9.6 2.745 10.07 2.975 ;
      RECT 7.82 2.79 8.295 2.975 ;
      RECT 7.82 2.745 8.11 2.975 ;
      RECT 9.6 2.735 9.965 2.99 ;
      RECT 8.445 2.45 8.765 2.71 ;
      RECT 8.445 2.45 8.91 2.695 ;
      RECT 8.77 2.07 8.91 2.695 ;
      RECT 8.77 2.07 9.035 2.21 ;
      RECT 9.3 1.905 9.59 2.135 ;
      RECT 8.895 1.95 9.59 2.09 ;
      RECT 8.34 3.29 8.63 3.815 ;
      RECT 8.325 3.29 8.645 3.55 ;
      RECT 8.065 1.89 8.385 2.15 ;
      RECT 8.065 1.905 8.63 2.135 ;
      RECT 7.34 3.585 7.63 3.815 ;
      RECT 7.535 2.23 7.675 3.77 ;
      RECT 7.58 2.185 7.87 2.415 ;
      RECT 7.175 2.23 7.87 2.37 ;
      RECT 7.175 2.07 7.315 2.37 ;
      RECT 5.715 2.07 7.315 2.21 ;
      RECT 5.625 1.89 5.945 2.15 ;
      RECT 5.625 1.905 6.19 2.15 ;
      RECT 4.735 2.93 7.315 3.07 ;
      RECT 7.1 2.745 7.39 2.975 ;
      RECT 4.66 2.745 5.325 2.975 ;
      RECT 5.005 2.73 5.325 3.07 ;
      RECT 6.005 2.45 6.325 2.71 ;
      RECT 6.005 2.465 6.43 2.695 ;
      RECT 4.645 2.17 4.965 2.43 ;
      RECT 5.14 2.185 5.43 2.415 ;
      RECT 4.645 2.23 5.43 2.37 ;
      RECT 4.765 3.29 5.085 3.55 ;
      RECT 3.925 3.29 4.245 3.55 ;
      RECT 4.765 3.305 5.19 3.535 ;
      RECT 3.925 3.35 5.19 3.49 ;
      RECT 3.46 3.025 3.75 3.255 ;
      RECT 3.535 1.95 3.675 3.255 ;
      RECT 3.185 2.45 3.675 2.71 ;
      RECT 2.94 2.465 3.675 2.695 ;
      RECT 3.94 1.905 4.23 2.135 ;
      RECT 3.535 1.95 4.23 2.09 ;
      RECT 2.7 3.305 2.99 3.535 ;
      RECT 2.7 3.305 3.155 3.49 ;
      RECT 3.015 2.93 3.155 3.49 ;
      RECT 2.655 2.93 3.155 3.07 ;
      RECT 2.655 1.95 2.795 3.07 ;
      RECT 2.445 1.89 2.765 2.15 ;
      RECT 2.205 3.57 2.525 3.83 ;
      RECT 1.5 3.585 1.79 3.815 ;
      RECT 1.5 3.63 2.525 3.77 ;
      RECT 1.575 3.58 1.835 3.77 ;
      RECT 1.965 2.45 2.285 2.71 ;
      RECT 1.965 2.465 2.51 2.695 ;
      RECT 1.965 3.01 2.285 3.27 ;
      RECT 1.965 3.025 2.51 3.255 ;
      RECT 1.005 3.01 1.325 3.27 ;
      RECT 1.095 1.95 1.235 3.27 ;
      RECT 1.5 1.905 1.79 2.135 ;
      RECT 1.095 1.95 1.79 2.09 ;
      RECT 0.01 8.575 81.625 8.88 ;
      RECT 71.895 2.45 72.215 2.71 ;
      RECT 69.455 2.45 69.775 2.71 ;
      RECT 55.57 2.45 55.89 2.71 ;
      RECT 53.13 2.45 53.45 2.71 ;
      RECT 39.25 2.45 39.57 2.71 ;
      RECT 36.81 2.45 37.13 2.71 ;
      RECT 22.925 2.45 23.245 2.71 ;
      RECT 20.485 2.45 20.805 2.71 ;
      RECT 6.605 2.45 6.925 2.71 ;
      RECT 4.165 2.45 4.485 2.71 ;
    LAYER mcon ;
      RECT 81.085 0.915 81.255 1.085 ;
      RECT 81.085 2.395 81.255 2.565 ;
      RECT 81.085 6.315 81.255 6.485 ;
      RECT 81.085 7.795 81.255 7.965 ;
      RECT 80.735 0.105 80.905 0.275 ;
      RECT 80.735 4.165 80.905 4.335 ;
      RECT 80.735 4.545 80.905 4.715 ;
      RECT 80.735 8.605 80.905 8.775 ;
      RECT 80.715 2.765 80.885 2.935 ;
      RECT 80.715 5.945 80.885 6.115 ;
      RECT 80.095 0.915 80.265 1.085 ;
      RECT 80.095 2.395 80.265 2.565 ;
      RECT 80.095 6.315 80.265 6.485 ;
      RECT 80.095 7.795 80.265 7.965 ;
      RECT 79.745 0.105 79.915 0.275 ;
      RECT 79.745 4.165 79.915 4.335 ;
      RECT 79.745 4.545 79.915 4.715 ;
      RECT 79.745 8.605 79.915 8.775 ;
      RECT 79.725 2.765 79.895 2.935 ;
      RECT 79.725 5.945 79.895 6.115 ;
      RECT 79.04 0.105 79.21 0.275 ;
      RECT 79.04 4.165 79.21 4.335 ;
      RECT 79.04 4.545 79.21 4.715 ;
      RECT 79.04 8.605 79.21 8.775 ;
      RECT 78.73 2.025 78.9 2.195 ;
      RECT 78.73 6.685 78.9 6.855 ;
      RECT 78.36 0.105 78.53 0.275 ;
      RECT 78.36 8.605 78.53 8.775 ;
      RECT 78.3 0.915 78.47 1.085 ;
      RECT 78.3 1.655 78.47 1.825 ;
      RECT 78.3 7.055 78.47 7.225 ;
      RECT 78.3 7.795 78.47 7.965 ;
      RECT 77.925 2.395 78.095 2.565 ;
      RECT 77.925 6.315 78.095 6.485 ;
      RECT 77.68 0.105 77.85 0.275 ;
      RECT 77.68 8.605 77.85 8.775 ;
      RECT 77 0.105 77.17 0.275 ;
      RECT 77 8.605 77.17 8.775 ;
      RECT 76.93 2.765 77.1 2.935 ;
      RECT 76.93 5.945 77.1 6.115 ;
      RECT 75.385 1.415 75.555 1.585 ;
      RECT 75.385 4.135 75.555 4.305 ;
      RECT 75.13 2.775 75.3 2.945 ;
      RECT 74.925 1.415 75.095 1.585 ;
      RECT 74.925 4.135 75.095 4.305 ;
      RECT 74.65 1.935 74.82 2.105 ;
      RECT 74.465 1.415 74.635 1.585 ;
      RECT 74.465 4.135 74.635 4.305 ;
      RECT 74.41 2.495 74.58 2.665 ;
      RECT 74.005 1.415 74.175 1.585 ;
      RECT 74.005 4.135 74.175 4.305 ;
      RECT 73.93 2.495 74.1 2.665 ;
      RECT 73.69 1.935 73.86 2.105 ;
      RECT 73.69 3.615 73.86 3.785 ;
      RECT 73.545 1.415 73.715 1.585 ;
      RECT 73.545 4.135 73.715 4.305 ;
      RECT 73.17 2.775 73.34 2.945 ;
      RECT 73.085 1.415 73.255 1.585 ;
      RECT 73.085 4.135 73.255 4.305 ;
      RECT 72.93 2.215 73.1 2.385 ;
      RECT 72.69 3.615 72.86 3.785 ;
      RECT 72.625 1.415 72.795 1.585 ;
      RECT 72.625 4.135 72.795 4.305 ;
      RECT 72.45 2.775 72.62 2.945 ;
      RECT 72.165 1.415 72.335 1.585 ;
      RECT 72.165 4.135 72.335 4.305 ;
      RECT 71.97 2.495 72.14 2.665 ;
      RECT 71.705 1.415 71.875 1.585 ;
      RECT 71.705 4.135 71.875 4.305 ;
      RECT 71.49 2.495 71.66 2.665 ;
      RECT 71.25 1.935 71.42 2.105 ;
      RECT 71.245 1.415 71.415 1.585 ;
      RECT 71.245 4.135 71.415 4.305 ;
      RECT 70.785 1.415 70.955 1.585 ;
      RECT 70.785 4.135 70.955 4.305 ;
      RECT 70.49 2.215 70.66 2.385 ;
      RECT 70.325 1.415 70.495 1.585 ;
      RECT 70.325 4.135 70.495 4.305 ;
      RECT 70.25 3.335 70.42 3.505 ;
      RECT 70.01 2.775 70.18 2.945 ;
      RECT 69.865 1.415 70.035 1.585 ;
      RECT 69.865 4.135 70.035 4.305 ;
      RECT 69.53 2.495 69.7 2.665 ;
      RECT 69.405 1.415 69.575 1.585 ;
      RECT 69.405 4.135 69.575 4.305 ;
      RECT 69.29 1.935 69.46 2.105 ;
      RECT 69.29 3.335 69.46 3.505 ;
      RECT 68.945 1.415 69.115 1.585 ;
      RECT 68.945 4.135 69.115 4.305 ;
      RECT 68.81 3.055 68.98 3.225 ;
      RECT 68.485 1.415 68.655 1.585 ;
      RECT 68.485 4.135 68.655 4.305 ;
      RECT 68.29 2.495 68.46 2.665 ;
      RECT 68.05 3.335 68.22 3.505 ;
      RECT 68.025 1.415 68.195 1.585 ;
      RECT 68.025 4.135 68.195 4.305 ;
      RECT 67.81 1.935 67.98 2.105 ;
      RECT 67.57 2.495 67.74 2.665 ;
      RECT 67.57 3.055 67.74 3.225 ;
      RECT 67.565 1.415 67.735 1.585 ;
      RECT 67.565 4.135 67.735 4.305 ;
      RECT 67.105 1.415 67.275 1.585 ;
      RECT 67.105 4.135 67.275 4.305 ;
      RECT 66.85 1.935 67.02 2.105 ;
      RECT 66.85 3.615 67.02 3.785 ;
      RECT 66.645 1.415 66.815 1.585 ;
      RECT 66.645 4.135 66.815 4.305 ;
      RECT 66.37 3.055 66.54 3.225 ;
      RECT 66.185 1.415 66.355 1.585 ;
      RECT 66.185 4.135 66.355 4.305 ;
      RECT 64.76 0.915 64.93 1.085 ;
      RECT 64.76 2.395 64.93 2.565 ;
      RECT 64.76 6.315 64.93 6.485 ;
      RECT 64.76 7.795 64.93 7.965 ;
      RECT 64.41 0.105 64.58 0.275 ;
      RECT 64.41 4.165 64.58 4.335 ;
      RECT 64.41 4.545 64.58 4.715 ;
      RECT 64.41 8.605 64.58 8.775 ;
      RECT 64.39 2.765 64.56 2.935 ;
      RECT 64.39 5.945 64.56 6.115 ;
      RECT 63.77 0.915 63.94 1.085 ;
      RECT 63.77 2.395 63.94 2.565 ;
      RECT 63.77 6.315 63.94 6.485 ;
      RECT 63.77 7.795 63.94 7.965 ;
      RECT 63.42 0.105 63.59 0.275 ;
      RECT 63.42 4.165 63.59 4.335 ;
      RECT 63.42 4.545 63.59 4.715 ;
      RECT 63.42 8.605 63.59 8.775 ;
      RECT 63.4 2.765 63.57 2.935 ;
      RECT 63.4 5.945 63.57 6.115 ;
      RECT 62.715 0.105 62.885 0.275 ;
      RECT 62.715 4.165 62.885 4.335 ;
      RECT 62.715 4.545 62.885 4.715 ;
      RECT 62.715 8.605 62.885 8.775 ;
      RECT 62.405 2.025 62.575 2.195 ;
      RECT 62.405 6.685 62.575 6.855 ;
      RECT 62.035 0.105 62.205 0.275 ;
      RECT 62.035 8.605 62.205 8.775 ;
      RECT 61.975 0.915 62.145 1.085 ;
      RECT 61.975 1.655 62.145 1.825 ;
      RECT 61.975 7.055 62.145 7.225 ;
      RECT 61.975 7.795 62.145 7.965 ;
      RECT 61.6 2.395 61.77 2.565 ;
      RECT 61.6 6.315 61.77 6.485 ;
      RECT 61.355 0.105 61.525 0.275 ;
      RECT 61.355 8.605 61.525 8.775 ;
      RECT 60.675 0.105 60.845 0.275 ;
      RECT 60.675 8.605 60.845 8.775 ;
      RECT 60.605 2.765 60.775 2.935 ;
      RECT 60.605 5.945 60.775 6.115 ;
      RECT 59.06 1.415 59.23 1.585 ;
      RECT 59.06 4.135 59.23 4.305 ;
      RECT 58.805 2.775 58.975 2.945 ;
      RECT 58.6 1.415 58.77 1.585 ;
      RECT 58.6 4.135 58.77 4.305 ;
      RECT 58.325 1.935 58.495 2.105 ;
      RECT 58.14 1.415 58.31 1.585 ;
      RECT 58.14 4.135 58.31 4.305 ;
      RECT 58.085 2.495 58.255 2.665 ;
      RECT 57.68 1.415 57.85 1.585 ;
      RECT 57.68 4.135 57.85 4.305 ;
      RECT 57.605 2.495 57.775 2.665 ;
      RECT 57.365 1.935 57.535 2.105 ;
      RECT 57.365 3.615 57.535 3.785 ;
      RECT 57.22 1.415 57.39 1.585 ;
      RECT 57.22 4.135 57.39 4.305 ;
      RECT 56.845 2.775 57.015 2.945 ;
      RECT 56.76 1.415 56.93 1.585 ;
      RECT 56.76 4.135 56.93 4.305 ;
      RECT 56.605 2.215 56.775 2.385 ;
      RECT 56.365 3.615 56.535 3.785 ;
      RECT 56.3 1.415 56.47 1.585 ;
      RECT 56.3 4.135 56.47 4.305 ;
      RECT 56.125 2.775 56.295 2.945 ;
      RECT 55.84 1.415 56.01 1.585 ;
      RECT 55.84 4.135 56.01 4.305 ;
      RECT 55.645 2.495 55.815 2.665 ;
      RECT 55.38 1.415 55.55 1.585 ;
      RECT 55.38 4.135 55.55 4.305 ;
      RECT 55.165 2.495 55.335 2.665 ;
      RECT 54.925 1.935 55.095 2.105 ;
      RECT 54.92 1.415 55.09 1.585 ;
      RECT 54.92 4.135 55.09 4.305 ;
      RECT 54.46 1.415 54.63 1.585 ;
      RECT 54.46 4.135 54.63 4.305 ;
      RECT 54.165 2.215 54.335 2.385 ;
      RECT 54 1.415 54.17 1.585 ;
      RECT 54 4.135 54.17 4.305 ;
      RECT 53.925 3.335 54.095 3.505 ;
      RECT 53.685 2.775 53.855 2.945 ;
      RECT 53.54 1.415 53.71 1.585 ;
      RECT 53.54 4.135 53.71 4.305 ;
      RECT 53.205 2.495 53.375 2.665 ;
      RECT 53.08 1.415 53.25 1.585 ;
      RECT 53.08 4.135 53.25 4.305 ;
      RECT 52.965 1.935 53.135 2.105 ;
      RECT 52.965 3.335 53.135 3.505 ;
      RECT 52.62 1.415 52.79 1.585 ;
      RECT 52.62 4.135 52.79 4.305 ;
      RECT 52.485 3.055 52.655 3.225 ;
      RECT 52.16 1.415 52.33 1.585 ;
      RECT 52.16 4.135 52.33 4.305 ;
      RECT 51.965 2.495 52.135 2.665 ;
      RECT 51.725 3.335 51.895 3.505 ;
      RECT 51.7 1.415 51.87 1.585 ;
      RECT 51.7 4.135 51.87 4.305 ;
      RECT 51.485 1.935 51.655 2.105 ;
      RECT 51.245 2.495 51.415 2.665 ;
      RECT 51.245 3.055 51.415 3.225 ;
      RECT 51.24 1.415 51.41 1.585 ;
      RECT 51.24 4.135 51.41 4.305 ;
      RECT 50.78 1.415 50.95 1.585 ;
      RECT 50.78 4.135 50.95 4.305 ;
      RECT 50.525 1.935 50.695 2.105 ;
      RECT 50.525 3.615 50.695 3.785 ;
      RECT 50.32 1.415 50.49 1.585 ;
      RECT 50.32 4.135 50.49 4.305 ;
      RECT 50.045 3.055 50.215 3.225 ;
      RECT 49.86 1.415 50.03 1.585 ;
      RECT 49.86 4.135 50.03 4.305 ;
      RECT 48.44 0.915 48.61 1.085 ;
      RECT 48.44 2.395 48.61 2.565 ;
      RECT 48.44 6.315 48.61 6.485 ;
      RECT 48.44 7.795 48.61 7.965 ;
      RECT 48.09 0.105 48.26 0.275 ;
      RECT 48.09 4.165 48.26 4.335 ;
      RECT 48.09 4.545 48.26 4.715 ;
      RECT 48.09 8.605 48.26 8.775 ;
      RECT 48.07 2.765 48.24 2.935 ;
      RECT 48.07 5.945 48.24 6.115 ;
      RECT 47.45 0.915 47.62 1.085 ;
      RECT 47.45 2.395 47.62 2.565 ;
      RECT 47.45 6.315 47.62 6.485 ;
      RECT 47.45 7.795 47.62 7.965 ;
      RECT 47.1 0.105 47.27 0.275 ;
      RECT 47.1 4.165 47.27 4.335 ;
      RECT 47.1 4.545 47.27 4.715 ;
      RECT 47.1 8.605 47.27 8.775 ;
      RECT 47.08 2.765 47.25 2.935 ;
      RECT 47.08 5.945 47.25 6.115 ;
      RECT 46.395 0.105 46.565 0.275 ;
      RECT 46.395 4.165 46.565 4.335 ;
      RECT 46.395 4.545 46.565 4.715 ;
      RECT 46.395 8.605 46.565 8.775 ;
      RECT 46.085 2.025 46.255 2.195 ;
      RECT 46.085 6.685 46.255 6.855 ;
      RECT 45.715 0.105 45.885 0.275 ;
      RECT 45.715 8.605 45.885 8.775 ;
      RECT 45.655 0.915 45.825 1.085 ;
      RECT 45.655 1.655 45.825 1.825 ;
      RECT 45.655 7.055 45.825 7.225 ;
      RECT 45.655 7.795 45.825 7.965 ;
      RECT 45.28 2.395 45.45 2.565 ;
      RECT 45.28 6.315 45.45 6.485 ;
      RECT 45.035 0.105 45.205 0.275 ;
      RECT 45.035 8.605 45.205 8.775 ;
      RECT 44.355 0.105 44.525 0.275 ;
      RECT 44.355 8.605 44.525 8.775 ;
      RECT 44.285 2.765 44.455 2.935 ;
      RECT 44.285 5.945 44.455 6.115 ;
      RECT 42.74 1.415 42.91 1.585 ;
      RECT 42.74 4.135 42.91 4.305 ;
      RECT 42.485 2.775 42.655 2.945 ;
      RECT 42.28 1.415 42.45 1.585 ;
      RECT 42.28 4.135 42.45 4.305 ;
      RECT 42.005 1.935 42.175 2.105 ;
      RECT 41.82 1.415 41.99 1.585 ;
      RECT 41.82 4.135 41.99 4.305 ;
      RECT 41.765 2.495 41.935 2.665 ;
      RECT 41.36 1.415 41.53 1.585 ;
      RECT 41.36 4.135 41.53 4.305 ;
      RECT 41.285 2.495 41.455 2.665 ;
      RECT 41.045 1.935 41.215 2.105 ;
      RECT 41.045 3.615 41.215 3.785 ;
      RECT 40.9 1.415 41.07 1.585 ;
      RECT 40.9 4.135 41.07 4.305 ;
      RECT 40.525 2.775 40.695 2.945 ;
      RECT 40.44 1.415 40.61 1.585 ;
      RECT 40.44 4.135 40.61 4.305 ;
      RECT 40.285 2.215 40.455 2.385 ;
      RECT 40.045 3.615 40.215 3.785 ;
      RECT 39.98 1.415 40.15 1.585 ;
      RECT 39.98 4.135 40.15 4.305 ;
      RECT 39.805 2.775 39.975 2.945 ;
      RECT 39.52 1.415 39.69 1.585 ;
      RECT 39.52 4.135 39.69 4.305 ;
      RECT 39.325 2.495 39.495 2.665 ;
      RECT 39.06 1.415 39.23 1.585 ;
      RECT 39.06 4.135 39.23 4.305 ;
      RECT 38.845 2.495 39.015 2.665 ;
      RECT 38.605 1.935 38.775 2.105 ;
      RECT 38.6 1.415 38.77 1.585 ;
      RECT 38.6 4.135 38.77 4.305 ;
      RECT 38.14 1.415 38.31 1.585 ;
      RECT 38.14 4.135 38.31 4.305 ;
      RECT 37.845 2.215 38.015 2.385 ;
      RECT 37.68 1.415 37.85 1.585 ;
      RECT 37.68 4.135 37.85 4.305 ;
      RECT 37.605 3.335 37.775 3.505 ;
      RECT 37.365 2.775 37.535 2.945 ;
      RECT 37.22 1.415 37.39 1.585 ;
      RECT 37.22 4.135 37.39 4.305 ;
      RECT 36.885 2.495 37.055 2.665 ;
      RECT 36.76 1.415 36.93 1.585 ;
      RECT 36.76 4.135 36.93 4.305 ;
      RECT 36.645 1.935 36.815 2.105 ;
      RECT 36.645 3.335 36.815 3.505 ;
      RECT 36.3 1.415 36.47 1.585 ;
      RECT 36.3 4.135 36.47 4.305 ;
      RECT 36.165 3.055 36.335 3.225 ;
      RECT 35.84 1.415 36.01 1.585 ;
      RECT 35.84 4.135 36.01 4.305 ;
      RECT 35.645 2.495 35.815 2.665 ;
      RECT 35.405 3.335 35.575 3.505 ;
      RECT 35.38 1.415 35.55 1.585 ;
      RECT 35.38 4.135 35.55 4.305 ;
      RECT 35.165 1.935 35.335 2.105 ;
      RECT 34.925 2.495 35.095 2.665 ;
      RECT 34.925 3.055 35.095 3.225 ;
      RECT 34.92 1.415 35.09 1.585 ;
      RECT 34.92 4.135 35.09 4.305 ;
      RECT 34.46 1.415 34.63 1.585 ;
      RECT 34.46 4.135 34.63 4.305 ;
      RECT 34.205 1.935 34.375 2.105 ;
      RECT 34.205 3.615 34.375 3.785 ;
      RECT 34 1.415 34.17 1.585 ;
      RECT 34 4.135 34.17 4.305 ;
      RECT 33.725 3.055 33.895 3.225 ;
      RECT 33.54 1.415 33.71 1.585 ;
      RECT 33.54 4.135 33.71 4.305 ;
      RECT 32.115 0.915 32.285 1.085 ;
      RECT 32.115 2.395 32.285 2.565 ;
      RECT 32.115 6.315 32.285 6.485 ;
      RECT 32.115 7.795 32.285 7.965 ;
      RECT 31.765 0.105 31.935 0.275 ;
      RECT 31.765 4.165 31.935 4.335 ;
      RECT 31.765 4.545 31.935 4.715 ;
      RECT 31.765 8.605 31.935 8.775 ;
      RECT 31.745 2.765 31.915 2.935 ;
      RECT 31.745 5.945 31.915 6.115 ;
      RECT 31.125 0.915 31.295 1.085 ;
      RECT 31.125 2.395 31.295 2.565 ;
      RECT 31.125 6.315 31.295 6.485 ;
      RECT 31.125 7.795 31.295 7.965 ;
      RECT 30.775 0.105 30.945 0.275 ;
      RECT 30.775 4.165 30.945 4.335 ;
      RECT 30.775 4.545 30.945 4.715 ;
      RECT 30.775 8.605 30.945 8.775 ;
      RECT 30.755 2.765 30.925 2.935 ;
      RECT 30.755 5.945 30.925 6.115 ;
      RECT 30.07 0.105 30.24 0.275 ;
      RECT 30.07 4.165 30.24 4.335 ;
      RECT 30.07 4.545 30.24 4.715 ;
      RECT 30.07 8.605 30.24 8.775 ;
      RECT 29.76 2.025 29.93 2.195 ;
      RECT 29.76 6.685 29.93 6.855 ;
      RECT 29.39 0.105 29.56 0.275 ;
      RECT 29.39 8.605 29.56 8.775 ;
      RECT 29.33 0.915 29.5 1.085 ;
      RECT 29.33 1.655 29.5 1.825 ;
      RECT 29.33 7.055 29.5 7.225 ;
      RECT 29.33 7.795 29.5 7.965 ;
      RECT 28.955 2.395 29.125 2.565 ;
      RECT 28.955 6.315 29.125 6.485 ;
      RECT 28.71 0.105 28.88 0.275 ;
      RECT 28.71 8.605 28.88 8.775 ;
      RECT 28.03 0.105 28.2 0.275 ;
      RECT 28.03 8.605 28.2 8.775 ;
      RECT 27.96 2.765 28.13 2.935 ;
      RECT 27.96 5.945 28.13 6.115 ;
      RECT 26.415 1.415 26.585 1.585 ;
      RECT 26.415 4.135 26.585 4.305 ;
      RECT 26.16 2.775 26.33 2.945 ;
      RECT 25.955 1.415 26.125 1.585 ;
      RECT 25.955 4.135 26.125 4.305 ;
      RECT 25.68 1.935 25.85 2.105 ;
      RECT 25.495 1.415 25.665 1.585 ;
      RECT 25.495 4.135 25.665 4.305 ;
      RECT 25.44 2.495 25.61 2.665 ;
      RECT 25.035 1.415 25.205 1.585 ;
      RECT 25.035 4.135 25.205 4.305 ;
      RECT 24.96 2.495 25.13 2.665 ;
      RECT 24.72 1.935 24.89 2.105 ;
      RECT 24.72 3.615 24.89 3.785 ;
      RECT 24.575 1.415 24.745 1.585 ;
      RECT 24.575 4.135 24.745 4.305 ;
      RECT 24.2 2.775 24.37 2.945 ;
      RECT 24.115 1.415 24.285 1.585 ;
      RECT 24.115 4.135 24.285 4.305 ;
      RECT 23.96 2.215 24.13 2.385 ;
      RECT 23.72 3.615 23.89 3.785 ;
      RECT 23.655 1.415 23.825 1.585 ;
      RECT 23.655 4.135 23.825 4.305 ;
      RECT 23.48 2.775 23.65 2.945 ;
      RECT 23.195 1.415 23.365 1.585 ;
      RECT 23.195 4.135 23.365 4.305 ;
      RECT 23 2.495 23.17 2.665 ;
      RECT 22.735 1.415 22.905 1.585 ;
      RECT 22.735 4.135 22.905 4.305 ;
      RECT 22.52 2.495 22.69 2.665 ;
      RECT 22.28 1.935 22.45 2.105 ;
      RECT 22.275 1.415 22.445 1.585 ;
      RECT 22.275 4.135 22.445 4.305 ;
      RECT 21.815 1.415 21.985 1.585 ;
      RECT 21.815 4.135 21.985 4.305 ;
      RECT 21.52 2.215 21.69 2.385 ;
      RECT 21.355 1.415 21.525 1.585 ;
      RECT 21.355 4.135 21.525 4.305 ;
      RECT 21.28 3.335 21.45 3.505 ;
      RECT 21.04 2.775 21.21 2.945 ;
      RECT 20.895 1.415 21.065 1.585 ;
      RECT 20.895 4.135 21.065 4.305 ;
      RECT 20.56 2.495 20.73 2.665 ;
      RECT 20.435 1.415 20.605 1.585 ;
      RECT 20.435 4.135 20.605 4.305 ;
      RECT 20.32 1.935 20.49 2.105 ;
      RECT 20.32 3.335 20.49 3.505 ;
      RECT 19.975 1.415 20.145 1.585 ;
      RECT 19.975 4.135 20.145 4.305 ;
      RECT 19.84 3.055 20.01 3.225 ;
      RECT 19.515 1.415 19.685 1.585 ;
      RECT 19.515 4.135 19.685 4.305 ;
      RECT 19.32 2.495 19.49 2.665 ;
      RECT 19.08 3.335 19.25 3.505 ;
      RECT 19.055 1.415 19.225 1.585 ;
      RECT 19.055 4.135 19.225 4.305 ;
      RECT 18.84 1.935 19.01 2.105 ;
      RECT 18.6 2.495 18.77 2.665 ;
      RECT 18.6 3.055 18.77 3.225 ;
      RECT 18.595 1.415 18.765 1.585 ;
      RECT 18.595 4.135 18.765 4.305 ;
      RECT 18.135 1.415 18.305 1.585 ;
      RECT 18.135 4.135 18.305 4.305 ;
      RECT 17.88 1.935 18.05 2.105 ;
      RECT 17.88 3.615 18.05 3.785 ;
      RECT 17.675 1.415 17.845 1.585 ;
      RECT 17.675 4.135 17.845 4.305 ;
      RECT 17.4 3.055 17.57 3.225 ;
      RECT 17.215 1.415 17.385 1.585 ;
      RECT 17.215 4.135 17.385 4.305 ;
      RECT 15.795 0.915 15.965 1.085 ;
      RECT 15.795 2.395 15.965 2.565 ;
      RECT 15.795 6.315 15.965 6.485 ;
      RECT 15.795 7.795 15.965 7.965 ;
      RECT 15.445 0.105 15.615 0.275 ;
      RECT 15.445 4.165 15.615 4.335 ;
      RECT 15.445 4.545 15.615 4.715 ;
      RECT 15.445 8.605 15.615 8.775 ;
      RECT 15.425 2.765 15.595 2.935 ;
      RECT 15.425 5.945 15.595 6.115 ;
      RECT 14.805 0.915 14.975 1.085 ;
      RECT 14.805 2.395 14.975 2.565 ;
      RECT 14.805 6.315 14.975 6.485 ;
      RECT 14.805 7.795 14.975 7.965 ;
      RECT 14.455 0.105 14.625 0.275 ;
      RECT 14.455 4.165 14.625 4.335 ;
      RECT 14.455 4.545 14.625 4.715 ;
      RECT 14.455 8.605 14.625 8.775 ;
      RECT 14.435 2.765 14.605 2.935 ;
      RECT 14.435 5.945 14.605 6.115 ;
      RECT 13.75 0.105 13.92 0.275 ;
      RECT 13.75 4.165 13.92 4.335 ;
      RECT 13.75 4.545 13.92 4.715 ;
      RECT 13.75 8.605 13.92 8.775 ;
      RECT 13.44 2.025 13.61 2.195 ;
      RECT 13.44 6.685 13.61 6.855 ;
      RECT 13.07 0.105 13.24 0.275 ;
      RECT 13.07 8.605 13.24 8.775 ;
      RECT 13.01 0.915 13.18 1.085 ;
      RECT 13.01 1.655 13.18 1.825 ;
      RECT 13.01 7.055 13.18 7.225 ;
      RECT 13.01 7.795 13.18 7.965 ;
      RECT 12.635 2.395 12.805 2.565 ;
      RECT 12.635 6.315 12.805 6.485 ;
      RECT 12.39 0.105 12.56 0.275 ;
      RECT 12.39 8.605 12.56 8.775 ;
      RECT 11.71 0.105 11.88 0.275 ;
      RECT 11.71 8.605 11.88 8.775 ;
      RECT 11.64 2.765 11.81 2.935 ;
      RECT 11.64 5.945 11.81 6.115 ;
      RECT 10.095 1.415 10.265 1.585 ;
      RECT 10.095 4.135 10.265 4.305 ;
      RECT 9.84 2.775 10.01 2.945 ;
      RECT 9.635 1.415 9.805 1.585 ;
      RECT 9.635 4.135 9.805 4.305 ;
      RECT 9.36 1.935 9.53 2.105 ;
      RECT 9.175 1.415 9.345 1.585 ;
      RECT 9.175 4.135 9.345 4.305 ;
      RECT 9.12 2.495 9.29 2.665 ;
      RECT 8.715 1.415 8.885 1.585 ;
      RECT 8.715 4.135 8.885 4.305 ;
      RECT 8.64 2.495 8.81 2.665 ;
      RECT 8.4 1.935 8.57 2.105 ;
      RECT 8.4 3.615 8.57 3.785 ;
      RECT 8.255 1.415 8.425 1.585 ;
      RECT 8.255 4.135 8.425 4.305 ;
      RECT 7.88 2.775 8.05 2.945 ;
      RECT 7.795 1.415 7.965 1.585 ;
      RECT 7.795 4.135 7.965 4.305 ;
      RECT 7.64 2.215 7.81 2.385 ;
      RECT 7.4 3.615 7.57 3.785 ;
      RECT 7.335 1.415 7.505 1.585 ;
      RECT 7.335 4.135 7.505 4.305 ;
      RECT 7.16 2.775 7.33 2.945 ;
      RECT 6.875 1.415 7.045 1.585 ;
      RECT 6.875 4.135 7.045 4.305 ;
      RECT 6.68 2.495 6.85 2.665 ;
      RECT 6.415 1.415 6.585 1.585 ;
      RECT 6.415 4.135 6.585 4.305 ;
      RECT 6.2 2.495 6.37 2.665 ;
      RECT 5.96 1.935 6.13 2.105 ;
      RECT 5.955 1.415 6.125 1.585 ;
      RECT 5.955 4.135 6.125 4.305 ;
      RECT 5.495 1.415 5.665 1.585 ;
      RECT 5.495 4.135 5.665 4.305 ;
      RECT 5.2 2.215 5.37 2.385 ;
      RECT 5.035 1.415 5.205 1.585 ;
      RECT 5.035 4.135 5.205 4.305 ;
      RECT 4.96 3.335 5.13 3.505 ;
      RECT 4.72 2.775 4.89 2.945 ;
      RECT 4.575 1.415 4.745 1.585 ;
      RECT 4.575 4.135 4.745 4.305 ;
      RECT 4.24 2.495 4.41 2.665 ;
      RECT 4.115 1.415 4.285 1.585 ;
      RECT 4.115 4.135 4.285 4.305 ;
      RECT 4 1.935 4.17 2.105 ;
      RECT 4 3.335 4.17 3.505 ;
      RECT 3.655 1.415 3.825 1.585 ;
      RECT 3.655 4.135 3.825 4.305 ;
      RECT 3.52 3.055 3.69 3.225 ;
      RECT 3.195 1.415 3.365 1.585 ;
      RECT 3.195 4.135 3.365 4.305 ;
      RECT 3 2.495 3.17 2.665 ;
      RECT 2.76 3.335 2.93 3.505 ;
      RECT 2.735 1.415 2.905 1.585 ;
      RECT 2.735 4.135 2.905 4.305 ;
      RECT 2.52 1.935 2.69 2.105 ;
      RECT 2.28 2.495 2.45 2.665 ;
      RECT 2.28 3.055 2.45 3.225 ;
      RECT 2.275 1.415 2.445 1.585 ;
      RECT 2.275 4.135 2.445 4.305 ;
      RECT 1.815 1.415 1.985 1.585 ;
      RECT 1.815 4.135 1.985 4.305 ;
      RECT 1.56 1.935 1.73 2.105 ;
      RECT 1.56 3.615 1.73 3.785 ;
      RECT 1.355 1.415 1.525 1.585 ;
      RECT 1.355 4.135 1.525 4.305 ;
      RECT 1.08 3.055 1.25 3.225 ;
      RECT 0.895 1.415 1.065 1.585 ;
      RECT 0.895 4.135 1.065 4.305 ;
    LAYER li ;
      RECT 74.17 0 74.34 2.085 ;
      RECT 72.21 0 72.38 2.085 ;
      RECT 69.77 0 69.94 2.085 ;
      RECT 68.81 0 68.98 2.085 ;
      RECT 68.29 0 68.46 2.085 ;
      RECT 67.33 0 67.5 2.085 ;
      RECT 66.37 0 66.54 2.085 ;
      RECT 57.845 0 58.015 2.085 ;
      RECT 55.885 0 56.055 2.085 ;
      RECT 53.445 0 53.615 2.085 ;
      RECT 52.485 0 52.655 2.085 ;
      RECT 51.965 0 52.135 2.085 ;
      RECT 51.005 0 51.175 2.085 ;
      RECT 50.045 0 50.215 2.085 ;
      RECT 41.525 0 41.695 2.085 ;
      RECT 39.565 0 39.735 2.085 ;
      RECT 37.125 0 37.295 2.085 ;
      RECT 36.165 0 36.335 2.085 ;
      RECT 35.645 0 35.815 2.085 ;
      RECT 34.685 0 34.855 2.085 ;
      RECT 33.725 0 33.895 2.085 ;
      RECT 25.2 0 25.37 2.085 ;
      RECT 23.24 0 23.41 2.085 ;
      RECT 20.8 0 20.97 2.085 ;
      RECT 19.84 0 20.01 2.085 ;
      RECT 19.32 0 19.49 2.085 ;
      RECT 18.36 0 18.53 2.085 ;
      RECT 17.4 0 17.57 2.085 ;
      RECT 8.88 0 9.05 2.085 ;
      RECT 6.92 0 7.09 2.085 ;
      RECT 4.48 0 4.65 2.085 ;
      RECT 3.52 0 3.69 2.085 ;
      RECT 3 0 3.17 2.085 ;
      RECT 2.04 0 2.21 2.085 ;
      RECT 1.08 0 1.25 2.085 ;
      RECT 72.14 0 72.38 1.595 ;
      RECT 70.59 0 70.785 1.595 ;
      RECT 68.465 0 68.66 1.595 ;
      RECT 66.165 0 66.36 1.595 ;
      RECT 55.815 0 56.055 1.595 ;
      RECT 54.265 0 54.46 1.595 ;
      RECT 52.14 0 52.335 1.595 ;
      RECT 49.84 0 50.035 1.595 ;
      RECT 39.495 0 39.735 1.595 ;
      RECT 37.945 0 38.14 1.595 ;
      RECT 35.82 0 36.015 1.595 ;
      RECT 33.52 0 33.715 1.595 ;
      RECT 23.17 0 23.41 1.595 ;
      RECT 21.62 0 21.815 1.595 ;
      RECT 19.495 0 19.69 1.595 ;
      RECT 17.195 0 17.39 1.595 ;
      RECT 6.85 0 7.09 1.595 ;
      RECT 5.3 0 5.495 1.595 ;
      RECT 3.175 0 3.37 1.595 ;
      RECT 0.875 0 1.07 1.595 ;
      RECT 66.04 0 75.855 1.585 ;
      RECT 49.715 0 59.53 1.585 ;
      RECT 33.395 0 43.21 1.585 ;
      RECT 17.07 0 26.885 1.585 ;
      RECT 0.75 0 10.565 1.585 ;
      RECT 80.655 0 80.825 0.935 ;
      RECT 79.665 0 79.835 0.935 ;
      RECT 76.92 0 77.09 0.935 ;
      RECT 64.33 0 64.5 0.935 ;
      RECT 63.34 0 63.51 0.935 ;
      RECT 60.595 0 60.765 0.935 ;
      RECT 48.01 0 48.18 0.935 ;
      RECT 47.02 0 47.19 0.935 ;
      RECT 44.275 0 44.445 0.935 ;
      RECT 31.685 0 31.855 0.935 ;
      RECT 30.695 0 30.865 0.935 ;
      RECT 27.95 0 28.12 0.935 ;
      RECT 15.365 0 15.535 0.935 ;
      RECT 14.375 0 14.545 0.935 ;
      RECT 11.63 0 11.8 0.935 ;
      RECT 0.005 0 81.625 0.305 ;
      RECT 80.655 3.405 80.825 5.475 ;
      RECT 79.665 3.405 79.835 5.475 ;
      RECT 76.92 3.405 77.09 5.475 ;
      RECT 64.33 3.405 64.5 5.475 ;
      RECT 63.34 3.405 63.51 5.475 ;
      RECT 60.595 3.405 60.765 5.475 ;
      RECT 48.01 3.405 48.18 5.475 ;
      RECT 47.02 3.405 47.19 5.475 ;
      RECT 44.275 3.405 44.445 5.475 ;
      RECT 31.685 3.405 31.855 5.475 ;
      RECT 30.695 3.405 30.865 5.475 ;
      RECT 27.95 3.405 28.12 5.475 ;
      RECT 15.365 3.405 15.535 5.475 ;
      RECT 14.375 3.405 14.545 5.475 ;
      RECT 11.63 3.405 11.8 5.475 ;
      RECT 0.005 4.135 81.625 4.745 ;
      RECT 75.13 3.635 75.3 4.745 ;
      RECT 74.17 3.635 74.34 4.745 ;
      RECT 71.73 3.635 71.9 4.745 ;
      RECT 70.73 3.635 70.9 4.745 ;
      RECT 69.77 3.635 69.94 4.745 ;
      RECT 67.33 3.635 67.5 4.745 ;
      RECT 58.805 3.635 58.975 4.745 ;
      RECT 57.845 3.635 58.015 4.745 ;
      RECT 55.405 3.635 55.575 4.745 ;
      RECT 54.405 3.635 54.575 4.745 ;
      RECT 53.445 3.635 53.615 4.745 ;
      RECT 51.005 3.635 51.175 4.745 ;
      RECT 42.485 3.635 42.655 4.745 ;
      RECT 41.525 3.635 41.695 4.745 ;
      RECT 39.085 3.635 39.255 4.745 ;
      RECT 38.085 3.635 38.255 4.745 ;
      RECT 37.125 3.635 37.295 4.745 ;
      RECT 34.685 3.635 34.855 4.745 ;
      RECT 26.16 3.635 26.33 4.745 ;
      RECT 25.2 3.635 25.37 4.745 ;
      RECT 22.76 3.635 22.93 4.745 ;
      RECT 21.76 3.635 21.93 4.745 ;
      RECT 20.8 3.635 20.97 4.745 ;
      RECT 18.36 3.635 18.53 4.745 ;
      RECT 9.84 3.635 10.01 4.745 ;
      RECT 8.88 3.635 9.05 4.745 ;
      RECT 6.44 3.635 6.61 4.745 ;
      RECT 5.44 3.635 5.61 4.745 ;
      RECT 4.48 3.635 4.65 4.745 ;
      RECT 2.04 3.635 2.21 4.745 ;
      RECT 0.01 8.575 81.625 8.88 ;
      RECT 80.655 7.945 80.825 8.88 ;
      RECT 79.665 7.945 79.835 8.88 ;
      RECT 76.92 7.945 77.09 8.88 ;
      RECT 64.33 7.945 64.5 8.88 ;
      RECT 63.34 7.945 63.51 8.88 ;
      RECT 60.595 7.945 60.765 8.88 ;
      RECT 48.01 7.945 48.18 8.88 ;
      RECT 47.02 7.945 47.19 8.88 ;
      RECT 44.275 7.945 44.445 8.88 ;
      RECT 31.685 7.945 31.855 8.88 ;
      RECT 30.695 7.945 30.865 8.88 ;
      RECT 27.95 7.945 28.12 8.88 ;
      RECT 15.365 7.945 15.535 8.88 ;
      RECT 14.375 7.945 14.545 8.88 ;
      RECT 11.63 7.945 11.8 8.88 ;
      RECT 80.715 1.74 80.885 2.935 ;
      RECT 80.715 1.74 81.18 1.91 ;
      RECT 80.715 6.97 81.18 7.14 ;
      RECT 80.715 5.945 80.885 7.14 ;
      RECT 79.725 1.74 79.895 2.935 ;
      RECT 79.725 1.74 80.19 1.91 ;
      RECT 79.725 6.97 80.19 7.14 ;
      RECT 79.725 5.945 79.895 7.14 ;
      RECT 77.87 2.635 78.04 3.865 ;
      RECT 77.925 0.855 78.095 2.805 ;
      RECT 77.87 0.575 78.04 1.025 ;
      RECT 77.87 7.855 78.04 8.305 ;
      RECT 77.925 6.075 78.095 8.025 ;
      RECT 77.87 5.015 78.04 6.245 ;
      RECT 77.35 0.575 77.52 3.865 ;
      RECT 77.35 2.075 77.755 2.405 ;
      RECT 77.35 1.235 77.755 1.565 ;
      RECT 77.35 5.015 77.52 8.305 ;
      RECT 77.35 7.315 77.755 7.645 ;
      RECT 77.35 6.475 77.755 6.805 ;
      RECT 74.65 1.835 74.82 2.105 ;
      RECT 74.65 1.835 75.38 2.005 ;
      RECT 75.13 2.575 75.3 2.945 ;
      RECT 74.81 2.575 75.3 2.745 ;
      RECT 74.57 3.225 74.9 3.395 ;
      RECT 73.81 3.055 74.82 3.225 ;
      RECT 73.81 2.575 73.98 3.225 ;
      RECT 73.93 2.495 74.1 2.825 ;
      RECT 73.09 3.225 73.42 3.395 ;
      RECT 71.17 3.225 72.46 3.395 ;
      RECT 72.21 3.14 73.34 3.31 ;
      RECT 72.93 2.215 73.34 2.385 ;
      RECT 73.17 1.755 73.34 2.385 ;
      RECT 73.17 2.575 73.34 2.945 ;
      RECT 72.85 2.575 73.34 2.745 ;
      RECT 70.41 2.575 71.74 2.745 ;
      RECT 71.49 2.495 71.66 2.745 ;
      RECT 70.49 2.175 70.66 2.385 ;
      RECT 70.49 2.175 70.98 2.345 ;
      RECT 69.17 3.335 69.46 3.505 ;
      RECT 69.17 2.575 69.34 3.505 ;
      RECT 68.97 2.575 69.34 2.745 ;
      RECT 67.97 2.575 68.46 2.745 ;
      RECT 68.29 2.495 68.46 2.745 ;
      RECT 68.05 3.335 68.46 3.505 ;
      RECT 68.29 3.145 68.46 3.505 ;
      RECT 67.09 3.055 67.74 3.225 ;
      RECT 67.09 2.495 67.26 3.225 ;
      RECT 66.73 3.615 67.02 3.785 ;
      RECT 66.73 2.575 66.9 3.785 ;
      RECT 66.53 2.575 66.9 2.745 ;
      RECT 64.39 1.74 64.56 2.935 ;
      RECT 64.39 1.74 64.855 1.91 ;
      RECT 64.39 6.97 64.855 7.14 ;
      RECT 64.39 5.945 64.56 7.14 ;
      RECT 63.4 1.74 63.57 2.935 ;
      RECT 63.4 1.74 63.865 1.91 ;
      RECT 63.4 6.97 63.865 7.14 ;
      RECT 63.4 5.945 63.57 7.14 ;
      RECT 61.545 2.635 61.715 3.865 ;
      RECT 61.6 0.855 61.77 2.805 ;
      RECT 61.545 0.575 61.715 1.025 ;
      RECT 61.545 7.855 61.715 8.305 ;
      RECT 61.6 6.075 61.77 8.025 ;
      RECT 61.545 5.015 61.715 6.245 ;
      RECT 61.025 0.575 61.195 3.865 ;
      RECT 61.025 2.075 61.43 2.405 ;
      RECT 61.025 1.235 61.43 1.565 ;
      RECT 61.025 5.015 61.195 8.305 ;
      RECT 61.025 7.315 61.43 7.645 ;
      RECT 61.025 6.475 61.43 6.805 ;
      RECT 58.325 1.835 58.495 2.105 ;
      RECT 58.325 1.835 59.055 2.005 ;
      RECT 58.805 2.575 58.975 2.945 ;
      RECT 58.485 2.575 58.975 2.745 ;
      RECT 58.245 3.225 58.575 3.395 ;
      RECT 57.485 3.055 58.495 3.225 ;
      RECT 57.485 2.575 57.655 3.225 ;
      RECT 57.605 2.495 57.775 2.825 ;
      RECT 56.765 3.225 57.095 3.395 ;
      RECT 54.845 3.225 56.135 3.395 ;
      RECT 55.885 3.14 57.015 3.31 ;
      RECT 56.605 2.215 57.015 2.385 ;
      RECT 56.845 1.755 57.015 2.385 ;
      RECT 56.845 2.575 57.015 2.945 ;
      RECT 56.525 2.575 57.015 2.745 ;
      RECT 54.085 2.575 55.415 2.745 ;
      RECT 55.165 2.495 55.335 2.745 ;
      RECT 54.165 2.175 54.335 2.385 ;
      RECT 54.165 2.175 54.655 2.345 ;
      RECT 52.845 3.335 53.135 3.505 ;
      RECT 52.845 2.575 53.015 3.505 ;
      RECT 52.645 2.575 53.015 2.745 ;
      RECT 51.645 2.575 52.135 2.745 ;
      RECT 51.965 2.495 52.135 2.745 ;
      RECT 51.725 3.335 52.135 3.505 ;
      RECT 51.965 3.145 52.135 3.505 ;
      RECT 50.765 3.055 51.415 3.225 ;
      RECT 50.765 2.495 50.935 3.225 ;
      RECT 50.405 3.615 50.695 3.785 ;
      RECT 50.405 2.575 50.575 3.785 ;
      RECT 50.205 2.575 50.575 2.745 ;
      RECT 48.07 1.74 48.24 2.935 ;
      RECT 48.07 1.74 48.535 1.91 ;
      RECT 48.07 6.97 48.535 7.14 ;
      RECT 48.07 5.945 48.24 7.14 ;
      RECT 47.08 1.74 47.25 2.935 ;
      RECT 47.08 1.74 47.545 1.91 ;
      RECT 47.08 6.97 47.545 7.14 ;
      RECT 47.08 5.945 47.25 7.14 ;
      RECT 45.225 2.635 45.395 3.865 ;
      RECT 45.28 0.855 45.45 2.805 ;
      RECT 45.225 0.575 45.395 1.025 ;
      RECT 45.225 7.855 45.395 8.305 ;
      RECT 45.28 6.075 45.45 8.025 ;
      RECT 45.225 5.015 45.395 6.245 ;
      RECT 44.705 0.575 44.875 3.865 ;
      RECT 44.705 2.075 45.11 2.405 ;
      RECT 44.705 1.235 45.11 1.565 ;
      RECT 44.705 5.015 44.875 8.305 ;
      RECT 44.705 7.315 45.11 7.645 ;
      RECT 44.705 6.475 45.11 6.805 ;
      RECT 42.005 1.835 42.175 2.105 ;
      RECT 42.005 1.835 42.735 2.005 ;
      RECT 42.485 2.575 42.655 2.945 ;
      RECT 42.165 2.575 42.655 2.745 ;
      RECT 41.925 3.225 42.255 3.395 ;
      RECT 41.165 3.055 42.175 3.225 ;
      RECT 41.165 2.575 41.335 3.225 ;
      RECT 41.285 2.495 41.455 2.825 ;
      RECT 40.445 3.225 40.775 3.395 ;
      RECT 38.525 3.225 39.815 3.395 ;
      RECT 39.565 3.14 40.695 3.31 ;
      RECT 40.285 2.215 40.695 2.385 ;
      RECT 40.525 1.755 40.695 2.385 ;
      RECT 40.525 2.575 40.695 2.945 ;
      RECT 40.205 2.575 40.695 2.745 ;
      RECT 37.765 2.575 39.095 2.745 ;
      RECT 38.845 2.495 39.015 2.745 ;
      RECT 37.845 2.175 38.015 2.385 ;
      RECT 37.845 2.175 38.335 2.345 ;
      RECT 36.525 3.335 36.815 3.505 ;
      RECT 36.525 2.575 36.695 3.505 ;
      RECT 36.325 2.575 36.695 2.745 ;
      RECT 35.325 2.575 35.815 2.745 ;
      RECT 35.645 2.495 35.815 2.745 ;
      RECT 35.405 3.335 35.815 3.505 ;
      RECT 35.645 3.145 35.815 3.505 ;
      RECT 34.445 3.055 35.095 3.225 ;
      RECT 34.445 2.495 34.615 3.225 ;
      RECT 34.085 3.615 34.375 3.785 ;
      RECT 34.085 2.575 34.255 3.785 ;
      RECT 33.885 2.575 34.255 2.745 ;
      RECT 31.745 1.74 31.915 2.935 ;
      RECT 31.745 1.74 32.21 1.91 ;
      RECT 31.745 6.97 32.21 7.14 ;
      RECT 31.745 5.945 31.915 7.14 ;
      RECT 30.755 1.74 30.925 2.935 ;
      RECT 30.755 1.74 31.22 1.91 ;
      RECT 30.755 6.97 31.22 7.14 ;
      RECT 30.755 5.945 30.925 7.14 ;
      RECT 28.9 2.635 29.07 3.865 ;
      RECT 28.955 0.855 29.125 2.805 ;
      RECT 28.9 0.575 29.07 1.025 ;
      RECT 28.9 7.855 29.07 8.305 ;
      RECT 28.955 6.075 29.125 8.025 ;
      RECT 28.9 5.015 29.07 6.245 ;
      RECT 28.38 0.575 28.55 3.865 ;
      RECT 28.38 2.075 28.785 2.405 ;
      RECT 28.38 1.235 28.785 1.565 ;
      RECT 28.38 5.015 28.55 8.305 ;
      RECT 28.38 7.315 28.785 7.645 ;
      RECT 28.38 6.475 28.785 6.805 ;
      RECT 25.68 1.835 25.85 2.105 ;
      RECT 25.68 1.835 26.41 2.005 ;
      RECT 26.16 2.575 26.33 2.945 ;
      RECT 25.84 2.575 26.33 2.745 ;
      RECT 25.6 3.225 25.93 3.395 ;
      RECT 24.84 3.055 25.85 3.225 ;
      RECT 24.84 2.575 25.01 3.225 ;
      RECT 24.96 2.495 25.13 2.825 ;
      RECT 24.12 3.225 24.45 3.395 ;
      RECT 22.2 3.225 23.49 3.395 ;
      RECT 23.24 3.14 24.37 3.31 ;
      RECT 23.96 2.215 24.37 2.385 ;
      RECT 24.2 1.755 24.37 2.385 ;
      RECT 24.2 2.575 24.37 2.945 ;
      RECT 23.88 2.575 24.37 2.745 ;
      RECT 21.44 2.575 22.77 2.745 ;
      RECT 22.52 2.495 22.69 2.745 ;
      RECT 21.52 2.175 21.69 2.385 ;
      RECT 21.52 2.175 22.01 2.345 ;
      RECT 20.2 3.335 20.49 3.505 ;
      RECT 20.2 2.575 20.37 3.505 ;
      RECT 20 2.575 20.37 2.745 ;
      RECT 19 2.575 19.49 2.745 ;
      RECT 19.32 2.495 19.49 2.745 ;
      RECT 19.08 3.335 19.49 3.505 ;
      RECT 19.32 3.145 19.49 3.505 ;
      RECT 18.12 3.055 18.77 3.225 ;
      RECT 18.12 2.495 18.29 3.225 ;
      RECT 17.76 3.615 18.05 3.785 ;
      RECT 17.76 2.575 17.93 3.785 ;
      RECT 17.56 2.575 17.93 2.745 ;
      RECT 15.425 1.74 15.595 2.935 ;
      RECT 15.425 1.74 15.89 1.91 ;
      RECT 15.425 6.97 15.89 7.14 ;
      RECT 15.425 5.945 15.595 7.14 ;
      RECT 14.435 1.74 14.605 2.935 ;
      RECT 14.435 1.74 14.9 1.91 ;
      RECT 14.435 6.97 14.9 7.14 ;
      RECT 14.435 5.945 14.605 7.14 ;
      RECT 12.58 2.635 12.75 3.865 ;
      RECT 12.635 0.855 12.805 2.805 ;
      RECT 12.58 0.575 12.75 1.025 ;
      RECT 12.58 7.855 12.75 8.305 ;
      RECT 12.635 6.075 12.805 8.025 ;
      RECT 12.58 5.015 12.75 6.245 ;
      RECT 12.06 0.575 12.23 3.865 ;
      RECT 12.06 2.075 12.465 2.405 ;
      RECT 12.06 1.235 12.465 1.565 ;
      RECT 12.06 5.015 12.23 8.305 ;
      RECT 12.06 7.315 12.465 7.645 ;
      RECT 12.06 6.475 12.465 6.805 ;
      RECT 9.36 1.835 9.53 2.105 ;
      RECT 9.36 1.835 10.09 2.005 ;
      RECT 9.84 2.575 10.01 2.945 ;
      RECT 9.52 2.575 10.01 2.745 ;
      RECT 9.28 3.225 9.61 3.395 ;
      RECT 8.52 3.055 9.53 3.225 ;
      RECT 8.52 2.575 8.69 3.225 ;
      RECT 8.64 2.495 8.81 2.825 ;
      RECT 7.8 3.225 8.13 3.395 ;
      RECT 5.88 3.225 7.17 3.395 ;
      RECT 6.92 3.14 8.05 3.31 ;
      RECT 7.64 2.215 8.05 2.385 ;
      RECT 7.88 1.755 8.05 2.385 ;
      RECT 7.88 2.575 8.05 2.945 ;
      RECT 7.56 2.575 8.05 2.745 ;
      RECT 5.12 2.575 6.45 2.745 ;
      RECT 6.2 2.495 6.37 2.745 ;
      RECT 5.2 2.175 5.37 2.385 ;
      RECT 5.2 2.175 5.69 2.345 ;
      RECT 3.88 3.335 4.17 3.505 ;
      RECT 3.88 2.575 4.05 3.505 ;
      RECT 3.68 2.575 4.05 2.745 ;
      RECT 2.68 2.575 3.17 2.745 ;
      RECT 3 2.495 3.17 2.745 ;
      RECT 2.76 3.335 3.17 3.505 ;
      RECT 3 3.145 3.17 3.505 ;
      RECT 1.8 3.055 2.45 3.225 ;
      RECT 1.8 2.495 1.97 3.225 ;
      RECT 1.44 3.615 1.73 3.785 ;
      RECT 1.44 2.575 1.61 3.785 ;
      RECT 1.24 2.575 1.61 2.745 ;
      RECT 81.085 0.575 81.255 1.085 ;
      RECT 81.085 2.395 81.255 3.865 ;
      RECT 81.085 5.015 81.255 6.485 ;
      RECT 81.085 7.795 81.255 8.305 ;
      RECT 80.095 0.575 80.265 1.085 ;
      RECT 80.095 2.395 80.265 3.865 ;
      RECT 80.095 5.015 80.265 6.485 ;
      RECT 80.095 7.795 80.265 8.305 ;
      RECT 78.73 0.575 78.9 3.865 ;
      RECT 78.73 5.015 78.9 8.305 ;
      RECT 78.3 0.575 78.47 1.085 ;
      RECT 78.3 1.655 78.47 3.865 ;
      RECT 78.3 5.015 78.47 7.225 ;
      RECT 78.3 7.795 78.47 8.305 ;
      RECT 76.93 1.66 77.1 2.935 ;
      RECT 76.93 5.945 77.1 7.22 ;
      RECT 74.41 2.495 74.58 2.825 ;
      RECT 73.69 1.755 73.86 2.105 ;
      RECT 73.69 3.485 73.86 3.815 ;
      RECT 72.69 3.485 72.86 3.815 ;
      RECT 72.45 2.495 72.62 2.945 ;
      RECT 71.97 2.495 72.14 2.825 ;
      RECT 71.25 1.755 71.42 2.105 ;
      RECT 70.25 3.145 70.42 3.505 ;
      RECT 70.01 2.495 70.18 2.945 ;
      RECT 69.53 2.495 69.7 2.825 ;
      RECT 69.29 1.755 69.46 2.105 ;
      RECT 68.81 3.055 68.98 3.475 ;
      RECT 67.81 1.755 67.98 2.105 ;
      RECT 67.57 2.495 67.74 2.825 ;
      RECT 66.85 1.755 67.02 2.105 ;
      RECT 66.37 3.055 66.54 3.475 ;
      RECT 64.76 0.575 64.93 1.085 ;
      RECT 64.76 2.395 64.93 3.865 ;
      RECT 64.76 5.015 64.93 6.485 ;
      RECT 64.76 7.795 64.93 8.305 ;
      RECT 63.77 0.575 63.94 1.085 ;
      RECT 63.77 2.395 63.94 3.865 ;
      RECT 63.77 5.015 63.94 6.485 ;
      RECT 63.77 7.795 63.94 8.305 ;
      RECT 62.405 0.575 62.575 3.865 ;
      RECT 62.405 5.015 62.575 8.305 ;
      RECT 61.975 0.575 62.145 1.085 ;
      RECT 61.975 1.655 62.145 3.865 ;
      RECT 61.975 5.015 62.145 7.225 ;
      RECT 61.975 7.795 62.145 8.305 ;
      RECT 60.605 1.66 60.775 2.935 ;
      RECT 60.605 5.945 60.775 7.22 ;
      RECT 58.085 2.495 58.255 2.825 ;
      RECT 57.365 1.755 57.535 2.105 ;
      RECT 57.365 3.485 57.535 3.815 ;
      RECT 56.365 3.485 56.535 3.815 ;
      RECT 56.125 2.495 56.295 2.945 ;
      RECT 55.645 2.495 55.815 2.825 ;
      RECT 54.925 1.755 55.095 2.105 ;
      RECT 53.925 3.145 54.095 3.505 ;
      RECT 53.685 2.495 53.855 2.945 ;
      RECT 53.205 2.495 53.375 2.825 ;
      RECT 52.965 1.755 53.135 2.105 ;
      RECT 52.485 3.055 52.655 3.475 ;
      RECT 51.485 1.755 51.655 2.105 ;
      RECT 51.245 2.495 51.415 2.825 ;
      RECT 50.525 1.755 50.695 2.105 ;
      RECT 50.045 3.055 50.215 3.475 ;
      RECT 48.44 0.575 48.61 1.085 ;
      RECT 48.44 2.395 48.61 3.865 ;
      RECT 48.44 5.015 48.61 6.485 ;
      RECT 48.44 7.795 48.61 8.305 ;
      RECT 47.45 0.575 47.62 1.085 ;
      RECT 47.45 2.395 47.62 3.865 ;
      RECT 47.45 5.015 47.62 6.485 ;
      RECT 47.45 7.795 47.62 8.305 ;
      RECT 46.085 0.575 46.255 3.865 ;
      RECT 46.085 5.015 46.255 8.305 ;
      RECT 45.655 0.575 45.825 1.085 ;
      RECT 45.655 1.655 45.825 3.865 ;
      RECT 45.655 5.015 45.825 7.225 ;
      RECT 45.655 7.795 45.825 8.305 ;
      RECT 44.285 1.66 44.455 2.935 ;
      RECT 44.285 5.945 44.455 7.22 ;
      RECT 41.765 2.495 41.935 2.825 ;
      RECT 41.045 1.755 41.215 2.105 ;
      RECT 41.045 3.485 41.215 3.815 ;
      RECT 40.045 3.485 40.215 3.815 ;
      RECT 39.805 2.495 39.975 2.945 ;
      RECT 39.325 2.495 39.495 2.825 ;
      RECT 38.605 1.755 38.775 2.105 ;
      RECT 37.605 3.145 37.775 3.505 ;
      RECT 37.365 2.495 37.535 2.945 ;
      RECT 36.885 2.495 37.055 2.825 ;
      RECT 36.645 1.755 36.815 2.105 ;
      RECT 36.165 3.055 36.335 3.475 ;
      RECT 35.165 1.755 35.335 2.105 ;
      RECT 34.925 2.495 35.095 2.825 ;
      RECT 34.205 1.755 34.375 2.105 ;
      RECT 33.725 3.055 33.895 3.475 ;
      RECT 32.115 0.575 32.285 1.085 ;
      RECT 32.115 2.395 32.285 3.865 ;
      RECT 32.115 5.015 32.285 6.485 ;
      RECT 32.115 7.795 32.285 8.305 ;
      RECT 31.125 0.575 31.295 1.085 ;
      RECT 31.125 2.395 31.295 3.865 ;
      RECT 31.125 5.015 31.295 6.485 ;
      RECT 31.125 7.795 31.295 8.305 ;
      RECT 29.76 0.575 29.93 3.865 ;
      RECT 29.76 5.015 29.93 8.305 ;
      RECT 29.33 0.575 29.5 1.085 ;
      RECT 29.33 1.655 29.5 3.865 ;
      RECT 29.33 5.015 29.5 7.225 ;
      RECT 29.33 7.795 29.5 8.305 ;
      RECT 27.96 1.66 28.13 2.935 ;
      RECT 27.96 5.945 28.13 7.22 ;
      RECT 25.44 2.495 25.61 2.825 ;
      RECT 24.72 1.755 24.89 2.105 ;
      RECT 24.72 3.485 24.89 3.815 ;
      RECT 23.72 3.485 23.89 3.815 ;
      RECT 23.48 2.495 23.65 2.945 ;
      RECT 23 2.495 23.17 2.825 ;
      RECT 22.28 1.755 22.45 2.105 ;
      RECT 21.28 3.145 21.45 3.505 ;
      RECT 21.04 2.495 21.21 2.945 ;
      RECT 20.56 2.495 20.73 2.825 ;
      RECT 20.32 1.755 20.49 2.105 ;
      RECT 19.84 3.055 20.01 3.475 ;
      RECT 18.84 1.755 19.01 2.105 ;
      RECT 18.6 2.495 18.77 2.825 ;
      RECT 17.88 1.755 18.05 2.105 ;
      RECT 17.4 3.055 17.57 3.475 ;
      RECT 15.795 0.575 15.965 1.085 ;
      RECT 15.795 2.395 15.965 3.865 ;
      RECT 15.795 5.015 15.965 6.485 ;
      RECT 15.795 7.795 15.965 8.305 ;
      RECT 14.805 0.575 14.975 1.085 ;
      RECT 14.805 2.395 14.975 3.865 ;
      RECT 14.805 5.015 14.975 6.485 ;
      RECT 14.805 7.795 14.975 8.305 ;
      RECT 13.44 0.575 13.61 3.865 ;
      RECT 13.44 5.015 13.61 8.305 ;
      RECT 13.01 0.575 13.18 1.085 ;
      RECT 13.01 1.655 13.18 3.865 ;
      RECT 13.01 5.015 13.18 7.225 ;
      RECT 13.01 7.795 13.18 8.305 ;
      RECT 11.64 1.66 11.81 2.935 ;
      RECT 11.64 5.945 11.81 7.22 ;
      RECT 9.12 2.495 9.29 2.825 ;
      RECT 8.4 1.755 8.57 2.105 ;
      RECT 8.4 3.485 8.57 3.815 ;
      RECT 7.4 3.485 7.57 3.815 ;
      RECT 7.16 2.495 7.33 2.945 ;
      RECT 6.68 2.495 6.85 2.825 ;
      RECT 5.96 1.755 6.13 2.105 ;
      RECT 4.96 3.145 5.13 3.505 ;
      RECT 4.72 2.495 4.89 2.945 ;
      RECT 4.24 2.495 4.41 2.825 ;
      RECT 4 1.755 4.17 2.105 ;
      RECT 3.52 3.055 3.69 3.475 ;
      RECT 2.52 1.755 2.69 2.105 ;
      RECT 2.28 2.495 2.45 2.825 ;
      RECT 1.56 1.755 1.73 2.105 ;
      RECT 1.08 3.055 1.25 3.475 ;
  END
END sky130_osu_ring_oscillator_mpr2ea_8

MACRO sky130_osu_ring_oscillator_mpr2et_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2et_8 0 0 ;
  SIZE 92.805 BY 8.88 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT 84.295 3.535 84.85 3.865 ;
      RECT 84.295 1.87 84.595 3.865 ;
      RECT 80.36 2.975 80.915 3.305 ;
      RECT 80.615 1.87 80.915 3.305 ;
      RECT 80.615 1.87 84.595 2.17 ;
      RECT 65.735 3.535 66.29 3.865 ;
      RECT 65.735 1.87 66.035 3.865 ;
      RECT 61.8 2.975 62.355 3.305 ;
      RECT 62.055 1.87 62.355 3.305 ;
      RECT 62.055 1.87 66.035 2.17 ;
      RECT 47.175 3.535 47.73 3.865 ;
      RECT 47.175 1.87 47.475 3.865 ;
      RECT 43.24 2.975 43.795 3.305 ;
      RECT 43.495 1.87 43.795 3.305 ;
      RECT 43.495 1.87 47.475 2.17 ;
      RECT 28.615 3.535 29.17 3.865 ;
      RECT 28.615 1.87 28.915 3.865 ;
      RECT 24.68 2.975 25.235 3.305 ;
      RECT 24.935 1.87 25.235 3.305 ;
      RECT 24.935 1.87 28.915 2.17 ;
      RECT 10.055 3.535 10.61 3.865 ;
      RECT 10.055 1.87 10.355 3.865 ;
      RECT 6.12 2.975 6.675 3.305 ;
      RECT 6.375 1.87 6.675 3.305 ;
      RECT 6.375 1.87 10.355 2.17 ;
      RECT 85.48 1.855 86.21 2.185 ;
      RECT 83.26 3.535 83.99 3.865 ;
      RECT 81.56 3.535 82.29 3.865 ;
      RECT 79.12 2.415 79.85 2.745 ;
      RECT 77.68 2.975 78.41 3.305 ;
      RECT 76.605 2.415 77.335 2.745 ;
      RECT 75.57 2.415 76.3 2.745 ;
      RECT 75.24 3.535 75.97 3.865 ;
      RECT 66.92 1.855 67.65 2.185 ;
      RECT 64.7 3.535 65.43 3.865 ;
      RECT 63 3.535 63.73 3.865 ;
      RECT 60.56 2.415 61.29 2.745 ;
      RECT 59.12 2.975 59.85 3.305 ;
      RECT 58.045 2.415 58.775 2.745 ;
      RECT 57.01 2.415 57.74 2.745 ;
      RECT 56.68 3.535 57.41 3.865 ;
      RECT 48.36 1.855 49.09 2.185 ;
      RECT 46.14 3.535 46.87 3.865 ;
      RECT 44.44 3.535 45.17 3.865 ;
      RECT 42 2.415 42.73 2.745 ;
      RECT 40.56 2.975 41.29 3.305 ;
      RECT 39.485 2.415 40.215 2.745 ;
      RECT 38.45 2.415 39.18 2.745 ;
      RECT 38.12 3.535 38.85 3.865 ;
      RECT 29.8 1.855 30.53 2.185 ;
      RECT 27.58 3.535 28.31 3.865 ;
      RECT 25.88 3.535 26.61 3.865 ;
      RECT 23.44 2.415 24.17 2.745 ;
      RECT 22 2.975 22.73 3.305 ;
      RECT 20.925 2.415 21.655 2.745 ;
      RECT 19.89 2.415 20.62 2.745 ;
      RECT 19.56 3.535 20.29 3.865 ;
      RECT 11.24 1.855 11.97 2.185 ;
      RECT 9.02 3.535 9.75 3.865 ;
      RECT 7.32 3.535 8.05 3.865 ;
      RECT 4.88 2.415 5.61 2.745 ;
      RECT 3.44 2.975 4.17 3.305 ;
      RECT 2.365 2.415 3.095 2.745 ;
      RECT 1.33 2.415 2.06 2.745 ;
      RECT 1 3.535 1.73 3.865 ;
    LAYER via2 ;
      RECT 85.545 1.92 85.745 2.12 ;
      RECT 84.585 3.6 84.785 3.8 ;
      RECT 83.585 3.6 83.785 3.8 ;
      RECT 81.625 3.6 81.825 3.8 ;
      RECT 80.425 3.04 80.625 3.24 ;
      RECT 79.185 2.48 79.385 2.68 ;
      RECT 77.745 3.04 77.945 3.24 ;
      RECT 77.005 2.48 77.205 2.68 ;
      RECT 75.785 2.48 75.985 2.68 ;
      RECT 75.305 3.6 75.505 3.8 ;
      RECT 66.985 1.92 67.185 2.12 ;
      RECT 66.025 3.6 66.225 3.8 ;
      RECT 65.025 3.6 65.225 3.8 ;
      RECT 63.065 3.6 63.265 3.8 ;
      RECT 61.865 3.04 62.065 3.24 ;
      RECT 60.625 2.48 60.825 2.68 ;
      RECT 59.185 3.04 59.385 3.24 ;
      RECT 58.445 2.48 58.645 2.68 ;
      RECT 57.225 2.48 57.425 2.68 ;
      RECT 56.745 3.6 56.945 3.8 ;
      RECT 48.425 1.92 48.625 2.12 ;
      RECT 47.465 3.6 47.665 3.8 ;
      RECT 46.465 3.6 46.665 3.8 ;
      RECT 44.505 3.6 44.705 3.8 ;
      RECT 43.305 3.04 43.505 3.24 ;
      RECT 42.065 2.48 42.265 2.68 ;
      RECT 40.625 3.04 40.825 3.24 ;
      RECT 39.885 2.48 40.085 2.68 ;
      RECT 38.665 2.48 38.865 2.68 ;
      RECT 38.185 3.6 38.385 3.8 ;
      RECT 29.865 1.92 30.065 2.12 ;
      RECT 28.905 3.6 29.105 3.8 ;
      RECT 27.905 3.6 28.105 3.8 ;
      RECT 25.945 3.6 26.145 3.8 ;
      RECT 24.745 3.04 24.945 3.24 ;
      RECT 23.505 2.48 23.705 2.68 ;
      RECT 22.065 3.04 22.265 3.24 ;
      RECT 21.325 2.48 21.525 2.68 ;
      RECT 20.105 2.48 20.305 2.68 ;
      RECT 19.625 3.6 19.825 3.8 ;
      RECT 11.305 1.92 11.505 2.12 ;
      RECT 10.345 3.6 10.545 3.8 ;
      RECT 9.345 3.6 9.545 3.8 ;
      RECT 7.385 3.6 7.585 3.8 ;
      RECT 6.185 3.04 6.385 3.24 ;
      RECT 4.945 2.48 5.145 2.68 ;
      RECT 3.505 3.04 3.705 3.24 ;
      RECT 2.765 2.48 2.965 2.68 ;
      RECT 1.545 2.48 1.745 2.68 ;
      RECT 1.065 3.6 1.265 3.8 ;
    LAYER met2 ;
      RECT 14.835 6.28 15.155 6.605 ;
      RECT 14.865 5.695 15.035 6.605 ;
      RECT 14.865 5.695 15.04 6.045 ;
      RECT 14.865 5.695 15.84 5.87 ;
      RECT 15.665 1.965 15.84 5.87 ;
      RECT 2.475 2.98 2.735 3.3 ;
      RECT 2.415 2.51 2.555 3.21 ;
      RECT 2.725 2.395 3.005 2.765 ;
      RECT 4.195 2.42 4.455 2.74 ;
      RECT 2.415 2.51 4.455 2.65 ;
      RECT 2.82 1.32 2.99 2.765 ;
      RECT 15.61 1.965 15.96 2.315 ;
      RECT 13.555 2.04 15.96 2.195 ;
      RECT 13.565 2.025 15.96 2.195 ;
      RECT 13.565 0.215 13.735 2.195 ;
      RECT 2.82 1.32 13.735 1.49 ;
      RECT 92.235 1.095 92.575 1.445 ;
      RECT 92.235 1.17 92.58 1.36 ;
      RECT 92.265 0.215 92.435 1.445 ;
      RECT 13.565 0.215 92.435 0.385 ;
      RECT 89.075 6.28 89.395 6.605 ;
      RECT 89.105 5.695 89.275 6.605 ;
      RECT 89.105 5.695 89.28 6.045 ;
      RECT 89.105 5.695 90.08 5.87 ;
      RECT 89.905 1.965 90.08 5.87 ;
      RECT 76.715 2.98 76.975 3.3 ;
      RECT 76.655 2.51 76.795 3.21 ;
      RECT 76.965 2.395 77.245 2.765 ;
      RECT 78.435 2.42 78.695 2.74 ;
      RECT 76.655 2.51 78.695 2.65 ;
      RECT 77.06 1.32 77.23 2.765 ;
      RECT 89.85 1.965 90.2 2.315 ;
      RECT 87.795 2.04 90.2 2.195 ;
      RECT 87.805 2.025 90.2 2.195 ;
      RECT 87.805 1.32 87.975 2.195 ;
      RECT 74.775 1.4 77.23 1.59 ;
      RECT 77.06 1.32 87.975 1.49 ;
      RECT 73.675 1.095 74.015 1.445 ;
      RECT 74.775 1.17 74.965 1.59 ;
      RECT 73.675 1.17 74.965 1.36 ;
      RECT 89.875 6.655 90.2 6.98 ;
      RECT 88.76 6.745 90.2 6.915 ;
      RECT 88.76 2.395 88.92 6.915 ;
      RECT 89.075 2.365 89.395 2.685 ;
      RECT 88.76 2.395 89.395 2.565 ;
      RECT 88.025 5.845 88.365 6.195 ;
      RECT 88.11 2.705 88.28 6.195 ;
      RECT 88.035 2.705 88.375 3.055 ;
      RECT 81.62 4.135 87.73 4.325 ;
      RECT 87.56 3.145 87.73 4.325 ;
      RECT 87.54 3.15 87.73 4.325 ;
      RECT 81.62 3.515 81.81 4.325 ;
      RECT 81.585 3.515 81.865 3.885 ;
      RECT 81.655 3.07 81.795 4.325 ;
      RECT 87.47 3.15 87.81 3.5 ;
      RECT 81.465 2.955 81.745 3.325 ;
      RECT 81.175 3.07 81.795 3.21 ;
      RECT 81.175 1.86 81.315 3.21 ;
      RECT 81.115 1.86 81.375 2.18 ;
      RECT 84.075 2.98 84.335 3.3 ;
      RECT 84.135 1.86 84.275 3.3 ;
      RECT 84.075 1.86 84.335 2.18 ;
      RECT 83.075 3.54 83.335 3.86 ;
      RECT 83.075 2.955 83.275 3.86 ;
      RECT 83.015 1.86 83.155 3.49 ;
      RECT 83.015 2.955 83.515 3.325 ;
      RECT 82.955 1.86 83.215 2.18 ;
      RECT 82.595 3.54 82.855 3.86 ;
      RECT 82.655 1.95 82.795 3.86 ;
      RECT 82.355 1.95 82.795 2.18 ;
      RECT 82.355 1.86 82.615 2.18 ;
      RECT 82.115 2.42 82.375 2.74 ;
      RECT 81.535 2.51 82.375 2.65 ;
      RECT 81.535 1.57 81.675 2.65 ;
      RECT 78.195 1.86 78.455 2.18 ;
      RECT 78.195 1.95 79.235 2.09 ;
      RECT 79.095 1.57 79.235 2.09 ;
      RECT 79.095 1.57 81.675 1.71 ;
      RECT 80.385 2.955 80.665 3.325 ;
      RECT 80.455 1.86 80.595 3.325 ;
      RECT 80.395 1.86 80.655 2.18 ;
      RECT 80.035 3.54 80.295 3.86 ;
      RECT 80.095 1.95 80.235 3.86 ;
      RECT 79.675 1.86 79.935 2.18 ;
      RECT 79.675 1.95 80.235 2.09 ;
      RECT 77.705 2.955 77.985 3.325 ;
      RECT 79.675 2.98 79.935 3.3 ;
      RECT 77.355 2.98 77.985 3.3 ;
      RECT 77.355 3.07 79.935 3.21 ;
      RECT 79.145 2.395 79.425 2.765 ;
      RECT 79.145 2.42 79.675 2.74 ;
      RECT 76.235 2.98 76.495 3.3 ;
      RECT 76.295 1.86 76.435 3.3 ;
      RECT 76.235 1.86 76.495 2.18 ;
      RECT 75.265 3.515 75.545 3.885 ;
      RECT 75.275 3.26 75.535 3.885 ;
      RECT 70.515 6.28 70.835 6.605 ;
      RECT 70.545 5.695 70.715 6.605 ;
      RECT 70.545 5.695 70.72 6.045 ;
      RECT 70.545 5.695 71.52 5.87 ;
      RECT 71.345 1.965 71.52 5.87 ;
      RECT 58.155 2.98 58.415 3.3 ;
      RECT 58.095 2.51 58.235 3.21 ;
      RECT 58.405 2.395 58.685 2.765 ;
      RECT 59.875 2.42 60.135 2.74 ;
      RECT 58.095 2.51 60.135 2.65 ;
      RECT 58.5 1.32 58.67 2.765 ;
      RECT 71.29 1.965 71.64 2.315 ;
      RECT 69.235 2.04 71.64 2.195 ;
      RECT 69.245 2.025 71.64 2.195 ;
      RECT 69.245 1.32 69.415 2.195 ;
      RECT 56.105 1.385 58.67 1.575 ;
      RECT 58.5 1.32 69.415 1.49 ;
      RECT 55.115 1.095 55.455 1.445 ;
      RECT 56.105 1.17 56.295 1.575 ;
      RECT 55.115 1.17 56.295 1.36 ;
      RECT 71.315 6.655 71.64 6.98 ;
      RECT 70.2 6.745 71.64 6.915 ;
      RECT 70.2 2.395 70.36 6.915 ;
      RECT 70.515 2.365 70.835 2.685 ;
      RECT 70.2 2.395 70.835 2.565 ;
      RECT 69.465 5.845 69.805 6.195 ;
      RECT 69.55 2.705 69.72 6.195 ;
      RECT 69.475 2.705 69.815 3.055 ;
      RECT 63.06 4.135 69.17 4.325 ;
      RECT 69 3.145 69.17 4.325 ;
      RECT 68.98 3.15 69.17 4.325 ;
      RECT 63.06 3.515 63.25 4.325 ;
      RECT 63.025 3.515 63.305 3.885 ;
      RECT 63.095 3.07 63.235 4.325 ;
      RECT 68.91 3.15 69.25 3.5 ;
      RECT 62.905 2.955 63.185 3.325 ;
      RECT 62.615 3.07 63.235 3.21 ;
      RECT 62.615 1.86 62.755 3.21 ;
      RECT 62.555 1.86 62.815 2.18 ;
      RECT 65.515 2.98 65.775 3.3 ;
      RECT 65.575 1.86 65.715 3.3 ;
      RECT 65.515 1.86 65.775 2.18 ;
      RECT 64.515 3.54 64.775 3.86 ;
      RECT 64.515 2.955 64.715 3.86 ;
      RECT 64.455 1.86 64.595 3.49 ;
      RECT 64.455 2.955 64.955 3.325 ;
      RECT 64.395 1.86 64.655 2.18 ;
      RECT 64.035 3.54 64.295 3.86 ;
      RECT 64.095 1.95 64.235 3.86 ;
      RECT 63.795 1.95 64.235 2.18 ;
      RECT 63.795 1.86 64.055 2.18 ;
      RECT 63.555 2.42 63.815 2.74 ;
      RECT 62.975 2.51 63.815 2.65 ;
      RECT 62.975 1.57 63.115 2.65 ;
      RECT 59.635 1.86 59.895 2.18 ;
      RECT 59.635 1.95 60.675 2.09 ;
      RECT 60.535 1.57 60.675 2.09 ;
      RECT 60.535 1.57 63.115 1.71 ;
      RECT 61.825 2.955 62.105 3.325 ;
      RECT 61.895 1.86 62.035 3.325 ;
      RECT 61.835 1.86 62.095 2.18 ;
      RECT 61.475 3.54 61.735 3.86 ;
      RECT 61.535 1.95 61.675 3.86 ;
      RECT 61.115 1.86 61.375 2.18 ;
      RECT 61.115 1.95 61.675 2.09 ;
      RECT 59.145 2.955 59.425 3.325 ;
      RECT 61.115 2.98 61.375 3.3 ;
      RECT 58.795 2.98 59.425 3.3 ;
      RECT 58.795 3.07 61.375 3.21 ;
      RECT 60.585 2.395 60.865 2.765 ;
      RECT 60.585 2.42 61.115 2.74 ;
      RECT 57.675 2.98 57.935 3.3 ;
      RECT 57.735 1.86 57.875 3.3 ;
      RECT 57.675 1.86 57.935 2.18 ;
      RECT 56.705 3.515 56.985 3.885 ;
      RECT 56.715 3.26 56.975 3.885 ;
      RECT 51.955 6.28 52.275 6.605 ;
      RECT 51.985 5.695 52.155 6.605 ;
      RECT 51.985 5.695 52.16 6.045 ;
      RECT 51.985 5.695 52.96 5.87 ;
      RECT 52.785 1.965 52.96 5.87 ;
      RECT 39.595 2.98 39.855 3.3 ;
      RECT 39.535 2.51 39.675 3.21 ;
      RECT 39.845 2.395 40.125 2.765 ;
      RECT 41.315 2.42 41.575 2.74 ;
      RECT 39.535 2.51 41.575 2.65 ;
      RECT 39.94 1.32 40.11 2.765 ;
      RECT 52.73 1.965 53.08 2.315 ;
      RECT 50.675 2.04 53.08 2.195 ;
      RECT 50.685 2.025 53.08 2.195 ;
      RECT 50.685 1.32 50.855 2.195 ;
      RECT 37.575 1.37 40.11 1.56 ;
      RECT 39.94 1.32 50.855 1.49 ;
      RECT 36.565 1.095 36.905 1.445 ;
      RECT 37.575 1.17 37.765 1.56 ;
      RECT 36.565 1.17 37.765 1.36 ;
      RECT 52.755 6.655 53.08 6.98 ;
      RECT 51.64 6.745 53.08 6.915 ;
      RECT 51.64 2.395 51.8 6.915 ;
      RECT 51.955 2.365 52.275 2.685 ;
      RECT 51.64 2.395 52.275 2.565 ;
      RECT 50.905 5.845 51.245 6.195 ;
      RECT 50.99 2.705 51.16 6.195 ;
      RECT 50.915 2.705 51.255 3.055 ;
      RECT 44.5 4.135 50.61 4.325 ;
      RECT 50.44 3.145 50.61 4.325 ;
      RECT 50.42 3.15 50.61 4.325 ;
      RECT 44.5 3.515 44.69 4.325 ;
      RECT 44.465 3.515 44.745 3.885 ;
      RECT 44.535 3.07 44.675 4.325 ;
      RECT 50.35 3.15 50.69 3.5 ;
      RECT 44.345 2.955 44.625 3.325 ;
      RECT 44.055 3.07 44.675 3.21 ;
      RECT 44.055 1.86 44.195 3.21 ;
      RECT 43.995 1.86 44.255 2.18 ;
      RECT 46.955 2.98 47.215 3.3 ;
      RECT 47.015 1.86 47.155 3.3 ;
      RECT 46.955 1.86 47.215 2.18 ;
      RECT 45.955 3.54 46.215 3.86 ;
      RECT 45.955 2.955 46.155 3.86 ;
      RECT 45.895 1.86 46.035 3.49 ;
      RECT 45.895 2.955 46.395 3.325 ;
      RECT 45.835 1.86 46.095 2.18 ;
      RECT 45.475 3.54 45.735 3.86 ;
      RECT 45.535 1.95 45.675 3.86 ;
      RECT 45.235 1.95 45.675 2.18 ;
      RECT 45.235 1.86 45.495 2.18 ;
      RECT 44.995 2.42 45.255 2.74 ;
      RECT 44.415 2.51 45.255 2.65 ;
      RECT 44.415 1.57 44.555 2.65 ;
      RECT 41.075 1.86 41.335 2.18 ;
      RECT 41.075 1.95 42.115 2.09 ;
      RECT 41.975 1.57 42.115 2.09 ;
      RECT 41.975 1.57 44.555 1.71 ;
      RECT 43.265 2.955 43.545 3.325 ;
      RECT 43.335 1.86 43.475 3.325 ;
      RECT 43.275 1.86 43.535 2.18 ;
      RECT 42.915 3.54 43.175 3.86 ;
      RECT 42.975 1.95 43.115 3.86 ;
      RECT 42.555 1.86 42.815 2.18 ;
      RECT 42.555 1.95 43.115 2.09 ;
      RECT 40.585 2.955 40.865 3.325 ;
      RECT 42.555 2.98 42.815 3.3 ;
      RECT 40.235 2.98 40.865 3.3 ;
      RECT 40.235 3.07 42.815 3.21 ;
      RECT 42.025 2.395 42.305 2.765 ;
      RECT 42.025 2.42 42.555 2.74 ;
      RECT 39.115 2.98 39.375 3.3 ;
      RECT 39.175 1.86 39.315 3.3 ;
      RECT 39.115 1.86 39.375 2.18 ;
      RECT 38.145 3.515 38.425 3.885 ;
      RECT 38.155 3.26 38.415 3.885 ;
      RECT 33.395 6.28 33.715 6.605 ;
      RECT 33.425 5.695 33.595 6.605 ;
      RECT 33.425 5.695 33.6 6.045 ;
      RECT 33.425 5.695 34.4 5.87 ;
      RECT 34.225 1.965 34.4 5.87 ;
      RECT 21.035 2.98 21.295 3.3 ;
      RECT 20.975 2.51 21.115 3.21 ;
      RECT 21.285 2.395 21.565 2.765 ;
      RECT 22.755 2.42 23.015 2.74 ;
      RECT 20.975 2.51 23.015 2.65 ;
      RECT 21.38 1.32 21.55 2.765 ;
      RECT 34.17 1.965 34.52 2.315 ;
      RECT 32.115 2.04 34.52 2.195 ;
      RECT 32.125 2.025 34.52 2.195 ;
      RECT 32.125 1.32 32.295 2.195 ;
      RECT 18.98 1.34 21.55 1.53 ;
      RECT 21.38 1.32 32.295 1.49 ;
      RECT 17.995 1.095 18.335 1.445 ;
      RECT 17.995 1.17 19.17 1.36 ;
      RECT 34.195 6.655 34.52 6.98 ;
      RECT 33.08 6.745 34.52 6.915 ;
      RECT 33.08 2.395 33.24 6.915 ;
      RECT 33.395 2.365 33.715 2.685 ;
      RECT 33.08 2.395 33.715 2.565 ;
      RECT 32.345 5.845 32.685 6.195 ;
      RECT 32.43 2.705 32.6 6.195 ;
      RECT 32.355 2.705 32.695 3.055 ;
      RECT 25.94 4.135 32.05 4.325 ;
      RECT 31.88 3.145 32.05 4.325 ;
      RECT 31.86 3.15 32.05 4.325 ;
      RECT 25.94 3.515 26.13 4.325 ;
      RECT 25.905 3.515 26.185 3.885 ;
      RECT 25.975 3.07 26.115 4.325 ;
      RECT 31.79 3.15 32.13 3.5 ;
      RECT 25.785 2.955 26.065 3.325 ;
      RECT 25.495 3.07 26.115 3.21 ;
      RECT 25.495 1.86 25.635 3.21 ;
      RECT 25.435 1.86 25.695 2.18 ;
      RECT 28.395 2.98 28.655 3.3 ;
      RECT 28.455 1.86 28.595 3.3 ;
      RECT 28.395 1.86 28.655 2.18 ;
      RECT 27.395 3.54 27.655 3.86 ;
      RECT 27.395 2.955 27.595 3.86 ;
      RECT 27.335 1.86 27.475 3.49 ;
      RECT 27.335 2.955 27.835 3.325 ;
      RECT 27.275 1.86 27.535 2.18 ;
      RECT 26.915 3.54 27.175 3.86 ;
      RECT 26.975 1.95 27.115 3.86 ;
      RECT 26.675 1.95 27.115 2.18 ;
      RECT 26.675 1.86 26.935 2.18 ;
      RECT 26.435 2.42 26.695 2.74 ;
      RECT 25.855 2.51 26.695 2.65 ;
      RECT 25.855 1.57 25.995 2.65 ;
      RECT 22.515 1.86 22.775 2.18 ;
      RECT 22.515 1.95 23.555 2.09 ;
      RECT 23.415 1.57 23.555 2.09 ;
      RECT 23.415 1.57 25.995 1.71 ;
      RECT 24.705 2.955 24.985 3.325 ;
      RECT 24.775 1.86 24.915 3.325 ;
      RECT 24.715 1.86 24.975 2.18 ;
      RECT 24.355 3.54 24.615 3.86 ;
      RECT 24.415 1.95 24.555 3.86 ;
      RECT 23.995 1.86 24.255 2.18 ;
      RECT 23.995 1.95 24.555 2.09 ;
      RECT 22.025 2.955 22.305 3.325 ;
      RECT 23.995 2.98 24.255 3.3 ;
      RECT 21.675 2.98 22.305 3.3 ;
      RECT 21.675 3.07 24.255 3.21 ;
      RECT 23.465 2.395 23.745 2.765 ;
      RECT 23.465 2.42 23.995 2.74 ;
      RECT 20.555 2.98 20.815 3.3 ;
      RECT 20.615 1.86 20.755 3.3 ;
      RECT 20.555 1.86 20.815 2.18 ;
      RECT 19.585 3.515 19.865 3.885 ;
      RECT 19.595 3.26 19.855 3.885 ;
      RECT 15.635 6.655 15.96 6.98 ;
      RECT 14.52 6.745 15.96 6.915 ;
      RECT 14.52 2.395 14.68 6.915 ;
      RECT 14.835 2.365 15.155 2.685 ;
      RECT 14.52 2.395 15.155 2.565 ;
      RECT 13.785 5.845 14.125 6.195 ;
      RECT 13.87 2.705 14.04 6.195 ;
      RECT 13.795 2.705 14.135 3.055 ;
      RECT 7.38 4.135 13.49 4.325 ;
      RECT 13.32 3.145 13.49 4.325 ;
      RECT 13.3 3.15 13.49 4.325 ;
      RECT 7.38 3.515 7.57 4.325 ;
      RECT 7.345 3.515 7.625 3.885 ;
      RECT 7.415 3.07 7.555 4.325 ;
      RECT 13.23 3.15 13.57 3.5 ;
      RECT 7.225 2.955 7.505 3.325 ;
      RECT 6.935 3.07 7.555 3.21 ;
      RECT 6.935 1.86 7.075 3.21 ;
      RECT 6.875 1.86 7.135 2.18 ;
      RECT 9.835 2.98 10.095 3.3 ;
      RECT 9.895 1.86 10.035 3.3 ;
      RECT 9.835 1.86 10.095 2.18 ;
      RECT 8.835 3.54 9.095 3.86 ;
      RECT 8.835 2.955 9.035 3.86 ;
      RECT 8.775 1.86 8.915 3.49 ;
      RECT 8.775 2.955 9.275 3.325 ;
      RECT 8.715 1.86 8.975 2.18 ;
      RECT 8.355 3.54 8.615 3.86 ;
      RECT 8.415 1.95 8.555 3.86 ;
      RECT 8.115 1.95 8.555 2.18 ;
      RECT 8.115 1.86 8.375 2.18 ;
      RECT 7.875 2.42 8.135 2.74 ;
      RECT 7.295 2.51 8.135 2.65 ;
      RECT 7.295 1.57 7.435 2.65 ;
      RECT 3.955 1.86 4.215 2.18 ;
      RECT 3.955 1.95 4.995 2.09 ;
      RECT 4.855 1.57 4.995 2.09 ;
      RECT 4.855 1.57 7.435 1.71 ;
      RECT 6.145 2.955 6.425 3.325 ;
      RECT 6.215 1.86 6.355 3.325 ;
      RECT 6.155 1.86 6.415 2.18 ;
      RECT 5.795 3.54 6.055 3.86 ;
      RECT 5.855 1.95 5.995 3.86 ;
      RECT 5.435 1.86 5.695 2.18 ;
      RECT 5.435 1.95 5.995 2.09 ;
      RECT 3.465 2.955 3.745 3.325 ;
      RECT 5.435 2.98 5.695 3.3 ;
      RECT 3.115 2.98 3.745 3.3 ;
      RECT 3.115 3.07 5.695 3.21 ;
      RECT 4.905 2.395 5.185 2.765 ;
      RECT 4.905 2.42 5.435 2.74 ;
      RECT 1.995 2.98 2.255 3.3 ;
      RECT 2.055 1.86 2.195 3.3 ;
      RECT 1.995 1.86 2.255 2.18 ;
      RECT 1.025 3.515 1.305 3.885 ;
      RECT 1.035 3.26 1.295 3.885 ;
      RECT 85.505 1.835 85.785 2.205 ;
      RECT 84.545 3.515 84.825 3.885 ;
      RECT 83.545 3.515 83.825 3.885 ;
      RECT 75.745 2.395 76.025 2.765 ;
      RECT 66.945 1.835 67.225 2.205 ;
      RECT 65.985 3.515 66.265 3.885 ;
      RECT 64.985 3.515 65.265 3.885 ;
      RECT 57.185 2.395 57.465 2.765 ;
      RECT 48.385 1.835 48.665 2.205 ;
      RECT 47.425 3.515 47.705 3.885 ;
      RECT 46.425 3.515 46.705 3.885 ;
      RECT 38.625 2.395 38.905 2.765 ;
      RECT 29.825 1.835 30.105 2.205 ;
      RECT 28.865 3.515 29.145 3.885 ;
      RECT 27.865 3.515 28.145 3.885 ;
      RECT 20.065 2.395 20.345 2.765 ;
      RECT 11.265 1.835 11.545 2.205 ;
      RECT 10.305 3.515 10.585 3.885 ;
      RECT 9.305 3.515 9.585 3.885 ;
      RECT 1.505 2.395 1.785 2.765 ;
    LAYER via1 ;
      RECT 92.335 1.195 92.485 1.345 ;
      RECT 89.965 6.74 90.115 6.89 ;
      RECT 89.95 2.065 90.1 2.215 ;
      RECT 89.16 2.45 89.31 2.6 ;
      RECT 89.16 6.37 89.31 6.52 ;
      RECT 88.135 2.805 88.285 2.955 ;
      RECT 88.125 5.945 88.275 6.095 ;
      RECT 87.57 3.25 87.72 3.4 ;
      RECT 85.57 1.945 85.72 2.095 ;
      RECT 84.61 3.625 84.76 3.775 ;
      RECT 84.13 1.945 84.28 2.095 ;
      RECT 84.13 3.065 84.28 3.215 ;
      RECT 83.61 3.625 83.76 3.775 ;
      RECT 83.13 3.625 83.28 3.775 ;
      RECT 83.01 1.945 83.16 2.095 ;
      RECT 82.65 3.625 82.8 3.775 ;
      RECT 82.41 1.945 82.56 2.095 ;
      RECT 82.17 2.505 82.32 2.655 ;
      RECT 81.65 3.625 81.8 3.775 ;
      RECT 81.17 1.945 81.32 2.095 ;
      RECT 80.45 1.945 80.6 2.095 ;
      RECT 80.45 3.065 80.6 3.215 ;
      RECT 80.09 3.625 80.24 3.775 ;
      RECT 79.73 1.945 79.88 2.095 ;
      RECT 79.73 3.065 79.88 3.215 ;
      RECT 79.47 2.505 79.62 2.655 ;
      RECT 78.49 2.505 78.64 2.655 ;
      RECT 78.25 1.945 78.4 2.095 ;
      RECT 77.41 3.065 77.56 3.215 ;
      RECT 76.77 3.065 76.92 3.215 ;
      RECT 76.29 1.945 76.44 2.095 ;
      RECT 76.29 3.065 76.44 3.215 ;
      RECT 75.81 2.505 75.96 2.655 ;
      RECT 75.33 3.345 75.48 3.495 ;
      RECT 73.775 1.195 73.925 1.345 ;
      RECT 71.405 6.74 71.555 6.89 ;
      RECT 71.39 2.065 71.54 2.215 ;
      RECT 70.6 2.45 70.75 2.6 ;
      RECT 70.6 6.37 70.75 6.52 ;
      RECT 69.575 2.805 69.725 2.955 ;
      RECT 69.565 5.945 69.715 6.095 ;
      RECT 69.01 3.25 69.16 3.4 ;
      RECT 67.01 1.945 67.16 2.095 ;
      RECT 66.05 3.625 66.2 3.775 ;
      RECT 65.57 1.945 65.72 2.095 ;
      RECT 65.57 3.065 65.72 3.215 ;
      RECT 65.05 3.625 65.2 3.775 ;
      RECT 64.57 3.625 64.72 3.775 ;
      RECT 64.45 1.945 64.6 2.095 ;
      RECT 64.09 3.625 64.24 3.775 ;
      RECT 63.85 1.945 64 2.095 ;
      RECT 63.61 2.505 63.76 2.655 ;
      RECT 63.09 3.625 63.24 3.775 ;
      RECT 62.61 1.945 62.76 2.095 ;
      RECT 61.89 1.945 62.04 2.095 ;
      RECT 61.89 3.065 62.04 3.215 ;
      RECT 61.53 3.625 61.68 3.775 ;
      RECT 61.17 1.945 61.32 2.095 ;
      RECT 61.17 3.065 61.32 3.215 ;
      RECT 60.91 2.505 61.06 2.655 ;
      RECT 59.93 2.505 60.08 2.655 ;
      RECT 59.69 1.945 59.84 2.095 ;
      RECT 58.85 3.065 59 3.215 ;
      RECT 58.21 3.065 58.36 3.215 ;
      RECT 57.73 1.945 57.88 2.095 ;
      RECT 57.73 3.065 57.88 3.215 ;
      RECT 57.25 2.505 57.4 2.655 ;
      RECT 56.77 3.345 56.92 3.495 ;
      RECT 55.215 1.195 55.365 1.345 ;
      RECT 52.845 6.74 52.995 6.89 ;
      RECT 52.83 2.065 52.98 2.215 ;
      RECT 52.04 2.45 52.19 2.6 ;
      RECT 52.04 6.37 52.19 6.52 ;
      RECT 51.015 2.805 51.165 2.955 ;
      RECT 51.005 5.945 51.155 6.095 ;
      RECT 50.45 3.25 50.6 3.4 ;
      RECT 48.45 1.945 48.6 2.095 ;
      RECT 47.49 3.625 47.64 3.775 ;
      RECT 47.01 1.945 47.16 2.095 ;
      RECT 47.01 3.065 47.16 3.215 ;
      RECT 46.49 3.625 46.64 3.775 ;
      RECT 46.01 3.625 46.16 3.775 ;
      RECT 45.89 1.945 46.04 2.095 ;
      RECT 45.53 3.625 45.68 3.775 ;
      RECT 45.29 1.945 45.44 2.095 ;
      RECT 45.05 2.505 45.2 2.655 ;
      RECT 44.53 3.625 44.68 3.775 ;
      RECT 44.05 1.945 44.2 2.095 ;
      RECT 43.33 1.945 43.48 2.095 ;
      RECT 43.33 3.065 43.48 3.215 ;
      RECT 42.97 3.625 43.12 3.775 ;
      RECT 42.61 1.945 42.76 2.095 ;
      RECT 42.61 3.065 42.76 3.215 ;
      RECT 42.35 2.505 42.5 2.655 ;
      RECT 41.37 2.505 41.52 2.655 ;
      RECT 41.13 1.945 41.28 2.095 ;
      RECT 40.29 3.065 40.44 3.215 ;
      RECT 39.65 3.065 39.8 3.215 ;
      RECT 39.17 1.945 39.32 2.095 ;
      RECT 39.17 3.065 39.32 3.215 ;
      RECT 38.69 2.505 38.84 2.655 ;
      RECT 38.21 3.345 38.36 3.495 ;
      RECT 36.665 1.195 36.815 1.345 ;
      RECT 34.285 6.74 34.435 6.89 ;
      RECT 34.27 2.065 34.42 2.215 ;
      RECT 33.48 2.45 33.63 2.6 ;
      RECT 33.48 6.37 33.63 6.52 ;
      RECT 32.455 2.805 32.605 2.955 ;
      RECT 32.445 5.945 32.595 6.095 ;
      RECT 31.89 3.25 32.04 3.4 ;
      RECT 29.89 1.945 30.04 2.095 ;
      RECT 28.93 3.625 29.08 3.775 ;
      RECT 28.45 1.945 28.6 2.095 ;
      RECT 28.45 3.065 28.6 3.215 ;
      RECT 27.93 3.625 28.08 3.775 ;
      RECT 27.45 3.625 27.6 3.775 ;
      RECT 27.33 1.945 27.48 2.095 ;
      RECT 26.97 3.625 27.12 3.775 ;
      RECT 26.73 1.945 26.88 2.095 ;
      RECT 26.49 2.505 26.64 2.655 ;
      RECT 25.97 3.625 26.12 3.775 ;
      RECT 25.49 1.945 25.64 2.095 ;
      RECT 24.77 1.945 24.92 2.095 ;
      RECT 24.77 3.065 24.92 3.215 ;
      RECT 24.41 3.625 24.56 3.775 ;
      RECT 24.05 1.945 24.2 2.095 ;
      RECT 24.05 3.065 24.2 3.215 ;
      RECT 23.79 2.505 23.94 2.655 ;
      RECT 22.81 2.505 22.96 2.655 ;
      RECT 22.57 1.945 22.72 2.095 ;
      RECT 21.73 3.065 21.88 3.215 ;
      RECT 21.09 3.065 21.24 3.215 ;
      RECT 20.61 1.945 20.76 2.095 ;
      RECT 20.61 3.065 20.76 3.215 ;
      RECT 20.13 2.505 20.28 2.655 ;
      RECT 19.65 3.345 19.8 3.495 ;
      RECT 18.095 1.195 18.245 1.345 ;
      RECT 15.725 6.74 15.875 6.89 ;
      RECT 15.71 2.065 15.86 2.215 ;
      RECT 14.92 2.45 15.07 2.6 ;
      RECT 14.92 6.37 15.07 6.52 ;
      RECT 13.895 2.805 14.045 2.955 ;
      RECT 13.885 5.945 14.035 6.095 ;
      RECT 13.33 3.25 13.48 3.4 ;
      RECT 11.33 1.945 11.48 2.095 ;
      RECT 10.37 3.625 10.52 3.775 ;
      RECT 9.89 1.945 10.04 2.095 ;
      RECT 9.89 3.065 10.04 3.215 ;
      RECT 9.37 3.625 9.52 3.775 ;
      RECT 8.89 3.625 9.04 3.775 ;
      RECT 8.77 1.945 8.92 2.095 ;
      RECT 8.41 3.625 8.56 3.775 ;
      RECT 8.17 1.945 8.32 2.095 ;
      RECT 7.93 2.505 8.08 2.655 ;
      RECT 7.41 3.625 7.56 3.775 ;
      RECT 6.93 1.945 7.08 2.095 ;
      RECT 6.21 1.945 6.36 2.095 ;
      RECT 6.21 3.065 6.36 3.215 ;
      RECT 5.85 3.625 6 3.775 ;
      RECT 5.49 1.945 5.64 2.095 ;
      RECT 5.49 3.065 5.64 3.215 ;
      RECT 5.23 2.505 5.38 2.655 ;
      RECT 4.25 2.505 4.4 2.655 ;
      RECT 4.01 1.945 4.16 2.095 ;
      RECT 3.17 3.065 3.32 3.215 ;
      RECT 2.53 3.065 2.68 3.215 ;
      RECT 2.05 1.945 2.2 2.095 ;
      RECT 2.05 3.065 2.2 3.215 ;
      RECT 1.57 2.505 1.72 2.655 ;
      RECT 1.09 3.345 1.24 3.495 ;
    LAYER met1 ;
      RECT 74.99 0 86.95 1.74 ;
      RECT 56.43 0 68.39 1.74 ;
      RECT 37.87 0 49.83 1.74 ;
      RECT 19.31 0 31.27 1.74 ;
      RECT 0.75 0 12.71 1.74 ;
      RECT 74.99 0 87.035 1.585 ;
      RECT 56.43 0 68.475 1.585 ;
      RECT 37.87 0 49.915 1.585 ;
      RECT 19.31 0 31.355 1.585 ;
      RECT 0.75 0 12.795 1.585 ;
      RECT 0 0 92.805 0.305 ;
      RECT 74.245 4.145 76.71 4.75 ;
      RECT 55.685 4.145 58.15 4.75 ;
      RECT 37.125 4.145 39.59 4.75 ;
      RECT 18.565 4.145 21.03 4.75 ;
      RECT 0.005 4.145 2.47 4.75 ;
      RECT 74.99 4.135 92.805 4.745 ;
      RECT 56.43 4.135 74.245 4.745 ;
      RECT 37.87 4.135 55.685 4.745 ;
      RECT 19.31 4.135 37.125 4.745 ;
      RECT 0.75 4.135 18.565 4.745 ;
      RECT 74.99 3.98 86.95 4.745 ;
      RECT 56.43 3.98 68.39 4.745 ;
      RECT 37.87 3.98 49.83 4.745 ;
      RECT 19.31 3.98 31.27 4.745 ;
      RECT 0.75 3.98 12.71 4.745 ;
      RECT 92.205 2.365 92.495 2.595 ;
      RECT 92.265 0.885 92.435 2.595 ;
      RECT 92.235 1.095 92.575 1.445 ;
      RECT 92.205 0.885 92.495 1.115 ;
      RECT 92.205 7.765 92.495 7.995 ;
      RECT 92.265 6.285 92.435 7.995 ;
      RECT 92.205 6.285 92.495 6.515 ;
      RECT 91.795 2.735 92.125 2.965 ;
      RECT 91.795 2.765 92.295 2.935 ;
      RECT 91.795 2.395 91.985 2.965 ;
      RECT 91.215 2.365 91.505 2.595 ;
      RECT 91.215 2.395 91.985 2.565 ;
      RECT 91.275 0.885 91.445 2.595 ;
      RECT 91.215 0.885 91.505 1.115 ;
      RECT 91.215 7.765 91.505 7.995 ;
      RECT 91.275 6.285 91.445 7.995 ;
      RECT 91.215 6.285 91.505 6.515 ;
      RECT 91.215 6.325 92.065 6.485 ;
      RECT 91.895 5.915 92.065 6.485 ;
      RECT 91.215 6.32 91.605 6.485 ;
      RECT 91.835 5.915 92.125 6.145 ;
      RECT 91.835 5.945 92.295 6.115 ;
      RECT 90.845 2.735 91.135 2.965 ;
      RECT 90.845 2.765 91.305 2.935 ;
      RECT 90.905 1.655 91.07 2.965 ;
      RECT 89.42 1.625 89.71 1.855 ;
      RECT 89.42 1.655 91.07 1.825 ;
      RECT 89.48 0.885 89.65 1.855 ;
      RECT 89.42 0.885 89.71 1.115 ;
      RECT 89.42 7.765 89.71 7.995 ;
      RECT 89.48 7.025 89.65 7.995 ;
      RECT 89.48 7.12 91.07 7.29 ;
      RECT 90.9 5.915 91.07 7.29 ;
      RECT 89.42 7.025 89.71 7.255 ;
      RECT 90.845 5.915 91.135 6.145 ;
      RECT 90.845 5.945 91.305 6.115 ;
      RECT 89.85 1.965 90.2 2.315 ;
      RECT 89.68 2.025 90.2 2.195 ;
      RECT 89.875 6.655 90.2 6.98 ;
      RECT 89.85 6.655 90.2 6.885 ;
      RECT 89.68 6.685 90.2 6.855 ;
      RECT 87.47 3.15 87.81 3.5 ;
      RECT 87.56 2.395 87.73 3.5 ;
      RECT 89.075 2.365 89.395 2.685 ;
      RECT 89.045 2.365 89.395 2.595 ;
      RECT 87.56 2.395 89.395 2.565 ;
      RECT 89.075 6.28 89.395 6.605 ;
      RECT 89.045 6.285 89.395 6.515 ;
      RECT 88.875 6.315 89.395 6.485 ;
      RECT 88.035 2.705 88.375 3.055 ;
      RECT 88.035 2.765 88.51 2.935 ;
      RECT 88.025 5.845 88.365 6.195 ;
      RECT 88.025 5.945 88.51 6.115 ;
      RECT 84.525 3.57 84.845 3.83 ;
      RECT 85.815 2.745 85.955 3.605 ;
      RECT 84.615 3.465 85.955 3.605 ;
      RECT 84.615 3.025 84.755 3.83 ;
      RECT 84.54 3.025 84.83 3.255 ;
      RECT 85.74 2.745 86.03 2.975 ;
      RECT 85.26 3.025 85.55 3.255 ;
      RECT 85.455 1.95 85.595 3.21 ;
      RECT 85.485 1.89 85.805 2.15 ;
      RECT 82.085 2.45 82.405 2.71 ;
      RECT 84.78 2.465 85.07 2.695 ;
      RECT 82.175 2.37 84.995 2.51 ;
      RECT 84.045 1.89 84.365 2.15 ;
      RECT 84.54 1.905 84.83 2.135 ;
      RECT 84.045 1.95 84.83 2.09 ;
      RECT 84.045 3.01 84.365 3.27 ;
      RECT 84.045 2.79 84.275 3.27 ;
      RECT 83.54 2.745 83.83 2.975 ;
      RECT 83.54 2.79 84.275 2.93 ;
      RECT 82.565 3.57 82.885 3.83 ;
      RECT 82.1 3.585 82.39 3.815 ;
      RECT 82.1 3.63 82.885 3.77 ;
      RECT 80.86 2.465 81.15 2.695 ;
      RECT 80.86 2.51 81.795 2.65 ;
      RECT 81.655 1.95 81.795 2.65 ;
      RECT 82.325 1.89 82.645 2.15 ;
      RECT 82.1 1.905 82.645 2.135 ;
      RECT 81.655 1.95 82.645 2.09 ;
      RECT 80.005 3.57 80.325 3.83 ;
      RECT 80.005 3.63 81.075 3.77 ;
      RECT 80.935 3.07 81.075 3.77 ;
      RECT 82.1 3.025 82.39 3.255 ;
      RECT 80.935 3.07 82.39 3.21 ;
      RECT 80.365 1.89 80.685 2.15 ;
      RECT 80.14 1.905 80.685 2.135 ;
      RECT 79.385 2.45 79.705 2.71 ;
      RECT 80.38 2.465 80.67 2.695 ;
      RECT 79.14 2.465 79.705 2.695 ;
      RECT 79.14 2.51 80.67 2.65 ;
      RECT 78.66 3.025 78.95 3.255 ;
      RECT 78.855 1.95 78.995 3.21 ;
      RECT 79.645 1.89 79.965 2.15 ;
      RECT 78.66 1.905 78.95 2.135 ;
      RECT 78.66 1.95 79.965 2.09 ;
      RECT 78.255 3.465 79.355 3.605 ;
      RECT 79.14 3.305 79.43 3.535 ;
      RECT 78.18 3.305 78.47 3.535 ;
      RECT 78.42 2.37 78.71 2.74 ;
      RECT 77.655 2.37 78.71 2.51 ;
      RECT 78.165 1.89 78.485 2.15 ;
      RECT 76.205 1.89 76.525 2.15 ;
      RECT 76.205 1.95 78.485 2.09 ;
      RECT 77.325 3.01 77.645 3.27 ;
      RECT 77.325 3.01 78.155 3.15 ;
      RECT 77.94 2.745 78.155 3.15 ;
      RECT 77.94 2.745 78.23 2.975 ;
      RECT 75.725 2.45 76.045 2.71 ;
      RECT 77.135 2.465 77.425 2.695 ;
      RECT 75.725 2.465 76.27 2.695 ;
      RECT 75.725 2.55 76.675 2.69 ;
      RECT 76.535 2.37 76.675 2.69 ;
      RECT 77.035 2.465 77.425 2.65 ;
      RECT 76.535 2.37 77.175 2.51 ;
      RECT 75.245 3.26 75.565 3.675 ;
      RECT 75.325 1.905 75.48 3.675 ;
      RECT 75.26 1.905 75.55 2.135 ;
      RECT 73.645 2.365 73.935 2.595 ;
      RECT 73.705 0.885 73.875 2.595 ;
      RECT 73.675 1.095 74.015 1.445 ;
      RECT 73.645 0.885 73.935 1.115 ;
      RECT 73.645 7.765 73.935 7.995 ;
      RECT 73.705 6.285 73.875 7.995 ;
      RECT 73.645 6.285 73.935 6.515 ;
      RECT 73.235 2.735 73.565 2.965 ;
      RECT 73.235 2.765 73.735 2.935 ;
      RECT 73.235 2.395 73.425 2.965 ;
      RECT 72.655 2.365 72.945 2.595 ;
      RECT 72.655 2.395 73.425 2.565 ;
      RECT 72.715 0.885 72.885 2.595 ;
      RECT 72.655 0.885 72.945 1.115 ;
      RECT 72.655 7.765 72.945 7.995 ;
      RECT 72.715 6.285 72.885 7.995 ;
      RECT 72.655 6.285 72.945 6.515 ;
      RECT 72.655 6.325 73.505 6.485 ;
      RECT 73.335 5.915 73.505 6.485 ;
      RECT 72.655 6.32 73.045 6.485 ;
      RECT 73.275 5.915 73.565 6.145 ;
      RECT 73.275 5.945 73.735 6.115 ;
      RECT 72.285 2.735 72.575 2.965 ;
      RECT 72.285 2.765 72.745 2.935 ;
      RECT 72.345 1.655 72.51 2.965 ;
      RECT 70.86 1.625 71.15 1.855 ;
      RECT 70.86 1.655 72.51 1.825 ;
      RECT 70.92 0.885 71.09 1.855 ;
      RECT 70.86 0.885 71.15 1.115 ;
      RECT 70.86 7.765 71.15 7.995 ;
      RECT 70.92 7.025 71.09 7.995 ;
      RECT 70.92 7.12 72.51 7.29 ;
      RECT 72.34 5.915 72.51 7.29 ;
      RECT 70.86 7.025 71.15 7.255 ;
      RECT 72.285 5.915 72.575 6.145 ;
      RECT 72.285 5.945 72.745 6.115 ;
      RECT 71.29 1.965 71.64 2.315 ;
      RECT 71.12 2.025 71.64 2.195 ;
      RECT 71.315 6.655 71.64 6.98 ;
      RECT 71.29 6.655 71.64 6.885 ;
      RECT 71.12 6.685 71.64 6.855 ;
      RECT 68.91 3.15 69.25 3.5 ;
      RECT 69 2.395 69.17 3.5 ;
      RECT 70.515 2.365 70.835 2.685 ;
      RECT 70.485 2.365 70.835 2.595 ;
      RECT 69 2.395 70.835 2.565 ;
      RECT 70.515 6.28 70.835 6.605 ;
      RECT 70.485 6.285 70.835 6.515 ;
      RECT 70.315 6.315 70.835 6.485 ;
      RECT 69.475 2.705 69.815 3.055 ;
      RECT 69.475 2.765 69.95 2.935 ;
      RECT 69.465 5.845 69.805 6.195 ;
      RECT 69.465 5.945 69.95 6.115 ;
      RECT 65.965 3.57 66.285 3.83 ;
      RECT 67.255 2.745 67.395 3.605 ;
      RECT 66.055 3.465 67.395 3.605 ;
      RECT 66.055 3.025 66.195 3.83 ;
      RECT 65.98 3.025 66.27 3.255 ;
      RECT 67.18 2.745 67.47 2.975 ;
      RECT 66.7 3.025 66.99 3.255 ;
      RECT 66.895 1.95 67.035 3.21 ;
      RECT 66.925 1.89 67.245 2.15 ;
      RECT 63.525 2.45 63.845 2.71 ;
      RECT 66.22 2.465 66.51 2.695 ;
      RECT 63.615 2.37 66.435 2.51 ;
      RECT 65.485 1.89 65.805 2.15 ;
      RECT 65.98 1.905 66.27 2.135 ;
      RECT 65.485 1.95 66.27 2.09 ;
      RECT 65.485 3.01 65.805 3.27 ;
      RECT 65.485 2.79 65.715 3.27 ;
      RECT 64.98 2.745 65.27 2.975 ;
      RECT 64.98 2.79 65.715 2.93 ;
      RECT 64.005 3.57 64.325 3.83 ;
      RECT 63.54 3.585 63.83 3.815 ;
      RECT 63.54 3.63 64.325 3.77 ;
      RECT 62.3 2.465 62.59 2.695 ;
      RECT 62.3 2.51 63.235 2.65 ;
      RECT 63.095 1.95 63.235 2.65 ;
      RECT 63.765 1.89 64.085 2.15 ;
      RECT 63.54 1.905 64.085 2.135 ;
      RECT 63.095 1.95 64.085 2.09 ;
      RECT 61.445 3.57 61.765 3.83 ;
      RECT 61.445 3.63 62.515 3.77 ;
      RECT 62.375 3.07 62.515 3.77 ;
      RECT 63.54 3.025 63.83 3.255 ;
      RECT 62.375 3.07 63.83 3.21 ;
      RECT 61.805 1.89 62.125 2.15 ;
      RECT 61.58 1.905 62.125 2.135 ;
      RECT 60.825 2.45 61.145 2.71 ;
      RECT 61.82 2.465 62.11 2.695 ;
      RECT 60.58 2.465 61.145 2.695 ;
      RECT 60.58 2.51 62.11 2.65 ;
      RECT 60.1 3.025 60.39 3.255 ;
      RECT 60.295 1.95 60.435 3.21 ;
      RECT 61.085 1.89 61.405 2.15 ;
      RECT 60.1 1.905 60.39 2.135 ;
      RECT 60.1 1.95 61.405 2.09 ;
      RECT 59.695 3.465 60.795 3.605 ;
      RECT 60.58 3.305 60.87 3.535 ;
      RECT 59.62 3.305 59.91 3.535 ;
      RECT 59.86 2.37 60.15 2.74 ;
      RECT 59.095 2.37 60.15 2.51 ;
      RECT 59.605 1.89 59.925 2.15 ;
      RECT 57.645 1.89 57.965 2.15 ;
      RECT 57.645 1.95 59.925 2.09 ;
      RECT 58.765 3.01 59.085 3.27 ;
      RECT 58.765 3.01 59.595 3.15 ;
      RECT 59.38 2.745 59.595 3.15 ;
      RECT 59.38 2.745 59.67 2.975 ;
      RECT 57.165 2.45 57.485 2.71 ;
      RECT 58.575 2.465 58.865 2.695 ;
      RECT 57.165 2.465 57.71 2.695 ;
      RECT 57.165 2.55 58.115 2.69 ;
      RECT 57.975 2.37 58.115 2.69 ;
      RECT 58.475 2.465 58.865 2.65 ;
      RECT 57.975 2.37 58.615 2.51 ;
      RECT 56.685 3.26 57.005 3.675 ;
      RECT 56.765 1.905 56.92 3.675 ;
      RECT 56.7 1.905 56.99 2.135 ;
      RECT 55.085 2.365 55.375 2.595 ;
      RECT 55.145 0.885 55.315 2.595 ;
      RECT 55.115 1.095 55.455 1.445 ;
      RECT 55.085 0.885 55.375 1.115 ;
      RECT 55.085 7.765 55.375 7.995 ;
      RECT 55.145 6.285 55.315 7.995 ;
      RECT 55.085 6.285 55.375 6.515 ;
      RECT 54.675 2.735 55.005 2.965 ;
      RECT 54.675 2.765 55.175 2.935 ;
      RECT 54.675 2.395 54.865 2.965 ;
      RECT 54.095 2.365 54.385 2.595 ;
      RECT 54.095 2.395 54.865 2.565 ;
      RECT 54.155 0.885 54.325 2.595 ;
      RECT 54.095 0.885 54.385 1.115 ;
      RECT 54.095 7.765 54.385 7.995 ;
      RECT 54.155 6.285 54.325 7.995 ;
      RECT 54.095 6.285 54.385 6.515 ;
      RECT 54.095 6.325 54.945 6.485 ;
      RECT 54.775 5.915 54.945 6.485 ;
      RECT 54.095 6.32 54.485 6.485 ;
      RECT 54.715 5.915 55.005 6.145 ;
      RECT 54.715 5.945 55.175 6.115 ;
      RECT 53.725 2.735 54.015 2.965 ;
      RECT 53.725 2.765 54.185 2.935 ;
      RECT 53.785 1.655 53.95 2.965 ;
      RECT 52.3 1.625 52.59 1.855 ;
      RECT 52.3 1.655 53.95 1.825 ;
      RECT 52.36 0.885 52.53 1.855 ;
      RECT 52.3 0.885 52.59 1.115 ;
      RECT 52.3 7.765 52.59 7.995 ;
      RECT 52.36 7.025 52.53 7.995 ;
      RECT 52.36 7.12 53.95 7.29 ;
      RECT 53.78 5.915 53.95 7.29 ;
      RECT 52.3 7.025 52.59 7.255 ;
      RECT 53.725 5.915 54.015 6.145 ;
      RECT 53.725 5.945 54.185 6.115 ;
      RECT 52.73 1.965 53.08 2.315 ;
      RECT 52.56 2.025 53.08 2.195 ;
      RECT 52.755 6.655 53.08 6.98 ;
      RECT 52.73 6.655 53.08 6.885 ;
      RECT 52.56 6.685 53.08 6.855 ;
      RECT 50.35 3.15 50.69 3.5 ;
      RECT 50.44 2.395 50.61 3.5 ;
      RECT 51.955 2.365 52.275 2.685 ;
      RECT 51.925 2.365 52.275 2.595 ;
      RECT 50.44 2.395 52.275 2.565 ;
      RECT 51.955 6.28 52.275 6.605 ;
      RECT 51.925 6.285 52.275 6.515 ;
      RECT 51.755 6.315 52.275 6.485 ;
      RECT 50.915 2.705 51.255 3.055 ;
      RECT 50.915 2.765 51.39 2.935 ;
      RECT 50.905 5.845 51.245 6.195 ;
      RECT 50.905 5.945 51.39 6.115 ;
      RECT 47.405 3.57 47.725 3.83 ;
      RECT 48.695 2.745 48.835 3.605 ;
      RECT 47.495 3.465 48.835 3.605 ;
      RECT 47.495 3.025 47.635 3.83 ;
      RECT 47.42 3.025 47.71 3.255 ;
      RECT 48.62 2.745 48.91 2.975 ;
      RECT 48.14 3.025 48.43 3.255 ;
      RECT 48.335 1.95 48.475 3.21 ;
      RECT 48.365 1.89 48.685 2.15 ;
      RECT 44.965 2.45 45.285 2.71 ;
      RECT 47.66 2.465 47.95 2.695 ;
      RECT 45.055 2.37 47.875 2.51 ;
      RECT 46.925 1.89 47.245 2.15 ;
      RECT 47.42 1.905 47.71 2.135 ;
      RECT 46.925 1.95 47.71 2.09 ;
      RECT 46.925 3.01 47.245 3.27 ;
      RECT 46.925 2.79 47.155 3.27 ;
      RECT 46.42 2.745 46.71 2.975 ;
      RECT 46.42 2.79 47.155 2.93 ;
      RECT 45.445 3.57 45.765 3.83 ;
      RECT 44.98 3.585 45.27 3.815 ;
      RECT 44.98 3.63 45.765 3.77 ;
      RECT 43.74 2.465 44.03 2.695 ;
      RECT 43.74 2.51 44.675 2.65 ;
      RECT 44.535 1.95 44.675 2.65 ;
      RECT 45.205 1.89 45.525 2.15 ;
      RECT 44.98 1.905 45.525 2.135 ;
      RECT 44.535 1.95 45.525 2.09 ;
      RECT 42.885 3.57 43.205 3.83 ;
      RECT 42.885 3.63 43.955 3.77 ;
      RECT 43.815 3.07 43.955 3.77 ;
      RECT 44.98 3.025 45.27 3.255 ;
      RECT 43.815 3.07 45.27 3.21 ;
      RECT 43.245 1.89 43.565 2.15 ;
      RECT 43.02 1.905 43.565 2.135 ;
      RECT 42.265 2.45 42.585 2.71 ;
      RECT 43.26 2.465 43.55 2.695 ;
      RECT 42.02 2.465 42.585 2.695 ;
      RECT 42.02 2.51 43.55 2.65 ;
      RECT 41.54 3.025 41.83 3.255 ;
      RECT 41.735 1.95 41.875 3.21 ;
      RECT 42.525 1.89 42.845 2.15 ;
      RECT 41.54 1.905 41.83 2.135 ;
      RECT 41.54 1.95 42.845 2.09 ;
      RECT 41.135 3.465 42.235 3.605 ;
      RECT 42.02 3.305 42.31 3.535 ;
      RECT 41.06 3.305 41.35 3.535 ;
      RECT 41.3 2.37 41.59 2.74 ;
      RECT 40.535 2.37 41.59 2.51 ;
      RECT 41.045 1.89 41.365 2.15 ;
      RECT 39.085 1.89 39.405 2.15 ;
      RECT 39.085 1.95 41.365 2.09 ;
      RECT 40.205 3.01 40.525 3.27 ;
      RECT 40.205 3.01 41.035 3.15 ;
      RECT 40.82 2.745 41.035 3.15 ;
      RECT 40.82 2.745 41.11 2.975 ;
      RECT 38.605 2.45 38.925 2.71 ;
      RECT 40.015 2.465 40.305 2.695 ;
      RECT 38.605 2.465 39.15 2.695 ;
      RECT 38.605 2.55 39.555 2.69 ;
      RECT 39.415 2.37 39.555 2.69 ;
      RECT 39.915 2.465 40.305 2.65 ;
      RECT 39.415 2.37 40.055 2.51 ;
      RECT 38.125 3.26 38.445 3.675 ;
      RECT 38.205 1.905 38.36 3.675 ;
      RECT 38.14 1.905 38.43 2.135 ;
      RECT 36.525 2.365 36.815 2.595 ;
      RECT 36.585 0.885 36.755 2.595 ;
      RECT 36.585 0.885 36.765 1.45 ;
      RECT 36.565 1.095 36.905 1.445 ;
      RECT 36.525 0.885 36.815 1.115 ;
      RECT 36.525 7.765 36.815 7.995 ;
      RECT 36.585 6.285 36.755 7.995 ;
      RECT 36.525 6.285 36.815 6.515 ;
      RECT 36.115 2.735 36.445 2.965 ;
      RECT 36.115 2.765 36.615 2.935 ;
      RECT 36.115 2.395 36.305 2.965 ;
      RECT 35.535 2.365 35.825 2.595 ;
      RECT 35.535 2.395 36.305 2.565 ;
      RECT 35.595 0.885 35.765 2.595 ;
      RECT 35.535 0.885 35.825 1.115 ;
      RECT 35.535 7.765 35.825 7.995 ;
      RECT 35.595 6.285 35.765 7.995 ;
      RECT 35.535 6.285 35.825 6.515 ;
      RECT 35.535 6.325 36.385 6.485 ;
      RECT 36.215 5.915 36.385 6.485 ;
      RECT 35.535 6.32 35.925 6.485 ;
      RECT 36.155 5.915 36.445 6.145 ;
      RECT 36.155 5.945 36.615 6.115 ;
      RECT 35.165 2.735 35.455 2.965 ;
      RECT 35.165 2.765 35.625 2.935 ;
      RECT 35.225 1.655 35.39 2.965 ;
      RECT 33.74 1.625 34.03 1.855 ;
      RECT 33.74 1.655 35.39 1.825 ;
      RECT 33.8 0.885 33.97 1.855 ;
      RECT 33.74 0.885 34.03 1.115 ;
      RECT 33.74 7.765 34.03 7.995 ;
      RECT 33.8 7.025 33.97 7.995 ;
      RECT 33.8 7.12 35.39 7.29 ;
      RECT 35.22 5.915 35.39 7.29 ;
      RECT 33.74 7.025 34.03 7.255 ;
      RECT 35.165 5.915 35.455 6.145 ;
      RECT 35.165 5.945 35.625 6.115 ;
      RECT 34.17 1.965 34.52 2.315 ;
      RECT 34 2.025 34.52 2.195 ;
      RECT 34.195 6.655 34.52 6.98 ;
      RECT 34.17 6.655 34.52 6.885 ;
      RECT 34 6.685 34.52 6.855 ;
      RECT 31.79 3.15 32.13 3.5 ;
      RECT 31.88 2.395 32.05 3.5 ;
      RECT 33.395 2.365 33.715 2.685 ;
      RECT 33.365 2.365 33.715 2.595 ;
      RECT 31.88 2.395 33.715 2.565 ;
      RECT 33.395 6.28 33.715 6.605 ;
      RECT 33.365 6.285 33.715 6.515 ;
      RECT 33.195 6.315 33.715 6.485 ;
      RECT 32.355 2.705 32.695 3.055 ;
      RECT 32.355 2.765 32.83 2.935 ;
      RECT 32.345 5.845 32.685 6.195 ;
      RECT 32.345 5.945 32.83 6.115 ;
      RECT 28.845 3.57 29.165 3.83 ;
      RECT 30.135 2.745 30.275 3.605 ;
      RECT 28.935 3.465 30.275 3.605 ;
      RECT 28.935 3.025 29.075 3.83 ;
      RECT 28.86 3.025 29.15 3.255 ;
      RECT 30.06 2.745 30.35 2.975 ;
      RECT 29.58 3.025 29.87 3.255 ;
      RECT 29.775 1.95 29.915 3.21 ;
      RECT 29.805 1.89 30.125 2.15 ;
      RECT 26.405 2.45 26.725 2.71 ;
      RECT 29.1 2.465 29.39 2.695 ;
      RECT 26.495 2.37 29.315 2.51 ;
      RECT 28.365 1.89 28.685 2.15 ;
      RECT 28.86 1.905 29.15 2.135 ;
      RECT 28.365 1.95 29.15 2.09 ;
      RECT 28.365 3.01 28.685 3.27 ;
      RECT 28.365 2.79 28.595 3.27 ;
      RECT 27.86 2.745 28.15 2.975 ;
      RECT 27.86 2.79 28.595 2.93 ;
      RECT 26.885 3.57 27.205 3.83 ;
      RECT 26.42 3.585 26.71 3.815 ;
      RECT 26.42 3.63 27.205 3.77 ;
      RECT 25.18 2.465 25.47 2.695 ;
      RECT 25.18 2.51 26.115 2.65 ;
      RECT 25.975 1.95 26.115 2.65 ;
      RECT 26.645 1.89 26.965 2.15 ;
      RECT 26.42 1.905 26.965 2.135 ;
      RECT 25.975 1.95 26.965 2.09 ;
      RECT 24.325 3.57 24.645 3.83 ;
      RECT 24.325 3.63 25.395 3.77 ;
      RECT 25.255 3.07 25.395 3.77 ;
      RECT 26.42 3.025 26.71 3.255 ;
      RECT 25.255 3.07 26.71 3.21 ;
      RECT 24.685 1.89 25.005 2.15 ;
      RECT 24.46 1.905 25.005 2.135 ;
      RECT 23.705 2.45 24.025 2.71 ;
      RECT 24.7 2.465 24.99 2.695 ;
      RECT 23.46 2.465 24.025 2.695 ;
      RECT 23.46 2.51 24.99 2.65 ;
      RECT 22.98 3.025 23.27 3.255 ;
      RECT 23.175 1.95 23.315 3.21 ;
      RECT 23.965 1.89 24.285 2.15 ;
      RECT 22.98 1.905 23.27 2.135 ;
      RECT 22.98 1.95 24.285 2.09 ;
      RECT 22.575 3.465 23.675 3.605 ;
      RECT 23.46 3.305 23.75 3.535 ;
      RECT 22.5 3.305 22.79 3.535 ;
      RECT 22.74 2.37 23.03 2.74 ;
      RECT 21.975 2.37 23.03 2.51 ;
      RECT 22.485 1.89 22.805 2.15 ;
      RECT 20.525 1.89 20.845 2.15 ;
      RECT 20.525 1.95 22.805 2.09 ;
      RECT 21.645 3.01 21.965 3.27 ;
      RECT 21.645 3.01 22.475 3.15 ;
      RECT 22.26 2.745 22.475 3.15 ;
      RECT 22.26 2.745 22.55 2.975 ;
      RECT 20.045 2.45 20.365 2.71 ;
      RECT 21.455 2.465 21.745 2.695 ;
      RECT 20.045 2.465 20.59 2.695 ;
      RECT 20.045 2.55 20.995 2.69 ;
      RECT 20.855 2.37 20.995 2.69 ;
      RECT 21.355 2.465 21.745 2.65 ;
      RECT 20.855 2.37 21.495 2.51 ;
      RECT 19.565 3.26 19.885 3.675 ;
      RECT 19.645 1.905 19.8 3.675 ;
      RECT 19.58 1.905 19.87 2.135 ;
      RECT 17.965 2.365 18.255 2.595 ;
      RECT 18.025 0.885 18.195 2.595 ;
      RECT 17.995 1.095 18.335 1.445 ;
      RECT 17.965 0.885 18.255 1.115 ;
      RECT 17.965 7.765 18.255 7.995 ;
      RECT 18.025 6.285 18.195 7.995 ;
      RECT 17.965 6.285 18.255 6.515 ;
      RECT 17.555 2.735 17.885 2.965 ;
      RECT 17.555 2.765 18.055 2.935 ;
      RECT 17.555 2.395 17.745 2.965 ;
      RECT 16.975 2.365 17.265 2.595 ;
      RECT 16.975 2.395 17.745 2.565 ;
      RECT 17.035 0.885 17.205 2.595 ;
      RECT 16.975 0.885 17.265 1.115 ;
      RECT 16.975 7.765 17.265 7.995 ;
      RECT 17.035 6.285 17.205 7.995 ;
      RECT 16.975 6.285 17.265 6.515 ;
      RECT 16.975 6.325 17.825 6.485 ;
      RECT 17.655 5.915 17.825 6.485 ;
      RECT 16.975 6.32 17.365 6.485 ;
      RECT 17.595 5.915 17.885 6.145 ;
      RECT 17.595 5.945 18.055 6.115 ;
      RECT 16.605 2.735 16.895 2.965 ;
      RECT 16.605 2.765 17.065 2.935 ;
      RECT 16.665 1.655 16.83 2.965 ;
      RECT 15.18 1.625 15.47 1.855 ;
      RECT 15.18 1.655 16.83 1.825 ;
      RECT 15.24 0.885 15.41 1.855 ;
      RECT 15.18 0.885 15.47 1.115 ;
      RECT 15.18 7.765 15.47 7.995 ;
      RECT 15.24 7.025 15.41 7.995 ;
      RECT 15.24 7.12 16.83 7.29 ;
      RECT 16.66 5.915 16.83 7.29 ;
      RECT 15.18 7.025 15.47 7.255 ;
      RECT 16.605 5.915 16.895 6.145 ;
      RECT 16.605 5.945 17.065 6.115 ;
      RECT 15.61 1.965 15.96 2.315 ;
      RECT 15.44 2.025 15.96 2.195 ;
      RECT 15.635 6.655 15.96 6.98 ;
      RECT 15.61 6.655 15.96 6.885 ;
      RECT 15.44 6.685 15.96 6.855 ;
      RECT 13.23 3.15 13.57 3.5 ;
      RECT 13.32 2.395 13.49 3.5 ;
      RECT 14.835 2.365 15.155 2.685 ;
      RECT 14.805 2.365 15.155 2.595 ;
      RECT 13.32 2.395 15.155 2.565 ;
      RECT 14.835 6.28 15.155 6.605 ;
      RECT 14.805 6.285 15.155 6.515 ;
      RECT 14.635 6.315 15.155 6.485 ;
      RECT 13.795 2.705 14.135 3.055 ;
      RECT 13.795 2.765 14.27 2.935 ;
      RECT 13.785 5.845 14.125 6.195 ;
      RECT 13.785 5.945 14.27 6.115 ;
      RECT 10.285 3.57 10.605 3.83 ;
      RECT 11.575 2.745 11.715 3.605 ;
      RECT 10.375 3.465 11.715 3.605 ;
      RECT 10.375 3.025 10.515 3.83 ;
      RECT 10.3 3.025 10.59 3.255 ;
      RECT 11.5 2.745 11.79 2.975 ;
      RECT 11.02 3.025 11.31 3.255 ;
      RECT 11.215 1.95 11.355 3.21 ;
      RECT 11.245 1.89 11.565 2.15 ;
      RECT 7.845 2.45 8.165 2.71 ;
      RECT 10.54 2.465 10.83 2.695 ;
      RECT 7.935 2.37 10.755 2.51 ;
      RECT 9.805 1.89 10.125 2.15 ;
      RECT 10.3 1.905 10.59 2.135 ;
      RECT 9.805 1.95 10.59 2.09 ;
      RECT 9.805 3.01 10.125 3.27 ;
      RECT 9.805 2.79 10.035 3.27 ;
      RECT 9.3 2.745 9.59 2.975 ;
      RECT 9.3 2.79 10.035 2.93 ;
      RECT 8.325 3.57 8.645 3.83 ;
      RECT 7.86 3.585 8.15 3.815 ;
      RECT 7.86 3.63 8.645 3.77 ;
      RECT 6.62 2.465 6.91 2.695 ;
      RECT 6.62 2.51 7.555 2.65 ;
      RECT 7.415 1.95 7.555 2.65 ;
      RECT 8.085 1.89 8.405 2.15 ;
      RECT 7.86 1.905 8.405 2.135 ;
      RECT 7.415 1.95 8.405 2.09 ;
      RECT 5.765 3.57 6.085 3.83 ;
      RECT 5.765 3.63 6.835 3.77 ;
      RECT 6.695 3.07 6.835 3.77 ;
      RECT 7.86 3.025 8.15 3.255 ;
      RECT 6.695 3.07 8.15 3.21 ;
      RECT 6.125 1.89 6.445 2.15 ;
      RECT 5.9 1.905 6.445 2.135 ;
      RECT 5.145 2.45 5.465 2.71 ;
      RECT 6.14 2.465 6.43 2.695 ;
      RECT 4.9 2.465 5.465 2.695 ;
      RECT 4.9 2.51 6.43 2.65 ;
      RECT 4.42 3.025 4.71 3.255 ;
      RECT 4.615 1.95 4.755 3.21 ;
      RECT 5.405 1.89 5.725 2.15 ;
      RECT 4.42 1.905 4.71 2.135 ;
      RECT 4.42 1.95 5.725 2.09 ;
      RECT 4.015 3.465 5.115 3.605 ;
      RECT 4.9 3.305 5.19 3.535 ;
      RECT 3.94 3.305 4.23 3.535 ;
      RECT 4.18 2.37 4.47 2.74 ;
      RECT 3.415 2.37 4.47 2.51 ;
      RECT 3.925 1.89 4.245 2.15 ;
      RECT 1.965 1.89 2.285 2.15 ;
      RECT 1.965 1.95 4.245 2.09 ;
      RECT 3.085 3.01 3.405 3.27 ;
      RECT 3.085 3.01 3.915 3.15 ;
      RECT 3.7 2.745 3.915 3.15 ;
      RECT 3.7 2.745 3.99 2.975 ;
      RECT 1.485 2.45 1.805 2.71 ;
      RECT 2.895 2.465 3.185 2.695 ;
      RECT 1.485 2.465 2.03 2.695 ;
      RECT 1.485 2.55 2.435 2.69 ;
      RECT 2.295 2.37 2.435 2.69 ;
      RECT 2.795 2.465 3.185 2.65 ;
      RECT 2.295 2.37 2.935 2.51 ;
      RECT 1.005 3.26 1.325 3.675 ;
      RECT 1.085 1.905 1.24 3.675 ;
      RECT 1.02 1.905 1.31 2.135 ;
      RECT 0.005 8.575 92.805 8.88 ;
      RECT 86.07 2.735 86.39 3.055 ;
      RECT 83.525 3.57 83.845 3.83 ;
      RECT 82.925 1.89 83.605 2.15 ;
      RECT 83.045 3.57 83.365 3.83 ;
      RECT 81.565 3.57 81.885 3.83 ;
      RECT 81.085 1.89 81.405 2.15 ;
      RECT 80.365 3.01 80.685 3.27 ;
      RECT 79.645 3.01 79.965 3.27 ;
      RECT 76.685 3.01 77.005 3.27 ;
      RECT 76.205 3.01 76.525 3.27 ;
      RECT 67.51 2.735 67.83 3.055 ;
      RECT 64.965 3.57 65.285 3.83 ;
      RECT 64.365 1.89 65.045 2.15 ;
      RECT 64.485 3.57 64.805 3.83 ;
      RECT 63.005 3.57 63.325 3.83 ;
      RECT 62.525 1.89 62.845 2.15 ;
      RECT 61.805 3.01 62.125 3.27 ;
      RECT 61.085 3.01 61.405 3.27 ;
      RECT 58.125 3.01 58.445 3.27 ;
      RECT 57.645 3.01 57.965 3.27 ;
      RECT 48.95 2.735 49.27 3.055 ;
      RECT 46.405 3.57 46.725 3.83 ;
      RECT 45.805 1.89 46.485 2.15 ;
      RECT 45.925 3.57 46.245 3.83 ;
      RECT 44.445 3.57 44.765 3.83 ;
      RECT 43.965 1.89 44.285 2.15 ;
      RECT 43.245 3.01 43.565 3.27 ;
      RECT 42.525 3.01 42.845 3.27 ;
      RECT 39.565 3.01 39.885 3.27 ;
      RECT 39.085 3.01 39.405 3.27 ;
      RECT 30.39 2.735 30.71 3.055 ;
      RECT 27.845 3.57 28.165 3.83 ;
      RECT 27.245 1.89 27.925 2.15 ;
      RECT 27.365 3.57 27.685 3.83 ;
      RECT 25.885 3.57 26.205 3.83 ;
      RECT 25.405 1.89 25.725 2.15 ;
      RECT 24.685 3.01 25.005 3.27 ;
      RECT 23.965 3.01 24.285 3.27 ;
      RECT 21.005 3.01 21.325 3.27 ;
      RECT 20.525 3.01 20.845 3.27 ;
      RECT 11.83 2.735 12.15 3.055 ;
      RECT 9.285 3.57 9.605 3.83 ;
      RECT 8.685 1.89 9.365 2.15 ;
      RECT 8.805 3.57 9.125 3.83 ;
      RECT 7.325 3.57 7.645 3.83 ;
      RECT 6.845 1.89 7.165 2.15 ;
      RECT 6.125 3.01 6.445 3.27 ;
      RECT 5.405 3.01 5.725 3.27 ;
      RECT 2.445 3.01 2.765 3.27 ;
      RECT 1.965 3.01 2.285 3.27 ;
    LAYER mcon ;
      RECT 92.265 0.915 92.435 1.085 ;
      RECT 92.265 2.395 92.435 2.565 ;
      RECT 92.265 6.315 92.435 6.485 ;
      RECT 92.265 7.795 92.435 7.965 ;
      RECT 91.915 0.105 92.085 0.275 ;
      RECT 91.915 4.165 92.085 4.335 ;
      RECT 91.915 4.545 92.085 4.715 ;
      RECT 91.915 8.605 92.085 8.775 ;
      RECT 91.895 2.765 92.065 2.935 ;
      RECT 91.895 5.945 92.065 6.115 ;
      RECT 91.275 0.915 91.445 1.085 ;
      RECT 91.275 2.395 91.445 2.565 ;
      RECT 91.275 6.315 91.445 6.485 ;
      RECT 91.275 7.795 91.445 7.965 ;
      RECT 90.925 0.105 91.095 0.275 ;
      RECT 90.925 4.165 91.095 4.335 ;
      RECT 90.925 4.545 91.095 4.715 ;
      RECT 90.925 8.605 91.095 8.775 ;
      RECT 90.905 2.765 91.075 2.935 ;
      RECT 90.905 5.945 91.075 6.115 ;
      RECT 90.22 0.105 90.39 0.275 ;
      RECT 90.22 4.165 90.39 4.335 ;
      RECT 90.22 4.545 90.39 4.715 ;
      RECT 90.22 8.605 90.39 8.775 ;
      RECT 89.91 2.025 90.08 2.195 ;
      RECT 89.91 6.685 90.08 6.855 ;
      RECT 89.54 0.105 89.71 0.275 ;
      RECT 89.54 8.605 89.71 8.775 ;
      RECT 89.48 0.915 89.65 1.085 ;
      RECT 89.48 1.655 89.65 1.825 ;
      RECT 89.48 7.055 89.65 7.225 ;
      RECT 89.48 7.795 89.65 7.965 ;
      RECT 89.105 2.395 89.275 2.565 ;
      RECT 89.105 6.315 89.275 6.485 ;
      RECT 88.86 0.105 89.03 0.275 ;
      RECT 88.86 8.605 89.03 8.775 ;
      RECT 88.18 0.105 88.35 0.275 ;
      RECT 88.18 8.605 88.35 8.775 ;
      RECT 88.11 2.765 88.28 2.935 ;
      RECT 88.11 5.945 88.28 6.115 ;
      RECT 86.635 1.415 86.805 1.585 ;
      RECT 86.635 4.135 86.805 4.305 ;
      RECT 86.175 1.415 86.345 1.585 ;
      RECT 86.175 4.135 86.345 4.305 ;
      RECT 85.8 2.775 85.97 2.945 ;
      RECT 85.715 1.415 85.885 1.585 ;
      RECT 85.715 4.135 85.885 4.305 ;
      RECT 85.56 1.935 85.73 2.105 ;
      RECT 85.32 3.055 85.49 3.225 ;
      RECT 85.255 1.415 85.425 1.585 ;
      RECT 85.255 4.135 85.425 4.305 ;
      RECT 84.84 2.495 85.01 2.665 ;
      RECT 84.795 1.415 84.965 1.585 ;
      RECT 84.795 4.135 84.965 4.305 ;
      RECT 84.6 1.935 84.77 2.105 ;
      RECT 84.6 3.055 84.77 3.225 ;
      RECT 84.6 3.615 84.77 3.785 ;
      RECT 84.335 1.415 84.505 1.585 ;
      RECT 84.335 4.135 84.505 4.305 ;
      RECT 84.12 3.055 84.29 3.225 ;
      RECT 83.875 1.415 84.045 1.585 ;
      RECT 83.875 4.135 84.045 4.305 ;
      RECT 83.6 2.775 83.77 2.945 ;
      RECT 83.6 3.615 83.77 3.785 ;
      RECT 83.415 1.415 83.585 1.585 ;
      RECT 83.415 4.135 83.585 4.305 ;
      RECT 83.12 1.935 83.29 2.105 ;
      RECT 83.12 3.615 83.29 3.785 ;
      RECT 82.955 1.415 83.125 1.585 ;
      RECT 82.955 4.135 83.125 4.305 ;
      RECT 82.495 1.415 82.665 1.585 ;
      RECT 82.495 4.135 82.665 4.305 ;
      RECT 82.16 1.935 82.33 2.105 ;
      RECT 82.16 2.495 82.33 2.665 ;
      RECT 82.16 3.055 82.33 3.225 ;
      RECT 82.16 3.615 82.33 3.785 ;
      RECT 82.035 1.415 82.205 1.585 ;
      RECT 82.035 4.135 82.205 4.305 ;
      RECT 81.64 3.615 81.81 3.785 ;
      RECT 81.575 1.415 81.745 1.585 ;
      RECT 81.575 4.135 81.745 4.305 ;
      RECT 81.16 1.935 81.33 2.105 ;
      RECT 81.115 1.415 81.285 1.585 ;
      RECT 81.115 4.135 81.285 4.305 ;
      RECT 80.92 2.495 81.09 2.665 ;
      RECT 80.655 1.415 80.825 1.585 ;
      RECT 80.655 4.135 80.825 4.305 ;
      RECT 80.44 2.495 80.61 2.665 ;
      RECT 80.44 3.055 80.61 3.225 ;
      RECT 80.2 1.935 80.37 2.105 ;
      RECT 80.195 1.415 80.365 1.585 ;
      RECT 80.195 4.135 80.365 4.305 ;
      RECT 79.735 1.415 79.905 1.585 ;
      RECT 79.735 4.135 79.905 4.305 ;
      RECT 79.72 3.055 79.89 3.225 ;
      RECT 79.275 1.415 79.445 1.585 ;
      RECT 79.275 4.135 79.445 4.305 ;
      RECT 79.2 2.495 79.37 2.665 ;
      RECT 79.2 3.335 79.37 3.505 ;
      RECT 78.815 1.415 78.985 1.585 ;
      RECT 78.815 4.135 78.985 4.305 ;
      RECT 78.72 1.935 78.89 2.105 ;
      RECT 78.72 3.055 78.89 3.225 ;
      RECT 78.48 2.495 78.65 2.665 ;
      RECT 78.355 1.415 78.525 1.585 ;
      RECT 78.355 4.135 78.525 4.305 ;
      RECT 78.24 3.335 78.41 3.505 ;
      RECT 78 2.775 78.17 2.945 ;
      RECT 77.895 1.415 78.065 1.585 ;
      RECT 77.895 4.135 78.065 4.305 ;
      RECT 77.435 1.415 77.605 1.585 ;
      RECT 77.435 4.135 77.605 4.305 ;
      RECT 77.195 2.495 77.365 2.665 ;
      RECT 76.975 1.415 77.145 1.585 ;
      RECT 76.975 4.135 77.145 4.305 ;
      RECT 76.76 3.055 76.93 3.225 ;
      RECT 76.515 1.415 76.685 1.585 ;
      RECT 76.515 4.135 76.685 4.305 ;
      RECT 76.28 1.935 76.45 2.105 ;
      RECT 76.28 3.055 76.45 3.225 ;
      RECT 76.055 1.415 76.225 1.585 ;
      RECT 76.055 4.135 76.225 4.305 ;
      RECT 76.04 2.495 76.21 2.665 ;
      RECT 75.595 1.415 75.765 1.585 ;
      RECT 75.595 4.135 75.765 4.305 ;
      RECT 75.32 1.935 75.49 2.105 ;
      RECT 75.32 3.475 75.49 3.645 ;
      RECT 75.135 1.415 75.305 1.585 ;
      RECT 75.135 4.135 75.305 4.305 ;
      RECT 73.705 0.915 73.875 1.085 ;
      RECT 73.705 2.395 73.875 2.565 ;
      RECT 73.705 6.315 73.875 6.485 ;
      RECT 73.705 7.795 73.875 7.965 ;
      RECT 73.355 0.105 73.525 0.275 ;
      RECT 73.355 4.165 73.525 4.335 ;
      RECT 73.355 4.545 73.525 4.715 ;
      RECT 73.355 8.605 73.525 8.775 ;
      RECT 73.335 2.765 73.505 2.935 ;
      RECT 73.335 5.945 73.505 6.115 ;
      RECT 72.715 0.915 72.885 1.085 ;
      RECT 72.715 2.395 72.885 2.565 ;
      RECT 72.715 6.315 72.885 6.485 ;
      RECT 72.715 7.795 72.885 7.965 ;
      RECT 72.365 0.105 72.535 0.275 ;
      RECT 72.365 4.165 72.535 4.335 ;
      RECT 72.365 4.545 72.535 4.715 ;
      RECT 72.365 8.605 72.535 8.775 ;
      RECT 72.345 2.765 72.515 2.935 ;
      RECT 72.345 5.945 72.515 6.115 ;
      RECT 71.66 0.105 71.83 0.275 ;
      RECT 71.66 4.165 71.83 4.335 ;
      RECT 71.66 4.545 71.83 4.715 ;
      RECT 71.66 8.605 71.83 8.775 ;
      RECT 71.35 2.025 71.52 2.195 ;
      RECT 71.35 6.685 71.52 6.855 ;
      RECT 70.98 0.105 71.15 0.275 ;
      RECT 70.98 8.605 71.15 8.775 ;
      RECT 70.92 0.915 71.09 1.085 ;
      RECT 70.92 1.655 71.09 1.825 ;
      RECT 70.92 7.055 71.09 7.225 ;
      RECT 70.92 7.795 71.09 7.965 ;
      RECT 70.545 2.395 70.715 2.565 ;
      RECT 70.545 6.315 70.715 6.485 ;
      RECT 70.3 0.105 70.47 0.275 ;
      RECT 70.3 8.605 70.47 8.775 ;
      RECT 69.62 0.105 69.79 0.275 ;
      RECT 69.62 8.605 69.79 8.775 ;
      RECT 69.55 2.765 69.72 2.935 ;
      RECT 69.55 5.945 69.72 6.115 ;
      RECT 68.075 1.415 68.245 1.585 ;
      RECT 68.075 4.135 68.245 4.305 ;
      RECT 67.615 1.415 67.785 1.585 ;
      RECT 67.615 4.135 67.785 4.305 ;
      RECT 67.24 2.775 67.41 2.945 ;
      RECT 67.155 1.415 67.325 1.585 ;
      RECT 67.155 4.135 67.325 4.305 ;
      RECT 67 1.935 67.17 2.105 ;
      RECT 66.76 3.055 66.93 3.225 ;
      RECT 66.695 1.415 66.865 1.585 ;
      RECT 66.695 4.135 66.865 4.305 ;
      RECT 66.28 2.495 66.45 2.665 ;
      RECT 66.235 1.415 66.405 1.585 ;
      RECT 66.235 4.135 66.405 4.305 ;
      RECT 66.04 1.935 66.21 2.105 ;
      RECT 66.04 3.055 66.21 3.225 ;
      RECT 66.04 3.615 66.21 3.785 ;
      RECT 65.775 1.415 65.945 1.585 ;
      RECT 65.775 4.135 65.945 4.305 ;
      RECT 65.56 3.055 65.73 3.225 ;
      RECT 65.315 1.415 65.485 1.585 ;
      RECT 65.315 4.135 65.485 4.305 ;
      RECT 65.04 2.775 65.21 2.945 ;
      RECT 65.04 3.615 65.21 3.785 ;
      RECT 64.855 1.415 65.025 1.585 ;
      RECT 64.855 4.135 65.025 4.305 ;
      RECT 64.56 1.935 64.73 2.105 ;
      RECT 64.56 3.615 64.73 3.785 ;
      RECT 64.395 1.415 64.565 1.585 ;
      RECT 64.395 4.135 64.565 4.305 ;
      RECT 63.935 1.415 64.105 1.585 ;
      RECT 63.935 4.135 64.105 4.305 ;
      RECT 63.6 1.935 63.77 2.105 ;
      RECT 63.6 2.495 63.77 2.665 ;
      RECT 63.6 3.055 63.77 3.225 ;
      RECT 63.6 3.615 63.77 3.785 ;
      RECT 63.475 1.415 63.645 1.585 ;
      RECT 63.475 4.135 63.645 4.305 ;
      RECT 63.08 3.615 63.25 3.785 ;
      RECT 63.015 1.415 63.185 1.585 ;
      RECT 63.015 4.135 63.185 4.305 ;
      RECT 62.6 1.935 62.77 2.105 ;
      RECT 62.555 1.415 62.725 1.585 ;
      RECT 62.555 4.135 62.725 4.305 ;
      RECT 62.36 2.495 62.53 2.665 ;
      RECT 62.095 1.415 62.265 1.585 ;
      RECT 62.095 4.135 62.265 4.305 ;
      RECT 61.88 2.495 62.05 2.665 ;
      RECT 61.88 3.055 62.05 3.225 ;
      RECT 61.64 1.935 61.81 2.105 ;
      RECT 61.635 1.415 61.805 1.585 ;
      RECT 61.635 4.135 61.805 4.305 ;
      RECT 61.175 1.415 61.345 1.585 ;
      RECT 61.175 4.135 61.345 4.305 ;
      RECT 61.16 3.055 61.33 3.225 ;
      RECT 60.715 1.415 60.885 1.585 ;
      RECT 60.715 4.135 60.885 4.305 ;
      RECT 60.64 2.495 60.81 2.665 ;
      RECT 60.64 3.335 60.81 3.505 ;
      RECT 60.255 1.415 60.425 1.585 ;
      RECT 60.255 4.135 60.425 4.305 ;
      RECT 60.16 1.935 60.33 2.105 ;
      RECT 60.16 3.055 60.33 3.225 ;
      RECT 59.92 2.495 60.09 2.665 ;
      RECT 59.795 1.415 59.965 1.585 ;
      RECT 59.795 4.135 59.965 4.305 ;
      RECT 59.68 3.335 59.85 3.505 ;
      RECT 59.44 2.775 59.61 2.945 ;
      RECT 59.335 1.415 59.505 1.585 ;
      RECT 59.335 4.135 59.505 4.305 ;
      RECT 58.875 1.415 59.045 1.585 ;
      RECT 58.875 4.135 59.045 4.305 ;
      RECT 58.635 2.495 58.805 2.665 ;
      RECT 58.415 1.415 58.585 1.585 ;
      RECT 58.415 4.135 58.585 4.305 ;
      RECT 58.2 3.055 58.37 3.225 ;
      RECT 57.955 1.415 58.125 1.585 ;
      RECT 57.955 4.135 58.125 4.305 ;
      RECT 57.72 1.935 57.89 2.105 ;
      RECT 57.72 3.055 57.89 3.225 ;
      RECT 57.495 1.415 57.665 1.585 ;
      RECT 57.495 4.135 57.665 4.305 ;
      RECT 57.48 2.495 57.65 2.665 ;
      RECT 57.035 1.415 57.205 1.585 ;
      RECT 57.035 4.135 57.205 4.305 ;
      RECT 56.76 1.935 56.93 2.105 ;
      RECT 56.76 3.475 56.93 3.645 ;
      RECT 56.575 1.415 56.745 1.585 ;
      RECT 56.575 4.135 56.745 4.305 ;
      RECT 55.145 0.915 55.315 1.085 ;
      RECT 55.145 2.395 55.315 2.565 ;
      RECT 55.145 6.315 55.315 6.485 ;
      RECT 55.145 7.795 55.315 7.965 ;
      RECT 54.795 0.105 54.965 0.275 ;
      RECT 54.795 4.165 54.965 4.335 ;
      RECT 54.795 4.545 54.965 4.715 ;
      RECT 54.795 8.605 54.965 8.775 ;
      RECT 54.775 2.765 54.945 2.935 ;
      RECT 54.775 5.945 54.945 6.115 ;
      RECT 54.155 0.915 54.325 1.085 ;
      RECT 54.155 2.395 54.325 2.565 ;
      RECT 54.155 6.315 54.325 6.485 ;
      RECT 54.155 7.795 54.325 7.965 ;
      RECT 53.805 0.105 53.975 0.275 ;
      RECT 53.805 4.165 53.975 4.335 ;
      RECT 53.805 4.545 53.975 4.715 ;
      RECT 53.805 8.605 53.975 8.775 ;
      RECT 53.785 2.765 53.955 2.935 ;
      RECT 53.785 5.945 53.955 6.115 ;
      RECT 53.1 0.105 53.27 0.275 ;
      RECT 53.1 4.165 53.27 4.335 ;
      RECT 53.1 4.545 53.27 4.715 ;
      RECT 53.1 8.605 53.27 8.775 ;
      RECT 52.79 2.025 52.96 2.195 ;
      RECT 52.79 6.685 52.96 6.855 ;
      RECT 52.42 0.105 52.59 0.275 ;
      RECT 52.42 8.605 52.59 8.775 ;
      RECT 52.36 0.915 52.53 1.085 ;
      RECT 52.36 1.655 52.53 1.825 ;
      RECT 52.36 7.055 52.53 7.225 ;
      RECT 52.36 7.795 52.53 7.965 ;
      RECT 51.985 2.395 52.155 2.565 ;
      RECT 51.985 6.315 52.155 6.485 ;
      RECT 51.74 0.105 51.91 0.275 ;
      RECT 51.74 8.605 51.91 8.775 ;
      RECT 51.06 0.105 51.23 0.275 ;
      RECT 51.06 8.605 51.23 8.775 ;
      RECT 50.99 2.765 51.16 2.935 ;
      RECT 50.99 5.945 51.16 6.115 ;
      RECT 49.515 1.415 49.685 1.585 ;
      RECT 49.515 4.135 49.685 4.305 ;
      RECT 49.055 1.415 49.225 1.585 ;
      RECT 49.055 4.135 49.225 4.305 ;
      RECT 48.68 2.775 48.85 2.945 ;
      RECT 48.595 1.415 48.765 1.585 ;
      RECT 48.595 4.135 48.765 4.305 ;
      RECT 48.44 1.935 48.61 2.105 ;
      RECT 48.2 3.055 48.37 3.225 ;
      RECT 48.135 1.415 48.305 1.585 ;
      RECT 48.135 4.135 48.305 4.305 ;
      RECT 47.72 2.495 47.89 2.665 ;
      RECT 47.675 1.415 47.845 1.585 ;
      RECT 47.675 4.135 47.845 4.305 ;
      RECT 47.48 1.935 47.65 2.105 ;
      RECT 47.48 3.055 47.65 3.225 ;
      RECT 47.48 3.615 47.65 3.785 ;
      RECT 47.215 1.415 47.385 1.585 ;
      RECT 47.215 4.135 47.385 4.305 ;
      RECT 47 3.055 47.17 3.225 ;
      RECT 46.755 1.415 46.925 1.585 ;
      RECT 46.755 4.135 46.925 4.305 ;
      RECT 46.48 2.775 46.65 2.945 ;
      RECT 46.48 3.615 46.65 3.785 ;
      RECT 46.295 1.415 46.465 1.585 ;
      RECT 46.295 4.135 46.465 4.305 ;
      RECT 46 1.935 46.17 2.105 ;
      RECT 46 3.615 46.17 3.785 ;
      RECT 45.835 1.415 46.005 1.585 ;
      RECT 45.835 4.135 46.005 4.305 ;
      RECT 45.375 1.415 45.545 1.585 ;
      RECT 45.375 4.135 45.545 4.305 ;
      RECT 45.04 1.935 45.21 2.105 ;
      RECT 45.04 2.495 45.21 2.665 ;
      RECT 45.04 3.055 45.21 3.225 ;
      RECT 45.04 3.615 45.21 3.785 ;
      RECT 44.915 1.415 45.085 1.585 ;
      RECT 44.915 4.135 45.085 4.305 ;
      RECT 44.52 3.615 44.69 3.785 ;
      RECT 44.455 1.415 44.625 1.585 ;
      RECT 44.455 4.135 44.625 4.305 ;
      RECT 44.04 1.935 44.21 2.105 ;
      RECT 43.995 1.415 44.165 1.585 ;
      RECT 43.995 4.135 44.165 4.305 ;
      RECT 43.8 2.495 43.97 2.665 ;
      RECT 43.535 1.415 43.705 1.585 ;
      RECT 43.535 4.135 43.705 4.305 ;
      RECT 43.32 2.495 43.49 2.665 ;
      RECT 43.32 3.055 43.49 3.225 ;
      RECT 43.08 1.935 43.25 2.105 ;
      RECT 43.075 1.415 43.245 1.585 ;
      RECT 43.075 4.135 43.245 4.305 ;
      RECT 42.615 1.415 42.785 1.585 ;
      RECT 42.615 4.135 42.785 4.305 ;
      RECT 42.6 3.055 42.77 3.225 ;
      RECT 42.155 1.415 42.325 1.585 ;
      RECT 42.155 4.135 42.325 4.305 ;
      RECT 42.08 2.495 42.25 2.665 ;
      RECT 42.08 3.335 42.25 3.505 ;
      RECT 41.695 1.415 41.865 1.585 ;
      RECT 41.695 4.135 41.865 4.305 ;
      RECT 41.6 1.935 41.77 2.105 ;
      RECT 41.6 3.055 41.77 3.225 ;
      RECT 41.36 2.495 41.53 2.665 ;
      RECT 41.235 1.415 41.405 1.585 ;
      RECT 41.235 4.135 41.405 4.305 ;
      RECT 41.12 3.335 41.29 3.505 ;
      RECT 40.88 2.775 41.05 2.945 ;
      RECT 40.775 1.415 40.945 1.585 ;
      RECT 40.775 4.135 40.945 4.305 ;
      RECT 40.315 1.415 40.485 1.585 ;
      RECT 40.315 4.135 40.485 4.305 ;
      RECT 40.075 2.495 40.245 2.665 ;
      RECT 39.855 1.415 40.025 1.585 ;
      RECT 39.855 4.135 40.025 4.305 ;
      RECT 39.64 3.055 39.81 3.225 ;
      RECT 39.395 1.415 39.565 1.585 ;
      RECT 39.395 4.135 39.565 4.305 ;
      RECT 39.16 1.935 39.33 2.105 ;
      RECT 39.16 3.055 39.33 3.225 ;
      RECT 38.935 1.415 39.105 1.585 ;
      RECT 38.935 4.135 39.105 4.305 ;
      RECT 38.92 2.495 39.09 2.665 ;
      RECT 38.475 1.415 38.645 1.585 ;
      RECT 38.475 4.135 38.645 4.305 ;
      RECT 38.2 1.935 38.37 2.105 ;
      RECT 38.2 3.475 38.37 3.645 ;
      RECT 38.015 1.415 38.185 1.585 ;
      RECT 38.015 4.135 38.185 4.305 ;
      RECT 36.585 0.915 36.755 1.085 ;
      RECT 36.585 2.395 36.755 2.565 ;
      RECT 36.585 6.315 36.755 6.485 ;
      RECT 36.585 7.795 36.755 7.965 ;
      RECT 36.235 0.105 36.405 0.275 ;
      RECT 36.235 4.165 36.405 4.335 ;
      RECT 36.235 4.545 36.405 4.715 ;
      RECT 36.235 8.605 36.405 8.775 ;
      RECT 36.215 2.765 36.385 2.935 ;
      RECT 36.215 5.945 36.385 6.115 ;
      RECT 35.595 0.915 35.765 1.085 ;
      RECT 35.595 2.395 35.765 2.565 ;
      RECT 35.595 6.315 35.765 6.485 ;
      RECT 35.595 7.795 35.765 7.965 ;
      RECT 35.245 0.105 35.415 0.275 ;
      RECT 35.245 4.165 35.415 4.335 ;
      RECT 35.245 4.545 35.415 4.715 ;
      RECT 35.245 8.605 35.415 8.775 ;
      RECT 35.225 2.765 35.395 2.935 ;
      RECT 35.225 5.945 35.395 6.115 ;
      RECT 34.54 0.105 34.71 0.275 ;
      RECT 34.54 4.165 34.71 4.335 ;
      RECT 34.54 4.545 34.71 4.715 ;
      RECT 34.54 8.605 34.71 8.775 ;
      RECT 34.23 2.025 34.4 2.195 ;
      RECT 34.23 6.685 34.4 6.855 ;
      RECT 33.86 0.105 34.03 0.275 ;
      RECT 33.86 8.605 34.03 8.775 ;
      RECT 33.8 0.915 33.97 1.085 ;
      RECT 33.8 1.655 33.97 1.825 ;
      RECT 33.8 7.055 33.97 7.225 ;
      RECT 33.8 7.795 33.97 7.965 ;
      RECT 33.425 2.395 33.595 2.565 ;
      RECT 33.425 6.315 33.595 6.485 ;
      RECT 33.18 0.105 33.35 0.275 ;
      RECT 33.18 8.605 33.35 8.775 ;
      RECT 32.5 0.105 32.67 0.275 ;
      RECT 32.5 8.605 32.67 8.775 ;
      RECT 32.43 2.765 32.6 2.935 ;
      RECT 32.43 5.945 32.6 6.115 ;
      RECT 30.955 1.415 31.125 1.585 ;
      RECT 30.955 4.135 31.125 4.305 ;
      RECT 30.495 1.415 30.665 1.585 ;
      RECT 30.495 4.135 30.665 4.305 ;
      RECT 30.12 2.775 30.29 2.945 ;
      RECT 30.035 1.415 30.205 1.585 ;
      RECT 30.035 4.135 30.205 4.305 ;
      RECT 29.88 1.935 30.05 2.105 ;
      RECT 29.64 3.055 29.81 3.225 ;
      RECT 29.575 1.415 29.745 1.585 ;
      RECT 29.575 4.135 29.745 4.305 ;
      RECT 29.16 2.495 29.33 2.665 ;
      RECT 29.115 1.415 29.285 1.585 ;
      RECT 29.115 4.135 29.285 4.305 ;
      RECT 28.92 1.935 29.09 2.105 ;
      RECT 28.92 3.055 29.09 3.225 ;
      RECT 28.92 3.615 29.09 3.785 ;
      RECT 28.655 1.415 28.825 1.585 ;
      RECT 28.655 4.135 28.825 4.305 ;
      RECT 28.44 3.055 28.61 3.225 ;
      RECT 28.195 1.415 28.365 1.585 ;
      RECT 28.195 4.135 28.365 4.305 ;
      RECT 27.92 2.775 28.09 2.945 ;
      RECT 27.92 3.615 28.09 3.785 ;
      RECT 27.735 1.415 27.905 1.585 ;
      RECT 27.735 4.135 27.905 4.305 ;
      RECT 27.44 1.935 27.61 2.105 ;
      RECT 27.44 3.615 27.61 3.785 ;
      RECT 27.275 1.415 27.445 1.585 ;
      RECT 27.275 4.135 27.445 4.305 ;
      RECT 26.815 1.415 26.985 1.585 ;
      RECT 26.815 4.135 26.985 4.305 ;
      RECT 26.48 1.935 26.65 2.105 ;
      RECT 26.48 2.495 26.65 2.665 ;
      RECT 26.48 3.055 26.65 3.225 ;
      RECT 26.48 3.615 26.65 3.785 ;
      RECT 26.355 1.415 26.525 1.585 ;
      RECT 26.355 4.135 26.525 4.305 ;
      RECT 25.96 3.615 26.13 3.785 ;
      RECT 25.895 1.415 26.065 1.585 ;
      RECT 25.895 4.135 26.065 4.305 ;
      RECT 25.48 1.935 25.65 2.105 ;
      RECT 25.435 1.415 25.605 1.585 ;
      RECT 25.435 4.135 25.605 4.305 ;
      RECT 25.24 2.495 25.41 2.665 ;
      RECT 24.975 1.415 25.145 1.585 ;
      RECT 24.975 4.135 25.145 4.305 ;
      RECT 24.76 2.495 24.93 2.665 ;
      RECT 24.76 3.055 24.93 3.225 ;
      RECT 24.52 1.935 24.69 2.105 ;
      RECT 24.515 1.415 24.685 1.585 ;
      RECT 24.515 4.135 24.685 4.305 ;
      RECT 24.055 1.415 24.225 1.585 ;
      RECT 24.055 4.135 24.225 4.305 ;
      RECT 24.04 3.055 24.21 3.225 ;
      RECT 23.595 1.415 23.765 1.585 ;
      RECT 23.595 4.135 23.765 4.305 ;
      RECT 23.52 2.495 23.69 2.665 ;
      RECT 23.52 3.335 23.69 3.505 ;
      RECT 23.135 1.415 23.305 1.585 ;
      RECT 23.135 4.135 23.305 4.305 ;
      RECT 23.04 1.935 23.21 2.105 ;
      RECT 23.04 3.055 23.21 3.225 ;
      RECT 22.8 2.495 22.97 2.665 ;
      RECT 22.675 1.415 22.845 1.585 ;
      RECT 22.675 4.135 22.845 4.305 ;
      RECT 22.56 3.335 22.73 3.505 ;
      RECT 22.32 2.775 22.49 2.945 ;
      RECT 22.215 1.415 22.385 1.585 ;
      RECT 22.215 4.135 22.385 4.305 ;
      RECT 21.755 1.415 21.925 1.585 ;
      RECT 21.755 4.135 21.925 4.305 ;
      RECT 21.515 2.495 21.685 2.665 ;
      RECT 21.295 1.415 21.465 1.585 ;
      RECT 21.295 4.135 21.465 4.305 ;
      RECT 21.08 3.055 21.25 3.225 ;
      RECT 20.835 1.415 21.005 1.585 ;
      RECT 20.835 4.135 21.005 4.305 ;
      RECT 20.6 1.935 20.77 2.105 ;
      RECT 20.6 3.055 20.77 3.225 ;
      RECT 20.375 1.415 20.545 1.585 ;
      RECT 20.375 4.135 20.545 4.305 ;
      RECT 20.36 2.495 20.53 2.665 ;
      RECT 19.915 1.415 20.085 1.585 ;
      RECT 19.915 4.135 20.085 4.305 ;
      RECT 19.64 1.935 19.81 2.105 ;
      RECT 19.64 3.475 19.81 3.645 ;
      RECT 19.455 1.415 19.625 1.585 ;
      RECT 19.455 4.135 19.625 4.305 ;
      RECT 18.025 0.915 18.195 1.085 ;
      RECT 18.025 2.395 18.195 2.565 ;
      RECT 18.025 6.315 18.195 6.485 ;
      RECT 18.025 7.795 18.195 7.965 ;
      RECT 17.675 0.105 17.845 0.275 ;
      RECT 17.675 4.165 17.845 4.335 ;
      RECT 17.675 4.545 17.845 4.715 ;
      RECT 17.675 8.605 17.845 8.775 ;
      RECT 17.655 2.765 17.825 2.935 ;
      RECT 17.655 5.945 17.825 6.115 ;
      RECT 17.035 0.915 17.205 1.085 ;
      RECT 17.035 2.395 17.205 2.565 ;
      RECT 17.035 6.315 17.205 6.485 ;
      RECT 17.035 7.795 17.205 7.965 ;
      RECT 16.685 0.105 16.855 0.275 ;
      RECT 16.685 4.165 16.855 4.335 ;
      RECT 16.685 4.545 16.855 4.715 ;
      RECT 16.685 8.605 16.855 8.775 ;
      RECT 16.665 2.765 16.835 2.935 ;
      RECT 16.665 5.945 16.835 6.115 ;
      RECT 15.98 0.105 16.15 0.275 ;
      RECT 15.98 4.165 16.15 4.335 ;
      RECT 15.98 4.545 16.15 4.715 ;
      RECT 15.98 8.605 16.15 8.775 ;
      RECT 15.67 2.025 15.84 2.195 ;
      RECT 15.67 6.685 15.84 6.855 ;
      RECT 15.3 0.105 15.47 0.275 ;
      RECT 15.3 8.605 15.47 8.775 ;
      RECT 15.24 0.915 15.41 1.085 ;
      RECT 15.24 1.655 15.41 1.825 ;
      RECT 15.24 7.055 15.41 7.225 ;
      RECT 15.24 7.795 15.41 7.965 ;
      RECT 14.865 2.395 15.035 2.565 ;
      RECT 14.865 6.315 15.035 6.485 ;
      RECT 14.62 0.105 14.79 0.275 ;
      RECT 14.62 8.605 14.79 8.775 ;
      RECT 13.94 0.105 14.11 0.275 ;
      RECT 13.94 8.605 14.11 8.775 ;
      RECT 13.87 2.765 14.04 2.935 ;
      RECT 13.87 5.945 14.04 6.115 ;
      RECT 12.395 1.415 12.565 1.585 ;
      RECT 12.395 4.135 12.565 4.305 ;
      RECT 11.935 1.415 12.105 1.585 ;
      RECT 11.935 4.135 12.105 4.305 ;
      RECT 11.56 2.775 11.73 2.945 ;
      RECT 11.475 1.415 11.645 1.585 ;
      RECT 11.475 4.135 11.645 4.305 ;
      RECT 11.32 1.935 11.49 2.105 ;
      RECT 11.08 3.055 11.25 3.225 ;
      RECT 11.015 1.415 11.185 1.585 ;
      RECT 11.015 4.135 11.185 4.305 ;
      RECT 10.6 2.495 10.77 2.665 ;
      RECT 10.555 1.415 10.725 1.585 ;
      RECT 10.555 4.135 10.725 4.305 ;
      RECT 10.36 1.935 10.53 2.105 ;
      RECT 10.36 3.055 10.53 3.225 ;
      RECT 10.36 3.615 10.53 3.785 ;
      RECT 10.095 1.415 10.265 1.585 ;
      RECT 10.095 4.135 10.265 4.305 ;
      RECT 9.88 3.055 10.05 3.225 ;
      RECT 9.635 1.415 9.805 1.585 ;
      RECT 9.635 4.135 9.805 4.305 ;
      RECT 9.36 2.775 9.53 2.945 ;
      RECT 9.36 3.615 9.53 3.785 ;
      RECT 9.175 1.415 9.345 1.585 ;
      RECT 9.175 4.135 9.345 4.305 ;
      RECT 8.88 1.935 9.05 2.105 ;
      RECT 8.88 3.615 9.05 3.785 ;
      RECT 8.715 1.415 8.885 1.585 ;
      RECT 8.715 4.135 8.885 4.305 ;
      RECT 8.255 1.415 8.425 1.585 ;
      RECT 8.255 4.135 8.425 4.305 ;
      RECT 7.92 1.935 8.09 2.105 ;
      RECT 7.92 2.495 8.09 2.665 ;
      RECT 7.92 3.055 8.09 3.225 ;
      RECT 7.92 3.615 8.09 3.785 ;
      RECT 7.795 1.415 7.965 1.585 ;
      RECT 7.795 4.135 7.965 4.305 ;
      RECT 7.4 3.615 7.57 3.785 ;
      RECT 7.335 1.415 7.505 1.585 ;
      RECT 7.335 4.135 7.505 4.305 ;
      RECT 6.92 1.935 7.09 2.105 ;
      RECT 6.875 1.415 7.045 1.585 ;
      RECT 6.875 4.135 7.045 4.305 ;
      RECT 6.68 2.495 6.85 2.665 ;
      RECT 6.415 1.415 6.585 1.585 ;
      RECT 6.415 4.135 6.585 4.305 ;
      RECT 6.2 2.495 6.37 2.665 ;
      RECT 6.2 3.055 6.37 3.225 ;
      RECT 5.96 1.935 6.13 2.105 ;
      RECT 5.955 1.415 6.125 1.585 ;
      RECT 5.955 4.135 6.125 4.305 ;
      RECT 5.495 1.415 5.665 1.585 ;
      RECT 5.495 4.135 5.665 4.305 ;
      RECT 5.48 3.055 5.65 3.225 ;
      RECT 5.035 1.415 5.205 1.585 ;
      RECT 5.035 4.135 5.205 4.305 ;
      RECT 4.96 2.495 5.13 2.665 ;
      RECT 4.96 3.335 5.13 3.505 ;
      RECT 4.575 1.415 4.745 1.585 ;
      RECT 4.575 4.135 4.745 4.305 ;
      RECT 4.48 1.935 4.65 2.105 ;
      RECT 4.48 3.055 4.65 3.225 ;
      RECT 4.24 2.495 4.41 2.665 ;
      RECT 4.115 1.415 4.285 1.585 ;
      RECT 4.115 4.135 4.285 4.305 ;
      RECT 4 3.335 4.17 3.505 ;
      RECT 3.76 2.775 3.93 2.945 ;
      RECT 3.655 1.415 3.825 1.585 ;
      RECT 3.655 4.135 3.825 4.305 ;
      RECT 3.195 1.415 3.365 1.585 ;
      RECT 3.195 4.135 3.365 4.305 ;
      RECT 2.955 2.495 3.125 2.665 ;
      RECT 2.735 1.415 2.905 1.585 ;
      RECT 2.735 4.135 2.905 4.305 ;
      RECT 2.52 3.055 2.69 3.225 ;
      RECT 2.275 1.415 2.445 1.585 ;
      RECT 2.275 4.135 2.445 4.305 ;
      RECT 2.04 1.935 2.21 2.105 ;
      RECT 2.04 3.055 2.21 3.225 ;
      RECT 1.815 1.415 1.985 1.585 ;
      RECT 1.815 4.135 1.985 4.305 ;
      RECT 1.8 2.495 1.97 2.665 ;
      RECT 1.355 1.415 1.525 1.585 ;
      RECT 1.355 4.135 1.525 4.305 ;
      RECT 1.08 1.935 1.25 2.105 ;
      RECT 1.08 3.475 1.25 3.645 ;
      RECT 0.895 1.415 1.065 1.585 ;
      RECT 0.895 4.135 1.065 4.305 ;
    LAYER li ;
      RECT 86.04 0 86.21 2.085 ;
      RECT 85.08 0 85.25 2.085 ;
      RECT 84.12 0 84.29 2.085 ;
      RECT 83.6 0 83.77 2.085 ;
      RECT 82.64 0 82.81 2.085 ;
      RECT 81.64 0 81.81 2.085 ;
      RECT 80.68 0 80.85 2.085 ;
      RECT 79.2 0 79.37 2.085 ;
      RECT 77.28 0 77.45 2.085 ;
      RECT 75.8 0 75.97 2.085 ;
      RECT 67.48 0 67.65 2.085 ;
      RECT 66.52 0 66.69 2.085 ;
      RECT 65.56 0 65.73 2.085 ;
      RECT 65.04 0 65.21 2.085 ;
      RECT 64.08 0 64.25 2.085 ;
      RECT 63.08 0 63.25 2.085 ;
      RECT 62.12 0 62.29 2.085 ;
      RECT 60.64 0 60.81 2.085 ;
      RECT 58.72 0 58.89 2.085 ;
      RECT 57.24 0 57.41 2.085 ;
      RECT 48.92 0 49.09 2.085 ;
      RECT 47.96 0 48.13 2.085 ;
      RECT 47 0 47.17 2.085 ;
      RECT 46.48 0 46.65 2.085 ;
      RECT 45.52 0 45.69 2.085 ;
      RECT 44.52 0 44.69 2.085 ;
      RECT 43.56 0 43.73 2.085 ;
      RECT 42.08 0 42.25 2.085 ;
      RECT 40.16 0 40.33 2.085 ;
      RECT 38.68 0 38.85 2.085 ;
      RECT 30.36 0 30.53 2.085 ;
      RECT 29.4 0 29.57 2.085 ;
      RECT 28.44 0 28.61 2.085 ;
      RECT 27.92 0 28.09 2.085 ;
      RECT 26.96 0 27.13 2.085 ;
      RECT 25.96 0 26.13 2.085 ;
      RECT 25 0 25.17 2.085 ;
      RECT 23.52 0 23.69 2.085 ;
      RECT 21.6 0 21.77 2.085 ;
      RECT 20.12 0 20.29 2.085 ;
      RECT 11.8 0 11.97 2.085 ;
      RECT 10.84 0 11.01 2.085 ;
      RECT 9.88 0 10.05 2.085 ;
      RECT 9.36 0 9.53 2.085 ;
      RECT 8.4 0 8.57 2.085 ;
      RECT 7.4 0 7.57 2.085 ;
      RECT 6.44 0 6.61 2.085 ;
      RECT 4.96 0 5.13 2.085 ;
      RECT 3.04 0 3.21 2.085 ;
      RECT 1.56 0 1.73 2.085 ;
      RECT 83.32 0 83.515 1.595 ;
      RECT 79.645 0 79.84 1.595 ;
      RECT 77.28 0 77.54 1.595 ;
      RECT 64.76 0 64.955 1.595 ;
      RECT 61.085 0 61.28 1.595 ;
      RECT 58.72 0 58.98 1.595 ;
      RECT 46.2 0 46.395 1.595 ;
      RECT 42.525 0 42.72 1.595 ;
      RECT 40.16 0 40.42 1.595 ;
      RECT 27.64 0 27.835 1.595 ;
      RECT 23.965 0 24.16 1.595 ;
      RECT 21.6 0 21.86 1.595 ;
      RECT 9.08 0 9.275 1.595 ;
      RECT 5.405 0 5.6 1.595 ;
      RECT 3.04 0 3.3 1.595 ;
      RECT 74.99 0 87.035 1.585 ;
      RECT 56.43 0 68.475 1.585 ;
      RECT 37.87 0 49.915 1.585 ;
      RECT 19.31 0 31.355 1.585 ;
      RECT 0.75 0 12.795 1.585 ;
      RECT 91.835 0 92.005 0.935 ;
      RECT 90.845 0 91.015 0.935 ;
      RECT 88.1 0 88.27 0.935 ;
      RECT 73.275 0 73.445 0.935 ;
      RECT 72.285 0 72.455 0.935 ;
      RECT 69.54 0 69.71 0.935 ;
      RECT 54.715 0 54.885 0.935 ;
      RECT 53.725 0 53.895 0.935 ;
      RECT 50.98 0 51.15 0.935 ;
      RECT 36.155 0 36.325 0.935 ;
      RECT 35.165 0 35.335 0.935 ;
      RECT 32.42 0 32.59 0.935 ;
      RECT 17.595 0 17.765 0.935 ;
      RECT 16.605 0 16.775 0.935 ;
      RECT 13.86 0 14.03 0.935 ;
      RECT 0 0 92.805 0.305 ;
      RECT 91.835 3.405 92.005 5.475 ;
      RECT 90.845 3.405 91.015 5.475 ;
      RECT 88.1 3.405 88.27 5.475 ;
      RECT 73.275 3.405 73.445 5.475 ;
      RECT 72.285 3.405 72.455 5.475 ;
      RECT 69.54 3.405 69.71 5.475 ;
      RECT 54.715 3.405 54.885 5.475 ;
      RECT 53.725 3.405 53.895 5.475 ;
      RECT 50.98 3.405 51.15 5.475 ;
      RECT 36.155 3.405 36.325 5.475 ;
      RECT 35.165 3.405 35.335 5.475 ;
      RECT 32.42 3.405 32.59 5.475 ;
      RECT 17.595 3.405 17.765 5.475 ;
      RECT 16.605 3.405 16.775 5.475 ;
      RECT 13.86 3.405 14.03 5.475 ;
      RECT 74.245 4.145 76.71 4.75 ;
      RECT 55.685 4.145 58.15 4.75 ;
      RECT 37.125 4.145 39.59 4.75 ;
      RECT 18.565 4.145 21.03 4.75 ;
      RECT 0.005 4.145 2.47 4.75 ;
      RECT 74.99 4.135 92.805 4.745 ;
      RECT 56.43 4.135 74.245 4.745 ;
      RECT 37.87 4.135 55.685 4.745 ;
      RECT 19.31 4.135 37.125 4.745 ;
      RECT 0.75 4.135 18.565 4.745 ;
      RECT 85.08 3.635 85.25 4.745 ;
      RECT 82.64 3.635 82.81 4.745 ;
      RECT 80.68 3.635 80.85 4.745 ;
      RECT 79.72 3.635 79.89 4.745 ;
      RECT 77.76 3.635 77.93 4.745 ;
      RECT 76.76 3.635 76.93 4.745 ;
      RECT 75.8 3.635 75.97 4.75 ;
      RECT 66.52 3.635 66.69 4.745 ;
      RECT 64.08 3.635 64.25 4.745 ;
      RECT 62.12 3.635 62.29 4.745 ;
      RECT 61.16 3.635 61.33 4.745 ;
      RECT 59.2 3.635 59.37 4.745 ;
      RECT 58.2 3.635 58.37 4.745 ;
      RECT 57.24 3.635 57.41 4.75 ;
      RECT 47.96 3.635 48.13 4.745 ;
      RECT 45.52 3.635 45.69 4.745 ;
      RECT 43.56 3.635 43.73 4.745 ;
      RECT 42.6 3.635 42.77 4.745 ;
      RECT 40.64 3.635 40.81 4.745 ;
      RECT 39.64 3.635 39.81 4.745 ;
      RECT 38.68 3.635 38.85 4.75 ;
      RECT 29.4 3.635 29.57 4.745 ;
      RECT 26.96 3.635 27.13 4.745 ;
      RECT 25 3.635 25.17 4.745 ;
      RECT 24.04 3.635 24.21 4.745 ;
      RECT 22.08 3.635 22.25 4.745 ;
      RECT 21.08 3.635 21.25 4.745 ;
      RECT 20.12 3.635 20.29 4.75 ;
      RECT 10.84 3.635 11.01 4.745 ;
      RECT 8.4 3.635 8.57 4.745 ;
      RECT 6.44 3.635 6.61 4.745 ;
      RECT 5.48 3.635 5.65 4.745 ;
      RECT 3.52 3.635 3.69 4.745 ;
      RECT 2.52 3.635 2.69 4.745 ;
      RECT 1.56 3.635 1.73 4.75 ;
      RECT 0.005 8.575 92.805 8.88 ;
      RECT 91.835 7.945 92.005 8.88 ;
      RECT 90.845 7.945 91.015 8.88 ;
      RECT 88.1 7.945 88.27 8.88 ;
      RECT 73.275 7.945 73.445 8.88 ;
      RECT 72.285 7.945 72.455 8.88 ;
      RECT 69.54 7.945 69.71 8.88 ;
      RECT 54.715 7.945 54.885 8.88 ;
      RECT 53.725 7.945 53.895 8.88 ;
      RECT 50.98 7.945 51.15 8.88 ;
      RECT 36.155 7.945 36.325 8.88 ;
      RECT 35.165 7.945 35.335 8.88 ;
      RECT 32.42 7.945 32.59 8.88 ;
      RECT 17.595 7.945 17.765 8.88 ;
      RECT 16.605 7.945 16.775 8.88 ;
      RECT 13.86 7.945 14.03 8.88 ;
      RECT 91.895 1.74 92.065 2.935 ;
      RECT 91.895 1.74 92.36 1.91 ;
      RECT 91.895 6.97 92.36 7.14 ;
      RECT 91.895 5.945 92.065 7.14 ;
      RECT 90.905 1.74 91.075 2.935 ;
      RECT 90.905 1.74 91.37 1.91 ;
      RECT 90.905 6.97 91.37 7.14 ;
      RECT 90.905 5.945 91.075 7.14 ;
      RECT 89.05 2.635 89.22 3.865 ;
      RECT 89.105 0.855 89.275 2.805 ;
      RECT 89.05 0.575 89.22 1.025 ;
      RECT 89.05 7.855 89.22 8.305 ;
      RECT 89.105 6.075 89.275 8.025 ;
      RECT 89.05 5.015 89.22 6.245 ;
      RECT 88.53 0.575 88.7 3.865 ;
      RECT 88.53 2.075 88.935 2.405 ;
      RECT 88.53 1.235 88.935 1.565 ;
      RECT 88.53 5.015 88.7 8.305 ;
      RECT 88.53 7.315 88.935 7.645 ;
      RECT 88.53 6.475 88.935 6.805 ;
      RECT 85.32 3.225 86.29 3.395 ;
      RECT 85.32 3.055 85.49 3.395 ;
      RECT 84.84 2.495 85.01 2.825 ;
      RECT 84.84 2.575 85.57 2.745 ;
      RECT 84.48 3.615 84.77 3.785 ;
      RECT 84.48 2.575 84.65 3.785 ;
      RECT 84.48 3.055 84.77 3.225 ;
      RECT 84.28 2.575 84.65 2.745 ;
      RECT 83.6 2.675 83.77 2.945 ;
      RECT 83.36 2.675 83.77 2.845 ;
      RECT 83.28 2.575 83.61 2.745 ;
      RECT 83.12 3.615 83.77 3.785 ;
      RECT 83.6 3.145 83.77 3.785 ;
      RECT 83.48 3.225 83.77 3.785 ;
      RECT 82.16 2.915 82.33 3.225 ;
      RECT 82.16 2.915 83.05 3.085 ;
      RECT 82.88 2.495 83.05 3.085 ;
      RECT 82.16 2.575 82.65 2.745 ;
      RECT 82.16 2.495 82.33 2.745 ;
      RECT 80.12 3.225 80.61 3.395 ;
      RECT 81.28 2.575 81.45 3.225 ;
      RECT 80.44 3.055 81.45 3.225 ;
      RECT 81.4 2.495 81.57 2.825 ;
      RECT 80.2 1.835 80.37 2.105 ;
      RECT 79.64 1.835 80.37 2.005 ;
      RECT 79.72 2.575 79.89 3.225 ;
      RECT 79.72 2.575 80.21 2.745 ;
      RECT 78.88 2.575 79.37 2.745 ;
      RECT 79.2 2.495 79.37 2.745 ;
      RECT 78.72 1.835 78.89 2.105 ;
      RECT 78.16 1.835 78.89 2.005 ;
      RECT 78.24 3.225 78.41 3.505 ;
      RECT 77.2 3.225 78.49 3.395 ;
      RECT 77.195 2.575 77.77 2.745 ;
      RECT 77.195 2.495 77.365 2.745 ;
      RECT 76.28 1.835 76.45 2.105 ;
      RECT 76.28 1.835 77.01 2.005 ;
      RECT 76.64 3.055 76.93 3.225 ;
      RECT 76.64 2.575 76.81 3.225 ;
      RECT 76.44 2.575 76.81 2.745 ;
      RECT 76.28 3.055 76.45 3.475 ;
      RECT 75.66 3.14 76.45 3.31 ;
      RECT 75.66 2.915 75.83 3.31 ;
      RECT 75.56 2.495 75.73 3.085 ;
      RECT 75.32 2.575 75.73 2.845 ;
      RECT 73.335 1.74 73.505 2.935 ;
      RECT 73.335 1.74 73.8 1.91 ;
      RECT 73.335 6.97 73.8 7.14 ;
      RECT 73.335 5.945 73.505 7.14 ;
      RECT 72.345 1.74 72.515 2.935 ;
      RECT 72.345 1.74 72.81 1.91 ;
      RECT 72.345 6.97 72.81 7.14 ;
      RECT 72.345 5.945 72.515 7.14 ;
      RECT 70.49 2.635 70.66 3.865 ;
      RECT 70.545 0.855 70.715 2.805 ;
      RECT 70.49 0.575 70.66 1.025 ;
      RECT 70.49 7.855 70.66 8.305 ;
      RECT 70.545 6.075 70.715 8.025 ;
      RECT 70.49 5.015 70.66 6.245 ;
      RECT 69.97 0.575 70.14 3.865 ;
      RECT 69.97 2.075 70.375 2.405 ;
      RECT 69.97 1.235 70.375 1.565 ;
      RECT 69.97 5.015 70.14 8.305 ;
      RECT 69.97 7.315 70.375 7.645 ;
      RECT 69.97 6.475 70.375 6.805 ;
      RECT 66.76 3.225 67.73 3.395 ;
      RECT 66.76 3.055 66.93 3.395 ;
      RECT 66.28 2.495 66.45 2.825 ;
      RECT 66.28 2.575 67.01 2.745 ;
      RECT 65.92 3.615 66.21 3.785 ;
      RECT 65.92 2.575 66.09 3.785 ;
      RECT 65.92 3.055 66.21 3.225 ;
      RECT 65.72 2.575 66.09 2.745 ;
      RECT 65.04 2.675 65.21 2.945 ;
      RECT 64.8 2.675 65.21 2.845 ;
      RECT 64.72 2.575 65.05 2.745 ;
      RECT 64.56 3.615 65.21 3.785 ;
      RECT 65.04 3.145 65.21 3.785 ;
      RECT 64.92 3.225 65.21 3.785 ;
      RECT 63.6 2.915 63.77 3.225 ;
      RECT 63.6 2.915 64.49 3.085 ;
      RECT 64.32 2.495 64.49 3.085 ;
      RECT 63.6 2.575 64.09 2.745 ;
      RECT 63.6 2.495 63.77 2.745 ;
      RECT 61.56 3.225 62.05 3.395 ;
      RECT 62.72 2.575 62.89 3.225 ;
      RECT 61.88 3.055 62.89 3.225 ;
      RECT 62.84 2.495 63.01 2.825 ;
      RECT 61.64 1.835 61.81 2.105 ;
      RECT 61.08 1.835 61.81 2.005 ;
      RECT 61.16 2.575 61.33 3.225 ;
      RECT 61.16 2.575 61.65 2.745 ;
      RECT 60.32 2.575 60.81 2.745 ;
      RECT 60.64 2.495 60.81 2.745 ;
      RECT 60.16 1.835 60.33 2.105 ;
      RECT 59.6 1.835 60.33 2.005 ;
      RECT 59.68 3.225 59.85 3.505 ;
      RECT 58.64 3.225 59.93 3.395 ;
      RECT 58.635 2.575 59.21 2.745 ;
      RECT 58.635 2.495 58.805 2.745 ;
      RECT 57.72 1.835 57.89 2.105 ;
      RECT 57.72 1.835 58.45 2.005 ;
      RECT 58.08 3.055 58.37 3.225 ;
      RECT 58.08 2.575 58.25 3.225 ;
      RECT 57.88 2.575 58.25 2.745 ;
      RECT 57.72 3.055 57.89 3.475 ;
      RECT 57.1 3.14 57.89 3.31 ;
      RECT 57.1 2.915 57.27 3.31 ;
      RECT 57 2.495 57.17 3.085 ;
      RECT 56.76 2.575 57.17 2.845 ;
      RECT 54.775 1.74 54.945 2.935 ;
      RECT 54.775 1.74 55.24 1.91 ;
      RECT 54.775 6.97 55.24 7.14 ;
      RECT 54.775 5.945 54.945 7.14 ;
      RECT 53.785 1.74 53.955 2.935 ;
      RECT 53.785 1.74 54.25 1.91 ;
      RECT 53.785 6.97 54.25 7.14 ;
      RECT 53.785 5.945 53.955 7.14 ;
      RECT 51.93 2.635 52.1 3.865 ;
      RECT 51.985 0.855 52.155 2.805 ;
      RECT 51.93 0.575 52.1 1.025 ;
      RECT 51.93 7.855 52.1 8.305 ;
      RECT 51.985 6.075 52.155 8.025 ;
      RECT 51.93 5.015 52.1 6.245 ;
      RECT 51.41 0.575 51.58 3.865 ;
      RECT 51.41 2.075 51.815 2.405 ;
      RECT 51.41 1.235 51.815 1.565 ;
      RECT 51.41 5.015 51.58 8.305 ;
      RECT 51.41 7.315 51.815 7.645 ;
      RECT 51.41 6.475 51.815 6.805 ;
      RECT 48.2 3.225 49.17 3.395 ;
      RECT 48.2 3.055 48.37 3.395 ;
      RECT 47.72 2.495 47.89 2.825 ;
      RECT 47.72 2.575 48.45 2.745 ;
      RECT 47.36 3.615 47.65 3.785 ;
      RECT 47.36 2.575 47.53 3.785 ;
      RECT 47.36 3.055 47.65 3.225 ;
      RECT 47.16 2.575 47.53 2.745 ;
      RECT 46.48 2.675 46.65 2.945 ;
      RECT 46.24 2.675 46.65 2.845 ;
      RECT 46.16 2.575 46.49 2.745 ;
      RECT 46 3.615 46.65 3.785 ;
      RECT 46.48 3.145 46.65 3.785 ;
      RECT 46.36 3.225 46.65 3.785 ;
      RECT 45.04 2.915 45.21 3.225 ;
      RECT 45.04 2.915 45.93 3.085 ;
      RECT 45.76 2.495 45.93 3.085 ;
      RECT 45.04 2.575 45.53 2.745 ;
      RECT 45.04 2.495 45.21 2.745 ;
      RECT 43 3.225 43.49 3.395 ;
      RECT 44.16 2.575 44.33 3.225 ;
      RECT 43.32 3.055 44.33 3.225 ;
      RECT 44.28 2.495 44.45 2.825 ;
      RECT 43.08 1.835 43.25 2.105 ;
      RECT 42.52 1.835 43.25 2.005 ;
      RECT 42.6 2.575 42.77 3.225 ;
      RECT 42.6 2.575 43.09 2.745 ;
      RECT 41.76 2.575 42.25 2.745 ;
      RECT 42.08 2.495 42.25 2.745 ;
      RECT 41.6 1.835 41.77 2.105 ;
      RECT 41.04 1.835 41.77 2.005 ;
      RECT 41.12 3.225 41.29 3.505 ;
      RECT 40.08 3.225 41.37 3.395 ;
      RECT 40.075 2.575 40.65 2.745 ;
      RECT 40.075 2.495 40.245 2.745 ;
      RECT 39.16 1.835 39.33 2.105 ;
      RECT 39.16 1.835 39.89 2.005 ;
      RECT 39.52 3.055 39.81 3.225 ;
      RECT 39.52 2.575 39.69 3.225 ;
      RECT 39.32 2.575 39.69 2.745 ;
      RECT 39.16 3.055 39.33 3.475 ;
      RECT 38.54 3.14 39.33 3.31 ;
      RECT 38.54 2.915 38.71 3.31 ;
      RECT 38.44 2.495 38.61 3.085 ;
      RECT 38.2 2.575 38.61 2.845 ;
      RECT 36.215 1.74 36.385 2.935 ;
      RECT 36.215 1.74 36.68 1.91 ;
      RECT 36.215 6.97 36.68 7.14 ;
      RECT 36.215 5.945 36.385 7.14 ;
      RECT 35.225 1.74 35.395 2.935 ;
      RECT 35.225 1.74 35.69 1.91 ;
      RECT 35.225 6.97 35.69 7.14 ;
      RECT 35.225 5.945 35.395 7.14 ;
      RECT 33.37 2.635 33.54 3.865 ;
      RECT 33.425 0.855 33.595 2.805 ;
      RECT 33.37 0.575 33.54 1.025 ;
      RECT 33.37 7.855 33.54 8.305 ;
      RECT 33.425 6.075 33.595 8.025 ;
      RECT 33.37 5.015 33.54 6.245 ;
      RECT 32.85 0.575 33.02 3.865 ;
      RECT 32.85 2.075 33.255 2.405 ;
      RECT 32.85 1.235 33.255 1.565 ;
      RECT 32.85 5.015 33.02 8.305 ;
      RECT 32.85 7.315 33.255 7.645 ;
      RECT 32.85 6.475 33.255 6.805 ;
      RECT 29.64 3.225 30.61 3.395 ;
      RECT 29.64 3.055 29.81 3.395 ;
      RECT 29.16 2.495 29.33 2.825 ;
      RECT 29.16 2.575 29.89 2.745 ;
      RECT 28.8 3.615 29.09 3.785 ;
      RECT 28.8 2.575 28.97 3.785 ;
      RECT 28.8 3.055 29.09 3.225 ;
      RECT 28.6 2.575 28.97 2.745 ;
      RECT 27.92 2.675 28.09 2.945 ;
      RECT 27.68 2.675 28.09 2.845 ;
      RECT 27.6 2.575 27.93 2.745 ;
      RECT 27.44 3.615 28.09 3.785 ;
      RECT 27.92 3.145 28.09 3.785 ;
      RECT 27.8 3.225 28.09 3.785 ;
      RECT 26.48 2.915 26.65 3.225 ;
      RECT 26.48 2.915 27.37 3.085 ;
      RECT 27.2 2.495 27.37 3.085 ;
      RECT 26.48 2.575 26.97 2.745 ;
      RECT 26.48 2.495 26.65 2.745 ;
      RECT 24.44 3.225 24.93 3.395 ;
      RECT 25.6 2.575 25.77 3.225 ;
      RECT 24.76 3.055 25.77 3.225 ;
      RECT 25.72 2.495 25.89 2.825 ;
      RECT 24.52 1.835 24.69 2.105 ;
      RECT 23.96 1.835 24.69 2.005 ;
      RECT 24.04 2.575 24.21 3.225 ;
      RECT 24.04 2.575 24.53 2.745 ;
      RECT 23.2 2.575 23.69 2.745 ;
      RECT 23.52 2.495 23.69 2.745 ;
      RECT 23.04 1.835 23.21 2.105 ;
      RECT 22.48 1.835 23.21 2.005 ;
      RECT 22.56 3.225 22.73 3.505 ;
      RECT 21.52 3.225 22.81 3.395 ;
      RECT 21.515 2.575 22.09 2.745 ;
      RECT 21.515 2.495 21.685 2.745 ;
      RECT 20.6 1.835 20.77 2.105 ;
      RECT 20.6 1.835 21.33 2.005 ;
      RECT 20.96 3.055 21.25 3.225 ;
      RECT 20.96 2.575 21.13 3.225 ;
      RECT 20.76 2.575 21.13 2.745 ;
      RECT 20.6 3.055 20.77 3.475 ;
      RECT 19.98 3.14 20.77 3.31 ;
      RECT 19.98 2.915 20.15 3.31 ;
      RECT 19.88 2.495 20.05 3.085 ;
      RECT 19.64 2.575 20.05 2.845 ;
      RECT 17.655 1.74 17.825 2.935 ;
      RECT 17.655 1.74 18.12 1.91 ;
      RECT 17.655 6.97 18.12 7.14 ;
      RECT 17.655 5.945 17.825 7.14 ;
      RECT 16.665 1.74 16.835 2.935 ;
      RECT 16.665 1.74 17.13 1.91 ;
      RECT 16.665 6.97 17.13 7.14 ;
      RECT 16.665 5.945 16.835 7.14 ;
      RECT 14.81 2.635 14.98 3.865 ;
      RECT 14.865 0.855 15.035 2.805 ;
      RECT 14.81 0.575 14.98 1.025 ;
      RECT 14.81 7.855 14.98 8.305 ;
      RECT 14.865 6.075 15.035 8.025 ;
      RECT 14.81 5.015 14.98 6.245 ;
      RECT 14.29 0.575 14.46 3.865 ;
      RECT 14.29 2.075 14.695 2.405 ;
      RECT 14.29 1.235 14.695 1.565 ;
      RECT 14.29 5.015 14.46 8.305 ;
      RECT 14.29 7.315 14.695 7.645 ;
      RECT 14.29 6.475 14.695 6.805 ;
      RECT 11.08 3.225 12.05 3.395 ;
      RECT 11.08 3.055 11.25 3.395 ;
      RECT 10.6 2.495 10.77 2.825 ;
      RECT 10.6 2.575 11.33 2.745 ;
      RECT 10.24 3.615 10.53 3.785 ;
      RECT 10.24 2.575 10.41 3.785 ;
      RECT 10.24 3.055 10.53 3.225 ;
      RECT 10.04 2.575 10.41 2.745 ;
      RECT 9.36 2.675 9.53 2.945 ;
      RECT 9.12 2.675 9.53 2.845 ;
      RECT 9.04 2.575 9.37 2.745 ;
      RECT 8.88 3.615 9.53 3.785 ;
      RECT 9.36 3.145 9.53 3.785 ;
      RECT 9.24 3.225 9.53 3.785 ;
      RECT 7.92 2.915 8.09 3.225 ;
      RECT 7.92 2.915 8.81 3.085 ;
      RECT 8.64 2.495 8.81 3.085 ;
      RECT 7.92 2.575 8.41 2.745 ;
      RECT 7.92 2.495 8.09 2.745 ;
      RECT 5.88 3.225 6.37 3.395 ;
      RECT 7.04 2.575 7.21 3.225 ;
      RECT 6.2 3.055 7.21 3.225 ;
      RECT 7.16 2.495 7.33 2.825 ;
      RECT 5.96 1.835 6.13 2.105 ;
      RECT 5.4 1.835 6.13 2.005 ;
      RECT 5.48 2.575 5.65 3.225 ;
      RECT 5.48 2.575 5.97 2.745 ;
      RECT 4.64 2.575 5.13 2.745 ;
      RECT 4.96 2.495 5.13 2.745 ;
      RECT 4.48 1.835 4.65 2.105 ;
      RECT 3.92 1.835 4.65 2.005 ;
      RECT 4 3.225 4.17 3.505 ;
      RECT 2.96 3.225 4.25 3.395 ;
      RECT 2.955 2.575 3.53 2.745 ;
      RECT 2.955 2.495 3.125 2.745 ;
      RECT 2.04 1.835 2.21 2.105 ;
      RECT 2.04 1.835 2.77 2.005 ;
      RECT 2.4 3.055 2.69 3.225 ;
      RECT 2.4 2.575 2.57 3.225 ;
      RECT 2.2 2.575 2.57 2.745 ;
      RECT 2.04 3.055 2.21 3.475 ;
      RECT 1.42 3.14 2.21 3.31 ;
      RECT 1.42 2.915 1.59 3.31 ;
      RECT 1.32 2.495 1.49 3.085 ;
      RECT 1.08 2.575 1.49 2.845 ;
      RECT 92.265 0.575 92.435 1.085 ;
      RECT 92.265 2.395 92.435 3.865 ;
      RECT 92.265 5.015 92.435 6.485 ;
      RECT 92.265 7.795 92.435 8.305 ;
      RECT 91.275 0.575 91.445 1.085 ;
      RECT 91.275 2.395 91.445 3.865 ;
      RECT 91.275 5.015 91.445 6.485 ;
      RECT 91.275 7.795 91.445 8.305 ;
      RECT 89.91 0.575 90.08 3.865 ;
      RECT 89.91 5.015 90.08 8.305 ;
      RECT 89.48 0.575 89.65 1.085 ;
      RECT 89.48 1.655 89.65 3.865 ;
      RECT 89.48 5.015 89.65 7.225 ;
      RECT 89.48 7.795 89.65 8.305 ;
      RECT 88.11 1.66 88.28 2.935 ;
      RECT 88.11 5.945 88.28 7.22 ;
      RECT 85.8 2.495 85.97 2.945 ;
      RECT 85.56 1.755 85.73 2.105 ;
      RECT 84.6 1.755 84.77 2.105 ;
      RECT 84.12 3.055 84.29 3.475 ;
      RECT 83.12 1.755 83.29 2.105 ;
      RECT 82.16 1.755 82.33 2.105 ;
      RECT 82.16 3.485 82.33 3.815 ;
      RECT 81.64 3.145 81.81 3.785 ;
      RECT 81.16 1.755 81.33 2.105 ;
      RECT 80.92 2.495 81.09 2.825 ;
      RECT 80.44 2.495 80.61 2.825 ;
      RECT 79.2 3.145 79.37 3.505 ;
      RECT 78.72 3.055 78.89 3.475 ;
      RECT 78.48 2.495 78.65 2.825 ;
      RECT 78 2.495 78.17 2.945 ;
      RECT 76.04 2.495 76.21 2.825 ;
      RECT 75.32 1.755 75.49 2.105 ;
      RECT 75.32 3.285 75.49 3.645 ;
      RECT 73.705 0.575 73.875 1.085 ;
      RECT 73.705 2.395 73.875 3.865 ;
      RECT 73.705 5.015 73.875 6.485 ;
      RECT 73.705 7.795 73.875 8.305 ;
      RECT 72.715 0.575 72.885 1.085 ;
      RECT 72.715 2.395 72.885 3.865 ;
      RECT 72.715 5.015 72.885 6.485 ;
      RECT 72.715 7.795 72.885 8.305 ;
      RECT 71.35 0.575 71.52 3.865 ;
      RECT 71.35 5.015 71.52 8.305 ;
      RECT 70.92 0.575 71.09 1.085 ;
      RECT 70.92 1.655 71.09 3.865 ;
      RECT 70.92 5.015 71.09 7.225 ;
      RECT 70.92 7.795 71.09 8.305 ;
      RECT 69.55 1.66 69.72 2.935 ;
      RECT 69.55 5.945 69.72 7.22 ;
      RECT 67.24 2.495 67.41 2.945 ;
      RECT 67 1.755 67.17 2.105 ;
      RECT 66.04 1.755 66.21 2.105 ;
      RECT 65.56 3.055 65.73 3.475 ;
      RECT 64.56 1.755 64.73 2.105 ;
      RECT 63.6 1.755 63.77 2.105 ;
      RECT 63.6 3.485 63.77 3.815 ;
      RECT 63.08 3.145 63.25 3.785 ;
      RECT 62.6 1.755 62.77 2.105 ;
      RECT 62.36 2.495 62.53 2.825 ;
      RECT 61.88 2.495 62.05 2.825 ;
      RECT 60.64 3.145 60.81 3.505 ;
      RECT 60.16 3.055 60.33 3.475 ;
      RECT 59.92 2.495 60.09 2.825 ;
      RECT 59.44 2.495 59.61 2.945 ;
      RECT 57.48 2.495 57.65 2.825 ;
      RECT 56.76 1.755 56.93 2.105 ;
      RECT 56.76 3.285 56.93 3.645 ;
      RECT 55.145 0.575 55.315 1.085 ;
      RECT 55.145 2.395 55.315 3.865 ;
      RECT 55.145 5.015 55.315 6.485 ;
      RECT 55.145 7.795 55.315 8.305 ;
      RECT 54.155 0.575 54.325 1.085 ;
      RECT 54.155 2.395 54.325 3.865 ;
      RECT 54.155 5.015 54.325 6.485 ;
      RECT 54.155 7.795 54.325 8.305 ;
      RECT 52.79 0.575 52.96 3.865 ;
      RECT 52.79 5.015 52.96 8.305 ;
      RECT 52.36 0.575 52.53 1.085 ;
      RECT 52.36 1.655 52.53 3.865 ;
      RECT 52.36 5.015 52.53 7.225 ;
      RECT 52.36 7.795 52.53 8.305 ;
      RECT 50.99 1.66 51.16 2.935 ;
      RECT 50.99 5.945 51.16 7.22 ;
      RECT 48.68 2.495 48.85 2.945 ;
      RECT 48.44 1.755 48.61 2.105 ;
      RECT 47.48 1.755 47.65 2.105 ;
      RECT 47 3.055 47.17 3.475 ;
      RECT 46 1.755 46.17 2.105 ;
      RECT 45.04 1.755 45.21 2.105 ;
      RECT 45.04 3.485 45.21 3.815 ;
      RECT 44.52 3.145 44.69 3.785 ;
      RECT 44.04 1.755 44.21 2.105 ;
      RECT 43.8 2.495 43.97 2.825 ;
      RECT 43.32 2.495 43.49 2.825 ;
      RECT 42.08 3.145 42.25 3.505 ;
      RECT 41.6 3.055 41.77 3.475 ;
      RECT 41.36 2.495 41.53 2.825 ;
      RECT 40.88 2.495 41.05 2.945 ;
      RECT 38.92 2.495 39.09 2.825 ;
      RECT 38.2 1.755 38.37 2.105 ;
      RECT 38.2 3.285 38.37 3.645 ;
      RECT 36.585 0.575 36.755 1.085 ;
      RECT 36.585 2.395 36.755 3.865 ;
      RECT 36.585 5.015 36.755 6.485 ;
      RECT 36.585 7.795 36.755 8.305 ;
      RECT 35.595 0.575 35.765 1.085 ;
      RECT 35.595 2.395 35.765 3.865 ;
      RECT 35.595 5.015 35.765 6.485 ;
      RECT 35.595 7.795 35.765 8.305 ;
      RECT 34.23 0.575 34.4 3.865 ;
      RECT 34.23 5.015 34.4 8.305 ;
      RECT 33.8 0.575 33.97 1.085 ;
      RECT 33.8 1.655 33.97 3.865 ;
      RECT 33.8 5.015 33.97 7.225 ;
      RECT 33.8 7.795 33.97 8.305 ;
      RECT 32.43 1.66 32.6 2.935 ;
      RECT 32.43 5.945 32.6 7.22 ;
      RECT 30.12 2.495 30.29 2.945 ;
      RECT 29.88 1.755 30.05 2.105 ;
      RECT 28.92 1.755 29.09 2.105 ;
      RECT 28.44 3.055 28.61 3.475 ;
      RECT 27.44 1.755 27.61 2.105 ;
      RECT 26.48 1.755 26.65 2.105 ;
      RECT 26.48 3.485 26.65 3.815 ;
      RECT 25.96 3.145 26.13 3.785 ;
      RECT 25.48 1.755 25.65 2.105 ;
      RECT 25.24 2.495 25.41 2.825 ;
      RECT 24.76 2.495 24.93 2.825 ;
      RECT 23.52 3.145 23.69 3.505 ;
      RECT 23.04 3.055 23.21 3.475 ;
      RECT 22.8 2.495 22.97 2.825 ;
      RECT 22.32 2.495 22.49 2.945 ;
      RECT 20.36 2.495 20.53 2.825 ;
      RECT 19.64 1.755 19.81 2.105 ;
      RECT 19.64 3.285 19.81 3.645 ;
      RECT 18.025 0.575 18.195 1.085 ;
      RECT 18.025 2.395 18.195 3.865 ;
      RECT 18.025 5.015 18.195 6.485 ;
      RECT 18.025 7.795 18.195 8.305 ;
      RECT 17.035 0.575 17.205 1.085 ;
      RECT 17.035 2.395 17.205 3.865 ;
      RECT 17.035 5.015 17.205 6.485 ;
      RECT 17.035 7.795 17.205 8.305 ;
      RECT 15.67 0.575 15.84 3.865 ;
      RECT 15.67 5.015 15.84 8.305 ;
      RECT 15.24 0.575 15.41 1.085 ;
      RECT 15.24 1.655 15.41 3.865 ;
      RECT 15.24 5.015 15.41 7.225 ;
      RECT 15.24 7.795 15.41 8.305 ;
      RECT 13.87 1.66 14.04 2.935 ;
      RECT 13.87 5.945 14.04 7.22 ;
      RECT 11.56 2.495 11.73 2.945 ;
      RECT 11.32 1.755 11.49 2.105 ;
      RECT 10.36 1.755 10.53 2.105 ;
      RECT 9.88 3.055 10.05 3.475 ;
      RECT 8.88 1.755 9.05 2.105 ;
      RECT 7.92 1.755 8.09 2.105 ;
      RECT 7.92 3.485 8.09 3.815 ;
      RECT 7.4 3.145 7.57 3.785 ;
      RECT 6.92 1.755 7.09 2.105 ;
      RECT 6.68 2.495 6.85 2.825 ;
      RECT 6.2 2.495 6.37 2.825 ;
      RECT 4.96 3.145 5.13 3.505 ;
      RECT 4.48 3.055 4.65 3.475 ;
      RECT 4.24 2.495 4.41 2.825 ;
      RECT 3.76 2.495 3.93 2.945 ;
      RECT 1.8 2.495 1.97 2.825 ;
      RECT 1.08 1.755 1.25 2.105 ;
      RECT 1.08 3.285 1.25 3.645 ;
  END
END sky130_osu_ring_oscillator_mpr2et_8

MACRO sky130_osu_ring_oscillator_mpr2xa_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2xa_8 0 0 ;
  SIZE 76.3 BY 8.88 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met4 ;
      RECT 63.94 2.975 64.27 3.305 ;
      RECT 63.955 2.5 64.27 3.305 ;
      RECT 66.1 2.485 66.43 2.84 ;
      RECT 63.955 2.5 66.43 2.8 ;
      RECT 48.68 2.975 49.01 3.305 ;
      RECT 48.695 2.5 49.01 3.305 ;
      RECT 50.84 2.485 51.17 2.84 ;
      RECT 48.695 2.5 51.17 2.8 ;
      RECT 33.42 2.975 33.75 3.305 ;
      RECT 33.435 2.5 33.75 3.305 ;
      RECT 35.58 2.485 35.91 2.84 ;
      RECT 33.435 2.5 35.91 2.8 ;
      RECT 18.16 2.975 18.49 3.305 ;
      RECT 18.175 2.5 18.49 3.305 ;
      RECT 20.32 2.485 20.65 2.84 ;
      RECT 18.175 2.5 20.65 2.8 ;
      RECT 2.9 2.975 3.23 3.305 ;
      RECT 2.915 2.5 3.23 3.305 ;
      RECT 5.06 2.485 5.39 2.84 ;
      RECT 2.915 2.5 5.39 2.8 ;
    LAYER via3 ;
      RECT 66.165 2.575 66.365 2.775 ;
      RECT 64.005 3.04 64.205 3.24 ;
      RECT 50.905 2.575 51.105 2.775 ;
      RECT 48.745 3.04 48.945 3.24 ;
      RECT 35.645 2.575 35.845 2.775 ;
      RECT 33.485 3.04 33.685 3.24 ;
      RECT 20.385 2.575 20.585 2.775 ;
      RECT 18.225 3.04 18.425 3.24 ;
      RECT 5.125 2.575 5.325 2.775 ;
      RECT 2.965 3.04 3.165 3.24 ;
    LAYER met3 ;
      RECT 66.58 3.51 66.91 3.865 ;
      RECT 64.675 3.55 66.91 3.85 ;
      RECT 64.675 2.415 64.975 3.85 ;
      RECT 64.66 2.415 64.99 2.745 ;
      RECT 65.65 2.52 66.43 2.865 ;
      RECT 66.125 2.485 66.43 2.865 ;
      RECT 66.105 2.515 66.43 2.865 ;
      RECT 65.225 1.88 65.955 2.21 ;
      RECT 65.37 1.06 65.675 2.21 ;
      RECT 65.34 1.06 65.715 1.43 ;
      RECT 63.945 2.415 64.265 3.33 ;
      RECT 63.945 2.415 64.275 2.95 ;
      RECT 51.32 3.51 51.65 3.865 ;
      RECT 49.415 3.55 51.65 3.85 ;
      RECT 49.415 2.415 49.715 3.85 ;
      RECT 49.4 2.415 49.73 2.745 ;
      RECT 50.39 2.52 51.17 2.865 ;
      RECT 50.865 2.485 51.17 2.865 ;
      RECT 50.845 2.515 51.17 2.865 ;
      RECT 49.965 1.88 50.695 2.21 ;
      RECT 50.11 1.06 50.415 2.21 ;
      RECT 50.08 1.06 50.455 1.43 ;
      RECT 48.685 2.415 49.005 3.33 ;
      RECT 48.685 2.415 49.015 2.95 ;
      RECT 36.06 3.51 36.39 3.865 ;
      RECT 34.155 3.55 36.39 3.85 ;
      RECT 34.155 2.415 34.455 3.85 ;
      RECT 34.14 2.415 34.47 2.745 ;
      RECT 35.13 2.52 35.91 2.865 ;
      RECT 35.605 2.485 35.91 2.865 ;
      RECT 35.585 2.515 35.91 2.865 ;
      RECT 34.705 1.88 35.435 2.21 ;
      RECT 34.85 1.06 35.155 2.21 ;
      RECT 34.82 1.06 35.195 1.43 ;
      RECT 33.425 2.415 33.745 3.33 ;
      RECT 33.425 2.415 33.755 2.95 ;
      RECT 20.8 3.51 21.13 3.865 ;
      RECT 18.895 3.55 21.13 3.85 ;
      RECT 18.895 2.415 19.195 3.85 ;
      RECT 18.88 2.415 19.21 2.745 ;
      RECT 19.87 2.52 20.65 2.865 ;
      RECT 20.345 2.485 20.65 2.865 ;
      RECT 20.325 2.515 20.65 2.865 ;
      RECT 19.445 1.88 20.175 2.21 ;
      RECT 19.59 1.06 19.895 2.21 ;
      RECT 19.56 1.06 19.935 1.43 ;
      RECT 18.165 2.415 18.485 3.33 ;
      RECT 18.165 2.415 18.495 2.95 ;
      RECT 5.54 3.51 5.87 3.865 ;
      RECT 3.635 3.55 5.87 3.85 ;
      RECT 3.635 2.415 3.935 3.85 ;
      RECT 3.62 2.415 3.95 2.745 ;
      RECT 4.61 2.52 5.39 2.865 ;
      RECT 5.085 2.485 5.39 2.865 ;
      RECT 5.065 2.515 5.39 2.865 ;
      RECT 4.185 1.88 4.915 2.21 ;
      RECT 4.33 1.06 4.635 2.21 ;
      RECT 4.3 1.06 4.675 1.43 ;
      RECT 2.905 2.415 3.225 3.33 ;
      RECT 2.905 2.415 3.235 2.95 ;
      RECT 69.5 1.855 70.23 2.185 ;
      RECT 67.81 1.87 68.54 2.2 ;
      RECT 66.775 1.855 67.505 2.205 ;
      RECT 62.755 2.975 63.485 3.305 ;
      RECT 62.62 1.855 63.35 2.185 ;
      RECT 54.24 1.855 54.97 2.185 ;
      RECT 52.55 1.87 53.28 2.2 ;
      RECT 51.515 1.855 52.245 2.205 ;
      RECT 47.495 2.975 48.225 3.305 ;
      RECT 47.36 1.855 48.09 2.185 ;
      RECT 38.98 1.855 39.71 2.185 ;
      RECT 37.29 1.87 38.02 2.2 ;
      RECT 36.255 1.855 36.985 2.205 ;
      RECT 32.235 2.975 32.965 3.305 ;
      RECT 32.1 1.855 32.83 2.185 ;
      RECT 23.72 1.855 24.45 2.185 ;
      RECT 22.03 1.87 22.76 2.2 ;
      RECT 20.995 1.855 21.725 2.205 ;
      RECT 16.975 2.975 17.705 3.305 ;
      RECT 16.84 1.855 17.57 2.185 ;
      RECT 8.46 1.855 9.19 2.185 ;
      RECT 6.77 1.87 7.5 2.2 ;
      RECT 5.735 1.855 6.465 2.205 ;
      RECT 1.715 2.975 2.445 3.305 ;
      RECT 1.58 1.855 2.31 2.185 ;
    LAYER via2 ;
      RECT 69.735 1.92 69.935 2.12 ;
      RECT 67.875 1.935 68.075 2.135 ;
      RECT 66.855 1.94 67.055 2.14 ;
      RECT 66.645 3.575 66.845 3.775 ;
      RECT 66.165 2.575 66.365 2.775 ;
      RECT 65.43 1.145 65.63 1.345 ;
      RECT 65.415 1.945 65.615 2.145 ;
      RECT 64.725 2.48 64.925 2.68 ;
      RECT 64.01 2.48 64.21 2.68 ;
      RECT 63.045 3.04 63.245 3.24 ;
      RECT 62.805 1.92 63.005 2.12 ;
      RECT 54.475 1.92 54.675 2.12 ;
      RECT 52.615 1.935 52.815 2.135 ;
      RECT 51.595 1.94 51.795 2.14 ;
      RECT 51.385 3.575 51.585 3.775 ;
      RECT 50.905 2.575 51.105 2.775 ;
      RECT 50.17 1.145 50.37 1.345 ;
      RECT 50.155 1.945 50.355 2.145 ;
      RECT 49.465 2.48 49.665 2.68 ;
      RECT 48.75 2.48 48.95 2.68 ;
      RECT 47.785 3.04 47.985 3.24 ;
      RECT 47.545 1.92 47.745 2.12 ;
      RECT 39.215 1.92 39.415 2.12 ;
      RECT 37.355 1.935 37.555 2.135 ;
      RECT 36.335 1.94 36.535 2.14 ;
      RECT 36.125 3.575 36.325 3.775 ;
      RECT 35.645 2.575 35.845 2.775 ;
      RECT 34.91 1.145 35.11 1.345 ;
      RECT 34.895 1.945 35.095 2.145 ;
      RECT 34.205 2.48 34.405 2.68 ;
      RECT 33.49 2.48 33.69 2.68 ;
      RECT 32.525 3.04 32.725 3.24 ;
      RECT 32.285 1.92 32.485 2.12 ;
      RECT 23.955 1.92 24.155 2.12 ;
      RECT 22.095 1.935 22.295 2.135 ;
      RECT 21.075 1.94 21.275 2.14 ;
      RECT 20.865 3.575 21.065 3.775 ;
      RECT 20.385 2.575 20.585 2.775 ;
      RECT 19.65 1.145 19.85 1.345 ;
      RECT 19.635 1.945 19.835 2.145 ;
      RECT 18.945 2.48 19.145 2.68 ;
      RECT 18.23 2.48 18.43 2.68 ;
      RECT 17.265 3.04 17.465 3.24 ;
      RECT 17.025 1.92 17.225 2.12 ;
      RECT 8.695 1.92 8.895 2.12 ;
      RECT 6.835 1.935 7.035 2.135 ;
      RECT 5.815 1.94 6.015 2.14 ;
      RECT 5.605 3.575 5.805 3.775 ;
      RECT 5.125 2.575 5.325 2.775 ;
      RECT 4.39 1.145 4.59 1.345 ;
      RECT 4.375 1.945 4.575 2.145 ;
      RECT 3.685 2.48 3.885 2.68 ;
      RECT 2.97 2.48 3.17 2.68 ;
      RECT 2.005 3.04 2.205 3.24 ;
      RECT 1.765 1.92 1.965 2.12 ;
    LAYER met2 ;
      RECT 11.53 6.28 11.85 6.605 ;
      RECT 11.56 5.695 11.73 6.605 ;
      RECT 11.56 5.695 11.735 6.045 ;
      RECT 11.56 5.695 12.535 5.87 ;
      RECT 12.36 1.965 12.535 5.87 ;
      RECT 12.305 1.965 12.655 2.315 ;
      RECT 1.725 1.835 2.005 2.205 ;
      RECT 9.895 2.025 12.655 2.195 ;
      RECT 1.725 1.86 2.115 2.18 ;
      RECT 9.895 0.745 10.065 2.195 ;
      RECT 1.875 0.745 2.045 2.18 ;
      RECT 9.89 0.23 10.06 1.53 ;
      RECT 75.74 1.09 76.08 1.44 ;
      RECT 75.74 1.16 76.085 1.36 ;
      RECT 75.76 0.23 75.93 1.44 ;
      RECT 1.875 0.745 10.065 0.915 ;
      RECT 9.89 0.23 75.93 0.4 ;
      RECT 72.57 6.28 72.89 6.605 ;
      RECT 72.6 5.695 72.77 6.605 ;
      RECT 72.6 5.695 72.775 6.045 ;
      RECT 72.6 5.695 73.575 5.87 ;
      RECT 73.4 1.965 73.575 5.87 ;
      RECT 73.345 1.965 73.695 2.315 ;
      RECT 62.765 1.835 63.045 2.205 ;
      RECT 70.935 2.025 73.695 2.195 ;
      RECT 62.765 1.86 63.155 2.18 ;
      RECT 70.935 0.745 71.105 2.195 ;
      RECT 62.915 0.745 63.085 2.18 ;
      RECT 61.64 1.26 63.085 1.46 ;
      RECT 60.475 1.095 60.815 1.445 ;
      RECT 60.475 1.165 61.78 1.365 ;
      RECT 62.915 0.745 71.105 0.915 ;
      RECT 73.37 6.655 73.695 6.98 ;
      RECT 72.255 6.745 73.695 6.915 ;
      RECT 72.255 2.395 72.415 6.915 ;
      RECT 72.57 2.365 72.89 2.685 ;
      RECT 72.255 2.395 72.89 2.565 ;
      RECT 71.525 5.86 71.865 6.21 ;
      RECT 71.605 2.705 71.775 6.21 ;
      RECT 71.525 2.705 71.865 3.055 ;
      RECT 70.965 2.7 71.305 3.05 ;
      RECT 70.455 2.77 71.305 2.97 ;
      RECT 70.455 1.18 70.655 2.97 ;
      RECT 71.055 2.695 71.225 3.05 ;
      RECT 65.34 1.06 65.715 1.43 ;
      RECT 65.34 1.18 70.655 1.38 ;
      RECT 69.705 3.54 69.965 3.86 ;
      RECT 69.765 1.835 69.905 3.86 ;
      RECT 69.59 2.395 69.905 2.765 ;
      RECT 69.66 1.95 69.905 2.765 ;
      RECT 69.695 1.835 69.975 2.205 ;
      RECT 69.015 2.42 69.275 2.74 ;
      RECT 68.355 2.51 69.275 2.65 ;
      RECT 68.355 1.57 68.495 2.65 ;
      RECT 64.815 1.86 65.075 2.18 ;
      RECT 64.995 1.57 65.135 2.09 ;
      RECT 64.995 1.57 68.495 1.71 ;
      RECT 67.845 3.26 68.105 3.58 ;
      RECT 67.905 1.85 68.045 3.58 ;
      RECT 67.835 1.85 68.115 2.22 ;
      RECT 65.235 4.01 67.67 4.15 ;
      RECT 67.53 2.7 67.67 4.15 ;
      RECT 65.235 3.63 65.375 4.15 ;
      RECT 64.935 3.63 65.375 3.86 ;
      RECT 62.595 3.63 65.375 3.77 ;
      RECT 64.935 3.54 65.195 3.86 ;
      RECT 62.595 3.35 62.735 3.77 ;
      RECT 62.085 3.26 62.345 3.58 ;
      RECT 62.085 3.35 62.735 3.49 ;
      RECT 62.145 1.86 62.285 3.58 ;
      RECT 67.47 2.7 67.73 3.02 ;
      RECT 62.085 1.86 62.345 2.18 ;
      RECT 67.095 3.54 67.355 3.86 ;
      RECT 67.155 1.95 67.295 3.86 ;
      RECT 66.815 1.95 67.295 2.225 ;
      RECT 66.615 1.855 67.095 2.2 ;
      RECT 66.605 3.49 66.885 3.86 ;
      RECT 66.675 2.395 66.815 3.86 ;
      RECT 66.615 2.395 66.875 3.02 ;
      RECT 66.605 2.395 66.885 2.765 ;
      RECT 65.535 3.54 65.795 3.86 ;
      RECT 65.535 3.35 65.735 3.86 ;
      RECT 65.34 3.35 65.735 3.49 ;
      RECT 65.34 1.86 65.48 3.49 ;
      RECT 65.34 1.86 65.655 2.23 ;
      RECT 65.28 1.86 65.655 2.18 ;
      RECT 63.005 2.955 63.285 3.325 ;
      RECT 64.455 2.98 64.715 3.3 ;
      RECT 62.835 3.07 64.715 3.21 ;
      RECT 62.835 2.955 63.285 3.21 ;
      RECT 62.775 2.395 63.035 3.02 ;
      RECT 62.765 2.395 63.045 2.765 ;
      RECT 63.845 2.395 64.255 2.765 ;
      RECT 63.255 2.42 63.515 2.74 ;
      RECT 63.255 2.51 64.255 2.65 ;
      RECT 57.31 6.28 57.63 6.605 ;
      RECT 57.34 5.695 57.51 6.605 ;
      RECT 57.34 5.695 57.515 6.045 ;
      RECT 57.34 5.695 58.315 5.87 ;
      RECT 58.14 1.965 58.315 5.87 ;
      RECT 58.085 1.965 58.435 2.315 ;
      RECT 47.505 1.835 47.785 2.205 ;
      RECT 55.675 2.025 58.435 2.195 ;
      RECT 47.505 1.86 47.895 2.18 ;
      RECT 55.675 0.745 55.845 2.195 ;
      RECT 47.655 0.745 47.825 2.18 ;
      RECT 46.39 1.255 47.825 1.455 ;
      RECT 45.215 1.095 45.555 1.445 ;
      RECT 45.215 1.165 46.53 1.365 ;
      RECT 47.655 0.745 55.845 0.915 ;
      RECT 58.11 6.655 58.435 6.98 ;
      RECT 56.995 6.745 58.435 6.915 ;
      RECT 56.995 2.395 57.155 6.915 ;
      RECT 57.31 2.365 57.63 2.685 ;
      RECT 56.995 2.395 57.63 2.565 ;
      RECT 56.265 5.86 56.605 6.21 ;
      RECT 56.345 2.705 56.515 6.21 ;
      RECT 56.265 2.705 56.605 3.055 ;
      RECT 55.705 2.7 56.045 3.05 ;
      RECT 55.195 2.77 56.045 2.97 ;
      RECT 55.195 1.18 55.395 2.97 ;
      RECT 55.795 2.695 55.965 3.05 ;
      RECT 50.08 1.06 50.455 1.43 ;
      RECT 50.08 1.18 55.395 1.38 ;
      RECT 54.445 3.54 54.705 3.86 ;
      RECT 54.505 1.835 54.645 3.86 ;
      RECT 54.33 2.395 54.645 2.765 ;
      RECT 54.4 1.95 54.645 2.765 ;
      RECT 54.435 1.835 54.715 2.205 ;
      RECT 53.755 2.42 54.015 2.74 ;
      RECT 53.095 2.51 54.015 2.65 ;
      RECT 53.095 1.57 53.235 2.65 ;
      RECT 49.555 1.86 49.815 2.18 ;
      RECT 49.735 1.57 49.875 2.09 ;
      RECT 49.735 1.57 53.235 1.71 ;
      RECT 52.585 3.26 52.845 3.58 ;
      RECT 52.645 1.85 52.785 3.58 ;
      RECT 52.575 1.85 52.855 2.22 ;
      RECT 49.975 4.01 52.41 4.15 ;
      RECT 52.27 2.7 52.41 4.15 ;
      RECT 49.975 3.63 50.115 4.15 ;
      RECT 49.675 3.63 50.115 3.86 ;
      RECT 47.335 3.63 50.115 3.77 ;
      RECT 49.675 3.54 49.935 3.86 ;
      RECT 47.335 3.35 47.475 3.77 ;
      RECT 46.825 3.26 47.085 3.58 ;
      RECT 46.825 3.35 47.475 3.49 ;
      RECT 46.885 1.86 47.025 3.58 ;
      RECT 52.21 2.7 52.47 3.02 ;
      RECT 46.825 1.86 47.085 2.18 ;
      RECT 51.835 3.54 52.095 3.86 ;
      RECT 51.895 1.95 52.035 3.86 ;
      RECT 51.555 1.95 52.035 2.225 ;
      RECT 51.355 1.855 51.835 2.2 ;
      RECT 51.345 3.49 51.625 3.86 ;
      RECT 51.415 2.395 51.555 3.86 ;
      RECT 51.355 2.395 51.615 3.02 ;
      RECT 51.345 2.395 51.625 2.765 ;
      RECT 50.275 3.54 50.535 3.86 ;
      RECT 50.275 3.35 50.475 3.86 ;
      RECT 50.08 3.35 50.475 3.49 ;
      RECT 50.08 1.86 50.22 3.49 ;
      RECT 50.08 1.86 50.395 2.23 ;
      RECT 50.02 1.86 50.395 2.18 ;
      RECT 47.745 2.955 48.025 3.325 ;
      RECT 49.195 2.98 49.455 3.3 ;
      RECT 47.575 3.07 49.455 3.21 ;
      RECT 47.575 2.955 48.025 3.21 ;
      RECT 47.515 2.395 47.775 3.02 ;
      RECT 47.505 2.395 47.785 2.765 ;
      RECT 48.585 2.395 48.995 2.765 ;
      RECT 47.995 2.42 48.255 2.74 ;
      RECT 47.995 2.51 48.995 2.65 ;
      RECT 42.05 6.28 42.37 6.605 ;
      RECT 42.08 5.695 42.25 6.605 ;
      RECT 42.08 5.695 42.255 6.045 ;
      RECT 42.08 5.695 43.055 5.87 ;
      RECT 42.88 1.965 43.055 5.87 ;
      RECT 42.825 1.965 43.175 2.315 ;
      RECT 32.245 1.835 32.525 2.205 ;
      RECT 40.415 2.025 43.175 2.195 ;
      RECT 32.245 1.86 32.635 2.18 ;
      RECT 40.415 0.745 40.585 2.195 ;
      RECT 32.395 0.745 32.565 2.18 ;
      RECT 31.13 1.255 32.565 1.455 ;
      RECT 29.955 1.095 30.295 1.445 ;
      RECT 29.955 1.165 31.27 1.365 ;
      RECT 32.395 0.745 40.585 0.915 ;
      RECT 42.85 6.655 43.175 6.98 ;
      RECT 41.735 6.745 43.175 6.915 ;
      RECT 41.735 2.395 41.895 6.915 ;
      RECT 42.05 2.365 42.37 2.685 ;
      RECT 41.735 2.395 42.37 2.565 ;
      RECT 41.005 5.86 41.345 6.21 ;
      RECT 41.085 2.705 41.255 6.21 ;
      RECT 41.005 2.705 41.345 3.055 ;
      RECT 40.445 2.7 40.785 3.05 ;
      RECT 39.935 2.77 40.785 2.97 ;
      RECT 39.935 1.18 40.135 2.97 ;
      RECT 40.535 2.695 40.705 3.05 ;
      RECT 34.82 1.06 35.195 1.43 ;
      RECT 34.82 1.18 40.135 1.38 ;
      RECT 39.185 3.54 39.445 3.86 ;
      RECT 39.245 1.835 39.385 3.86 ;
      RECT 39.07 2.395 39.385 2.765 ;
      RECT 39.14 1.95 39.385 2.765 ;
      RECT 39.175 1.835 39.455 2.205 ;
      RECT 38.495 2.42 38.755 2.74 ;
      RECT 37.835 2.51 38.755 2.65 ;
      RECT 37.835 1.57 37.975 2.65 ;
      RECT 34.295 1.86 34.555 2.18 ;
      RECT 34.475 1.57 34.615 2.09 ;
      RECT 34.475 1.57 37.975 1.71 ;
      RECT 37.325 3.26 37.585 3.58 ;
      RECT 37.385 1.85 37.525 3.58 ;
      RECT 37.315 1.85 37.595 2.22 ;
      RECT 34.715 4.01 37.15 4.15 ;
      RECT 37.01 2.7 37.15 4.15 ;
      RECT 34.715 3.63 34.855 4.15 ;
      RECT 34.415 3.63 34.855 3.86 ;
      RECT 32.075 3.63 34.855 3.77 ;
      RECT 34.415 3.54 34.675 3.86 ;
      RECT 32.075 3.35 32.215 3.77 ;
      RECT 31.565 3.26 31.825 3.58 ;
      RECT 31.565 3.35 32.215 3.49 ;
      RECT 31.625 1.86 31.765 3.58 ;
      RECT 36.95 2.7 37.21 3.02 ;
      RECT 31.565 1.86 31.825 2.18 ;
      RECT 36.575 3.54 36.835 3.86 ;
      RECT 36.635 1.95 36.775 3.86 ;
      RECT 36.295 1.95 36.775 2.225 ;
      RECT 36.095 1.855 36.575 2.2 ;
      RECT 36.085 3.49 36.365 3.86 ;
      RECT 36.155 2.395 36.295 3.86 ;
      RECT 36.095 2.395 36.355 3.02 ;
      RECT 36.085 2.395 36.365 2.765 ;
      RECT 35.015 3.54 35.275 3.86 ;
      RECT 35.015 3.35 35.215 3.86 ;
      RECT 34.82 3.35 35.215 3.49 ;
      RECT 34.82 1.86 34.96 3.49 ;
      RECT 34.82 1.86 35.135 2.23 ;
      RECT 34.76 1.86 35.135 2.18 ;
      RECT 32.485 2.955 32.765 3.325 ;
      RECT 33.935 2.98 34.195 3.3 ;
      RECT 32.315 3.07 34.195 3.21 ;
      RECT 32.315 2.955 32.765 3.21 ;
      RECT 32.255 2.395 32.515 3.02 ;
      RECT 32.245 2.395 32.525 2.765 ;
      RECT 33.325 2.395 33.735 2.765 ;
      RECT 32.735 2.42 32.995 2.74 ;
      RECT 32.735 2.51 33.735 2.65 ;
      RECT 26.79 6.28 27.11 6.605 ;
      RECT 26.82 5.695 26.99 6.605 ;
      RECT 26.82 5.695 26.995 6.045 ;
      RECT 26.82 5.695 27.795 5.87 ;
      RECT 27.62 1.965 27.795 5.87 ;
      RECT 27.565 1.965 27.915 2.315 ;
      RECT 16.985 1.835 17.265 2.205 ;
      RECT 25.155 2.025 27.915 2.195 ;
      RECT 16.985 1.86 17.375 2.18 ;
      RECT 25.155 0.745 25.325 2.195 ;
      RECT 17.135 0.745 17.305 2.18 ;
      RECT 15.87 1.26 17.305 1.46 ;
      RECT 14.7 1.1 15.04 1.45 ;
      RECT 14.7 1.17 16.01 1.37 ;
      RECT 17.135 0.745 25.325 0.915 ;
      RECT 27.59 6.655 27.915 6.98 ;
      RECT 26.475 6.745 27.915 6.915 ;
      RECT 26.475 2.395 26.635 6.915 ;
      RECT 26.79 2.365 27.11 2.685 ;
      RECT 26.475 2.395 27.11 2.565 ;
      RECT 25.745 5.86 26.085 6.21 ;
      RECT 25.825 2.705 25.995 6.21 ;
      RECT 25.745 2.705 26.085 3.055 ;
      RECT 25.185 2.7 25.525 3.05 ;
      RECT 24.675 2.77 25.525 2.97 ;
      RECT 24.675 1.18 24.875 2.97 ;
      RECT 25.275 2.695 25.445 3.05 ;
      RECT 19.56 1.06 19.935 1.43 ;
      RECT 19.56 1.18 24.875 1.38 ;
      RECT 23.925 3.54 24.185 3.86 ;
      RECT 23.985 1.835 24.125 3.86 ;
      RECT 23.81 2.395 24.125 2.765 ;
      RECT 23.88 1.95 24.125 2.765 ;
      RECT 23.915 1.835 24.195 2.205 ;
      RECT 23.235 2.42 23.495 2.74 ;
      RECT 22.575 2.51 23.495 2.65 ;
      RECT 22.575 1.57 22.715 2.65 ;
      RECT 19.035 1.86 19.295 2.18 ;
      RECT 19.215 1.57 19.355 2.09 ;
      RECT 19.215 1.57 22.715 1.71 ;
      RECT 22.065 3.26 22.325 3.58 ;
      RECT 22.125 1.85 22.265 3.58 ;
      RECT 22.055 1.85 22.335 2.22 ;
      RECT 19.455 4.01 21.89 4.15 ;
      RECT 21.75 2.7 21.89 4.15 ;
      RECT 19.455 3.63 19.595 4.15 ;
      RECT 19.155 3.63 19.595 3.86 ;
      RECT 16.815 3.63 19.595 3.77 ;
      RECT 19.155 3.54 19.415 3.86 ;
      RECT 16.815 3.35 16.955 3.77 ;
      RECT 16.305 3.26 16.565 3.58 ;
      RECT 16.305 3.35 16.955 3.49 ;
      RECT 16.365 1.86 16.505 3.58 ;
      RECT 21.69 2.7 21.95 3.02 ;
      RECT 16.305 1.86 16.565 2.18 ;
      RECT 21.315 3.54 21.575 3.86 ;
      RECT 21.375 1.95 21.515 3.86 ;
      RECT 21.035 1.95 21.515 2.225 ;
      RECT 20.835 1.855 21.315 2.2 ;
      RECT 20.825 3.49 21.105 3.86 ;
      RECT 20.895 2.395 21.035 3.86 ;
      RECT 20.835 2.395 21.095 3.02 ;
      RECT 20.825 2.395 21.105 2.765 ;
      RECT 19.755 3.54 20.015 3.86 ;
      RECT 19.755 3.35 19.955 3.86 ;
      RECT 19.56 3.35 19.955 3.49 ;
      RECT 19.56 1.86 19.7 3.49 ;
      RECT 19.56 1.86 19.875 2.23 ;
      RECT 19.5 1.86 19.875 2.18 ;
      RECT 17.225 2.955 17.505 3.325 ;
      RECT 18.675 2.98 18.935 3.3 ;
      RECT 17.055 3.07 18.935 3.21 ;
      RECT 17.055 2.955 17.505 3.21 ;
      RECT 16.995 2.395 17.255 3.02 ;
      RECT 16.985 2.395 17.265 2.765 ;
      RECT 18.065 2.395 18.475 2.765 ;
      RECT 17.475 2.42 17.735 2.74 ;
      RECT 17.475 2.51 18.475 2.65 ;
      RECT 12.33 6.655 12.655 6.98 ;
      RECT 11.215 6.745 12.655 6.915 ;
      RECT 11.215 2.395 11.375 6.915 ;
      RECT 11.53 2.365 11.85 2.685 ;
      RECT 11.215 2.395 11.85 2.565 ;
      RECT 10.485 5.86 10.825 6.21 ;
      RECT 10.565 2.705 10.735 6.21 ;
      RECT 10.485 2.705 10.825 3.055 ;
      RECT 9.925 2.7 10.265 3.05 ;
      RECT 9.415 2.77 10.265 2.97 ;
      RECT 9.415 1.18 9.615 2.97 ;
      RECT 10.015 2.695 10.185 3.05 ;
      RECT 4.3 1.06 4.675 1.43 ;
      RECT 4.3 1.18 9.615 1.38 ;
      RECT 8.665 3.54 8.925 3.86 ;
      RECT 8.725 1.835 8.865 3.86 ;
      RECT 8.55 2.395 8.865 2.765 ;
      RECT 8.62 1.95 8.865 2.765 ;
      RECT 8.655 1.835 8.935 2.205 ;
      RECT 7.975 2.42 8.235 2.74 ;
      RECT 7.315 2.51 8.235 2.65 ;
      RECT 7.315 1.57 7.455 2.65 ;
      RECT 3.775 1.86 4.035 2.18 ;
      RECT 3.955 1.57 4.095 2.09 ;
      RECT 3.955 1.57 7.455 1.71 ;
      RECT 6.805 3.26 7.065 3.58 ;
      RECT 6.865 1.85 7.005 3.58 ;
      RECT 6.795 1.85 7.075 2.22 ;
      RECT 4.195 4.01 6.63 4.15 ;
      RECT 6.49 2.7 6.63 4.15 ;
      RECT 4.195 3.63 4.335 4.15 ;
      RECT 3.895 3.63 4.335 3.86 ;
      RECT 1.555 3.63 4.335 3.77 ;
      RECT 3.895 3.54 4.155 3.86 ;
      RECT 1.555 3.35 1.695 3.77 ;
      RECT 1.045 3.26 1.305 3.58 ;
      RECT 1.045 3.35 1.695 3.49 ;
      RECT 1.105 1.86 1.245 3.58 ;
      RECT 6.43 2.7 6.69 3.02 ;
      RECT 1.045 1.86 1.305 2.18 ;
      RECT 6.055 3.54 6.315 3.86 ;
      RECT 6.115 1.95 6.255 3.86 ;
      RECT 5.775 1.95 6.255 2.225 ;
      RECT 5.575 1.855 6.055 2.2 ;
      RECT 5.565 3.49 5.845 3.86 ;
      RECT 5.635 2.395 5.775 3.86 ;
      RECT 5.575 2.395 5.835 3.02 ;
      RECT 5.565 2.395 5.845 2.765 ;
      RECT 4.495 3.54 4.755 3.86 ;
      RECT 4.495 3.35 4.695 3.86 ;
      RECT 4.3 3.35 4.695 3.49 ;
      RECT 4.3 1.86 4.44 3.49 ;
      RECT 4.3 1.86 4.615 2.23 ;
      RECT 4.24 1.86 4.615 2.18 ;
      RECT 1.965 2.955 2.245 3.325 ;
      RECT 3.415 2.98 3.675 3.3 ;
      RECT 1.795 3.07 3.675 3.21 ;
      RECT 1.795 2.955 2.245 3.21 ;
      RECT 1.735 2.395 1.995 3.02 ;
      RECT 1.725 2.395 2.005 2.765 ;
      RECT 2.805 2.395 3.215 2.765 ;
      RECT 2.215 2.42 2.475 2.74 ;
      RECT 2.215 2.51 3.215 2.65 ;
      RECT 66.125 2.395 66.405 2.86 ;
      RECT 65.885 1.86 66.165 2.205 ;
      RECT 64.685 2.395 64.965 2.765 ;
      RECT 50.865 2.395 51.145 2.86 ;
      RECT 50.625 1.86 50.905 2.205 ;
      RECT 49.425 2.395 49.705 2.765 ;
      RECT 35.605 2.395 35.885 2.86 ;
      RECT 35.365 1.86 35.645 2.205 ;
      RECT 34.165 2.395 34.445 2.765 ;
      RECT 20.345 2.395 20.625 2.86 ;
      RECT 20.105 1.86 20.385 2.205 ;
      RECT 18.905 2.395 19.185 2.765 ;
      RECT 5.085 2.395 5.365 2.86 ;
      RECT 4.845 1.86 5.125 2.205 ;
      RECT 3.645 2.395 3.925 2.765 ;
    LAYER via1 ;
      RECT 75.83 1.19 75.98 1.34 ;
      RECT 73.46 6.74 73.61 6.89 ;
      RECT 73.445 2.065 73.595 2.215 ;
      RECT 72.655 2.45 72.805 2.6 ;
      RECT 72.655 6.37 72.805 6.52 ;
      RECT 71.625 2.805 71.775 2.955 ;
      RECT 71.625 5.96 71.775 6.11 ;
      RECT 71.065 2.8 71.215 2.95 ;
      RECT 69.76 1.945 69.91 2.095 ;
      RECT 69.76 3.625 69.91 3.775 ;
      RECT 69.07 2.505 69.22 2.655 ;
      RECT 67.9 1.945 68.05 2.095 ;
      RECT 67.9 3.345 68.05 3.495 ;
      RECT 67.525 2.785 67.675 2.935 ;
      RECT 67.15 3.625 67.3 3.775 ;
      RECT 66.67 1.945 66.82 2.095 ;
      RECT 66.67 2.785 66.82 2.935 ;
      RECT 66.19 2.505 66.34 2.655 ;
      RECT 65.95 1.945 66.1 2.095 ;
      RECT 65.59 3.625 65.74 3.775 ;
      RECT 65.335 1.945 65.485 2.095 ;
      RECT 64.99 3.625 65.14 3.775 ;
      RECT 64.87 1.945 65.02 2.095 ;
      RECT 64.75 2.505 64.9 2.655 ;
      RECT 64.51 3.065 64.66 3.215 ;
      RECT 63.31 2.505 63.46 2.655 ;
      RECT 62.95 1.945 63.1 2.095 ;
      RECT 62.83 2.785 62.98 2.935 ;
      RECT 62.14 1.945 62.29 2.095 ;
      RECT 62.14 3.345 62.29 3.495 ;
      RECT 60.565 1.195 60.715 1.345 ;
      RECT 58.2 6.74 58.35 6.89 ;
      RECT 58.185 2.065 58.335 2.215 ;
      RECT 57.395 2.45 57.545 2.6 ;
      RECT 57.395 6.37 57.545 6.52 ;
      RECT 56.365 2.805 56.515 2.955 ;
      RECT 56.365 5.96 56.515 6.11 ;
      RECT 55.805 2.8 55.955 2.95 ;
      RECT 54.5 1.945 54.65 2.095 ;
      RECT 54.5 3.625 54.65 3.775 ;
      RECT 53.81 2.505 53.96 2.655 ;
      RECT 52.64 1.945 52.79 2.095 ;
      RECT 52.64 3.345 52.79 3.495 ;
      RECT 52.265 2.785 52.415 2.935 ;
      RECT 51.89 3.625 52.04 3.775 ;
      RECT 51.41 1.945 51.56 2.095 ;
      RECT 51.41 2.785 51.56 2.935 ;
      RECT 50.93 2.505 51.08 2.655 ;
      RECT 50.69 1.945 50.84 2.095 ;
      RECT 50.33 3.625 50.48 3.775 ;
      RECT 50.075 1.945 50.225 2.095 ;
      RECT 49.73 3.625 49.88 3.775 ;
      RECT 49.61 1.945 49.76 2.095 ;
      RECT 49.49 2.505 49.64 2.655 ;
      RECT 49.25 3.065 49.4 3.215 ;
      RECT 48.05 2.505 48.2 2.655 ;
      RECT 47.69 1.945 47.84 2.095 ;
      RECT 47.57 2.785 47.72 2.935 ;
      RECT 46.88 1.945 47.03 2.095 ;
      RECT 46.88 3.345 47.03 3.495 ;
      RECT 45.305 1.195 45.455 1.345 ;
      RECT 42.94 6.74 43.09 6.89 ;
      RECT 42.925 2.065 43.075 2.215 ;
      RECT 42.135 2.45 42.285 2.6 ;
      RECT 42.135 6.37 42.285 6.52 ;
      RECT 41.105 2.805 41.255 2.955 ;
      RECT 41.105 5.96 41.255 6.11 ;
      RECT 40.545 2.8 40.695 2.95 ;
      RECT 39.24 1.945 39.39 2.095 ;
      RECT 39.24 3.625 39.39 3.775 ;
      RECT 38.55 2.505 38.7 2.655 ;
      RECT 37.38 1.945 37.53 2.095 ;
      RECT 37.38 3.345 37.53 3.495 ;
      RECT 37.005 2.785 37.155 2.935 ;
      RECT 36.63 3.625 36.78 3.775 ;
      RECT 36.15 1.945 36.3 2.095 ;
      RECT 36.15 2.785 36.3 2.935 ;
      RECT 35.67 2.505 35.82 2.655 ;
      RECT 35.43 1.945 35.58 2.095 ;
      RECT 35.07 3.625 35.22 3.775 ;
      RECT 34.815 1.945 34.965 2.095 ;
      RECT 34.47 3.625 34.62 3.775 ;
      RECT 34.35 1.945 34.5 2.095 ;
      RECT 34.23 2.505 34.38 2.655 ;
      RECT 33.99 3.065 34.14 3.215 ;
      RECT 32.79 2.505 32.94 2.655 ;
      RECT 32.43 1.945 32.58 2.095 ;
      RECT 32.31 2.785 32.46 2.935 ;
      RECT 31.62 1.945 31.77 2.095 ;
      RECT 31.62 3.345 31.77 3.495 ;
      RECT 30.045 1.195 30.195 1.345 ;
      RECT 27.68 6.74 27.83 6.89 ;
      RECT 27.665 2.065 27.815 2.215 ;
      RECT 26.875 2.45 27.025 2.6 ;
      RECT 26.875 6.37 27.025 6.52 ;
      RECT 25.845 2.805 25.995 2.955 ;
      RECT 25.845 5.96 25.995 6.11 ;
      RECT 25.285 2.8 25.435 2.95 ;
      RECT 23.98 1.945 24.13 2.095 ;
      RECT 23.98 3.625 24.13 3.775 ;
      RECT 23.29 2.505 23.44 2.655 ;
      RECT 22.12 1.945 22.27 2.095 ;
      RECT 22.12 3.345 22.27 3.495 ;
      RECT 21.745 2.785 21.895 2.935 ;
      RECT 21.37 3.625 21.52 3.775 ;
      RECT 20.89 1.945 21.04 2.095 ;
      RECT 20.89 2.785 21.04 2.935 ;
      RECT 20.41 2.505 20.56 2.655 ;
      RECT 20.17 1.945 20.32 2.095 ;
      RECT 19.81 3.625 19.96 3.775 ;
      RECT 19.555 1.945 19.705 2.095 ;
      RECT 19.21 3.625 19.36 3.775 ;
      RECT 19.09 1.945 19.24 2.095 ;
      RECT 18.97 2.505 19.12 2.655 ;
      RECT 18.73 3.065 18.88 3.215 ;
      RECT 17.53 2.505 17.68 2.655 ;
      RECT 17.17 1.945 17.32 2.095 ;
      RECT 17.05 2.785 17.2 2.935 ;
      RECT 16.36 1.945 16.51 2.095 ;
      RECT 16.36 3.345 16.51 3.495 ;
      RECT 14.79 1.2 14.94 1.35 ;
      RECT 12.42 6.74 12.57 6.89 ;
      RECT 12.405 2.065 12.555 2.215 ;
      RECT 11.615 2.45 11.765 2.6 ;
      RECT 11.615 6.37 11.765 6.52 ;
      RECT 10.585 2.805 10.735 2.955 ;
      RECT 10.585 5.96 10.735 6.11 ;
      RECT 10.025 2.8 10.175 2.95 ;
      RECT 8.72 1.945 8.87 2.095 ;
      RECT 8.72 3.625 8.87 3.775 ;
      RECT 8.03 2.505 8.18 2.655 ;
      RECT 6.86 1.945 7.01 2.095 ;
      RECT 6.86 3.345 7.01 3.495 ;
      RECT 6.485 2.785 6.635 2.935 ;
      RECT 6.11 3.625 6.26 3.775 ;
      RECT 5.63 1.945 5.78 2.095 ;
      RECT 5.63 2.785 5.78 2.935 ;
      RECT 5.15 2.505 5.3 2.655 ;
      RECT 4.91 1.945 5.06 2.095 ;
      RECT 4.55 3.625 4.7 3.775 ;
      RECT 4.295 1.945 4.445 2.095 ;
      RECT 3.95 3.625 4.1 3.775 ;
      RECT 3.83 1.945 3.98 2.095 ;
      RECT 3.71 2.505 3.86 2.655 ;
      RECT 3.47 3.065 3.62 3.215 ;
      RECT 2.27 2.505 2.42 2.655 ;
      RECT 1.91 1.945 2.06 2.095 ;
      RECT 1.79 2.785 1.94 2.935 ;
      RECT 1.1 1.945 1.25 2.095 ;
      RECT 1.1 3.345 1.25 3.495 ;
    LAYER met1 ;
      RECT 61.79 0 70.53 1.74 ;
      RECT 46.53 0 55.27 1.74 ;
      RECT 31.27 0 40.01 1.74 ;
      RECT 16.01 0 24.75 1.74 ;
      RECT 0.75 0 9.49 1.74 ;
      RECT 0 0 76.3 0.305 ;
      RECT 0 4.14 76.3 4.745 ;
      RECT 61.79 4.135 76.3 4.745 ;
      RECT 46.53 4.135 61.04 4.745 ;
      RECT 31.27 4.135 45.78 4.745 ;
      RECT 16.01 4.135 30.52 4.745 ;
      RECT 0.75 4.135 15.26 4.745 ;
      RECT 61.79 3.98 70.53 4.745 ;
      RECT 46.53 3.98 55.27 4.745 ;
      RECT 31.27 3.98 40.01 4.745 ;
      RECT 16.01 3.98 24.75 4.745 ;
      RECT 0.75 3.98 9.49 4.745 ;
      RECT 75.7 2.365 75.99 2.595 ;
      RECT 75.76 0.885 75.93 2.595 ;
      RECT 75.76 0.885 75.935 1.445 ;
      RECT 75.74 1.09 76.08 1.44 ;
      RECT 75.7 0.885 75.99 1.115 ;
      RECT 75.7 1.085 75.995 1.115 ;
      RECT 75.7 7.765 75.99 7.995 ;
      RECT 75.76 6.285 75.93 7.995 ;
      RECT 75.7 6.285 75.99 6.515 ;
      RECT 75.29 2.735 75.62 2.965 ;
      RECT 75.29 2.765 75.79 2.935 ;
      RECT 75.29 2.395 75.48 2.965 ;
      RECT 74.71 2.365 75 2.595 ;
      RECT 74.71 2.395 75.48 2.565 ;
      RECT 74.77 0.885 74.94 2.595 ;
      RECT 74.71 0.885 75 1.115 ;
      RECT 74.71 7.765 75 7.995 ;
      RECT 74.77 6.285 74.94 7.995 ;
      RECT 74.71 6.285 75 6.515 ;
      RECT 74.71 6.325 75.56 6.485 ;
      RECT 75.39 5.915 75.56 6.485 ;
      RECT 74.71 6.32 75.1 6.485 ;
      RECT 75.33 5.915 75.62 6.145 ;
      RECT 75.33 5.945 75.79 6.115 ;
      RECT 74.34 2.735 74.63 2.965 ;
      RECT 74.34 2.765 74.8 2.935 ;
      RECT 74.4 1.655 74.565 2.965 ;
      RECT 72.915 1.625 73.205 1.855 ;
      RECT 72.915 1.655 74.565 1.825 ;
      RECT 72.975 0.885 73.145 1.855 ;
      RECT 72.915 0.885 73.205 1.115 ;
      RECT 72.915 7.765 73.205 7.995 ;
      RECT 72.975 7.025 73.145 7.995 ;
      RECT 72.975 7.12 74.565 7.29 ;
      RECT 74.395 5.915 74.565 7.29 ;
      RECT 72.915 7.025 73.205 7.255 ;
      RECT 74.34 5.915 74.63 6.145 ;
      RECT 74.34 5.945 74.8 6.115 ;
      RECT 73.345 1.965 73.695 2.315 ;
      RECT 73.175 2.025 73.695 2.195 ;
      RECT 73.37 6.655 73.695 6.98 ;
      RECT 73.345 6.655 73.695 6.885 ;
      RECT 73.175 6.685 73.695 6.855 ;
      RECT 70.965 2.7 71.305 3.05 ;
      RECT 71.055 2.395 71.225 3.05 ;
      RECT 72.57 2.365 72.89 2.685 ;
      RECT 72.54 2.365 72.89 2.595 ;
      RECT 71.055 2.395 72.89 2.565 ;
      RECT 72.57 6.28 72.89 6.605 ;
      RECT 72.54 6.285 72.89 6.515 ;
      RECT 72.37 6.315 72.89 6.485 ;
      RECT 71.525 2.705 71.865 3.055 ;
      RECT 71.525 2.765 72.005 2.935 ;
      RECT 71.525 5.86 71.865 6.21 ;
      RECT 71.525 5.945 72.005 6.115 ;
      RECT 69.675 1.89 69.995 2.15 ;
      RECT 69.24 1.905 69.53 2.135 ;
      RECT 69.24 1.95 69.995 2.09 ;
      RECT 69.675 3.57 69.995 3.83 ;
      RECT 69.24 3.585 69.53 3.815 ;
      RECT 69.24 3.63 69.995 3.77 ;
      RECT 69 3.025 69.29 3.255 ;
      RECT 69 3.07 69.575 3.21 ;
      RECT 69.435 2.93 69.695 3.07 ;
      RECT 69.48 2.745 69.575 3.21 ;
      RECT 69.565 2.735 69.885 3.055 ;
      RECT 67.635 2.93 68.735 3.07 ;
      RECT 67.44 2.73 67.76 2.99 ;
      RECT 68.52 2.745 68.81 2.975 ;
      RECT 67.44 2.745 67.85 2.99 ;
      RECT 67.815 1.89 68.135 2.15 ;
      RECT 68.28 1.905 68.57 2.135 ;
      RECT 67.815 1.95 68.57 2.09 ;
      RECT 65.115 3.155 67.295 3.295 ;
      RECT 67.155 2.165 67.295 3.295 ;
      RECT 65.115 3.07 66.41 3.295 ;
      RECT 66.12 3.025 66.41 3.295 ;
      RECT 65.115 2.79 65.45 3.295 ;
      RECT 65.16 2.745 65.45 3.295 ;
      RECT 68.04 2.465 68.33 2.695 ;
      RECT 67.155 2.37 68.255 2.51 ;
      RECT 67.08 2.165 67.37 2.415 ;
      RECT 67.065 3.57 67.385 3.83 ;
      RECT 67.065 3.585 67.58 3.815 ;
      RECT 65.64 2.465 65.93 2.695 ;
      RECT 65.79 2.07 65.93 2.695 ;
      RECT 65.79 2.07 66.095 2.21 ;
      RECT 66.585 1.89 66.905 2.15 ;
      RECT 65.865 1.89 66.185 2.15 ;
      RECT 66.36 1.905 66.905 2.135 ;
      RECT 65.865 1.95 66.905 2.09 ;
      RECT 65.505 3.57 65.825 3.83 ;
      RECT 65.4 3.585 65.825 3.815 ;
      RECT 63.48 3.025 63.77 3.255 ;
      RECT 63.48 3.025 63.935 3.21 ;
      RECT 63.795 2.55 63.935 3.21 ;
      RECT 63.915 1.95 64.055 2.69 ;
      RECT 64.785 1.89 65.105 2.15 ;
      RECT 63.96 1.905 64.25 2.135 ;
      RECT 63.915 1.95 65.105 2.09 ;
      RECT 64.665 2.45 64.985 2.71 ;
      RECT 64.2 2.465 64.49 2.695 ;
      RECT 64.2 2.51 64.985 2.65 ;
      RECT 64.425 3.01 64.745 3.27 ;
      RECT 64.425 3.025 64.97 3.255 ;
      RECT 63.96 3.585 64.25 3.815 ;
      RECT 63.075 3.465 64.175 3.605 ;
      RECT 63 3.305 63.29 3.535 ;
      RECT 62.28 2.745 62.57 2.975 ;
      RECT 62.355 2.37 62.495 2.975 ;
      RECT 62.355 2.37 62.975 2.51 ;
      RECT 62.835 1.95 62.975 2.51 ;
      RECT 62.595 1.95 62.975 2.21 ;
      RECT 62.865 1.89 63.185 2.15 ;
      RECT 63.48 1.905 63.77 2.135 ;
      RECT 62.595 1.95 63.77 2.09 ;
      RECT 60.44 2.365 60.73 2.595 ;
      RECT 60.5 0.885 60.67 2.595 ;
      RECT 60.475 1.095 60.815 1.445 ;
      RECT 60.44 0.885 60.73 1.115 ;
      RECT 60.44 7.765 60.73 7.995 ;
      RECT 60.5 6.285 60.67 7.995 ;
      RECT 60.44 6.285 60.73 6.515 ;
      RECT 60.03 2.735 60.36 2.965 ;
      RECT 60.03 2.765 60.53 2.935 ;
      RECT 60.03 2.395 60.22 2.965 ;
      RECT 59.45 2.365 59.74 2.595 ;
      RECT 59.45 2.395 60.22 2.565 ;
      RECT 59.51 0.885 59.68 2.595 ;
      RECT 59.45 0.885 59.74 1.115 ;
      RECT 59.45 7.765 59.74 7.995 ;
      RECT 59.51 6.285 59.68 7.995 ;
      RECT 59.45 6.285 59.74 6.515 ;
      RECT 59.45 6.325 60.3 6.485 ;
      RECT 60.13 5.915 60.3 6.485 ;
      RECT 59.45 6.32 59.84 6.485 ;
      RECT 60.07 5.915 60.36 6.145 ;
      RECT 60.07 5.945 60.53 6.115 ;
      RECT 59.08 2.735 59.37 2.965 ;
      RECT 59.08 2.765 59.54 2.935 ;
      RECT 59.14 1.655 59.305 2.965 ;
      RECT 57.655 1.625 57.945 1.855 ;
      RECT 57.655 1.655 59.305 1.825 ;
      RECT 57.715 0.885 57.885 1.855 ;
      RECT 57.655 0.885 57.945 1.115 ;
      RECT 57.655 7.765 57.945 7.995 ;
      RECT 57.715 7.025 57.885 7.995 ;
      RECT 57.715 7.12 59.305 7.29 ;
      RECT 59.135 5.915 59.305 7.29 ;
      RECT 57.655 7.025 57.945 7.255 ;
      RECT 59.08 5.915 59.37 6.145 ;
      RECT 59.08 5.945 59.54 6.115 ;
      RECT 58.085 1.965 58.435 2.315 ;
      RECT 57.915 2.025 58.435 2.195 ;
      RECT 58.11 6.655 58.435 6.98 ;
      RECT 58.085 6.655 58.435 6.885 ;
      RECT 57.915 6.685 58.435 6.855 ;
      RECT 55.705 2.7 56.045 3.05 ;
      RECT 55.795 2.395 55.965 3.05 ;
      RECT 57.31 2.365 57.63 2.685 ;
      RECT 57.28 2.365 57.63 2.595 ;
      RECT 55.795 2.395 57.63 2.565 ;
      RECT 57.31 6.28 57.63 6.605 ;
      RECT 57.28 6.285 57.63 6.515 ;
      RECT 57.11 6.315 57.63 6.485 ;
      RECT 56.265 2.705 56.605 3.055 ;
      RECT 56.265 2.765 56.745 2.935 ;
      RECT 56.265 5.86 56.605 6.21 ;
      RECT 56.265 5.945 56.745 6.115 ;
      RECT 54.415 1.89 54.735 2.15 ;
      RECT 53.98 1.905 54.27 2.135 ;
      RECT 53.98 1.95 54.735 2.09 ;
      RECT 54.415 3.57 54.735 3.83 ;
      RECT 53.98 3.585 54.27 3.815 ;
      RECT 53.98 3.63 54.735 3.77 ;
      RECT 53.74 3.025 54.03 3.255 ;
      RECT 53.74 3.07 54.315 3.21 ;
      RECT 54.175 2.93 54.435 3.07 ;
      RECT 54.22 2.745 54.315 3.21 ;
      RECT 54.305 2.735 54.625 3.055 ;
      RECT 52.375 2.93 53.475 3.07 ;
      RECT 52.18 2.73 52.5 2.99 ;
      RECT 53.26 2.745 53.55 2.975 ;
      RECT 52.18 2.745 52.59 2.99 ;
      RECT 52.555 1.89 52.875 2.15 ;
      RECT 53.02 1.905 53.31 2.135 ;
      RECT 52.555 1.95 53.31 2.09 ;
      RECT 49.855 3.155 52.035 3.295 ;
      RECT 51.895 2.165 52.035 3.295 ;
      RECT 49.855 3.07 51.15 3.295 ;
      RECT 50.86 3.025 51.15 3.295 ;
      RECT 49.855 2.79 50.19 3.295 ;
      RECT 49.9 2.745 50.19 3.295 ;
      RECT 52.78 2.465 53.07 2.695 ;
      RECT 51.895 2.37 52.995 2.51 ;
      RECT 51.82 2.165 52.11 2.415 ;
      RECT 51.805 3.57 52.125 3.83 ;
      RECT 51.805 3.585 52.32 3.815 ;
      RECT 50.38 2.465 50.67 2.695 ;
      RECT 50.53 2.07 50.67 2.695 ;
      RECT 50.53 2.07 50.835 2.21 ;
      RECT 51.325 1.89 51.645 2.15 ;
      RECT 50.605 1.89 50.925 2.15 ;
      RECT 51.1 1.905 51.645 2.135 ;
      RECT 50.605 1.95 51.645 2.09 ;
      RECT 50.245 3.57 50.565 3.83 ;
      RECT 50.14 3.585 50.565 3.815 ;
      RECT 48.22 3.025 48.51 3.255 ;
      RECT 48.22 3.025 48.675 3.21 ;
      RECT 48.535 2.55 48.675 3.21 ;
      RECT 48.655 1.95 48.795 2.69 ;
      RECT 49.525 1.89 49.845 2.15 ;
      RECT 48.7 1.905 48.99 2.135 ;
      RECT 48.655 1.95 49.845 2.09 ;
      RECT 49.405 2.45 49.725 2.71 ;
      RECT 48.94 2.465 49.23 2.695 ;
      RECT 48.94 2.51 49.725 2.65 ;
      RECT 49.165 3.01 49.485 3.27 ;
      RECT 49.165 3.025 49.71 3.255 ;
      RECT 48.7 3.585 48.99 3.815 ;
      RECT 47.815 3.465 48.915 3.605 ;
      RECT 47.74 3.305 48.03 3.535 ;
      RECT 47.02 2.745 47.31 2.975 ;
      RECT 47.095 2.37 47.235 2.975 ;
      RECT 47.095 2.37 47.715 2.51 ;
      RECT 47.575 1.95 47.715 2.51 ;
      RECT 47.335 1.95 47.715 2.21 ;
      RECT 47.605 1.89 47.925 2.15 ;
      RECT 48.22 1.905 48.51 2.135 ;
      RECT 47.335 1.95 48.51 2.09 ;
      RECT 45.18 2.365 45.47 2.595 ;
      RECT 45.24 0.885 45.41 2.595 ;
      RECT 45.215 1.095 45.555 1.445 ;
      RECT 45.18 0.885 45.47 1.115 ;
      RECT 45.18 7.765 45.47 7.995 ;
      RECT 45.24 6.285 45.41 7.995 ;
      RECT 45.18 6.285 45.47 6.515 ;
      RECT 44.77 2.735 45.1 2.965 ;
      RECT 44.77 2.765 45.27 2.935 ;
      RECT 44.77 2.395 44.96 2.965 ;
      RECT 44.19 2.365 44.48 2.595 ;
      RECT 44.19 2.395 44.96 2.565 ;
      RECT 44.25 0.885 44.42 2.595 ;
      RECT 44.19 0.885 44.48 1.115 ;
      RECT 44.19 7.765 44.48 7.995 ;
      RECT 44.25 6.285 44.42 7.995 ;
      RECT 44.19 6.285 44.48 6.515 ;
      RECT 44.19 6.325 45.04 6.485 ;
      RECT 44.87 5.915 45.04 6.485 ;
      RECT 44.19 6.32 44.58 6.485 ;
      RECT 44.81 5.915 45.1 6.145 ;
      RECT 44.81 5.945 45.27 6.115 ;
      RECT 43.82 2.735 44.11 2.965 ;
      RECT 43.82 2.765 44.28 2.935 ;
      RECT 43.88 1.655 44.045 2.965 ;
      RECT 42.395 1.625 42.685 1.855 ;
      RECT 42.395 1.655 44.045 1.825 ;
      RECT 42.455 0.885 42.625 1.855 ;
      RECT 42.395 0.885 42.685 1.115 ;
      RECT 42.395 7.765 42.685 7.995 ;
      RECT 42.455 7.025 42.625 7.995 ;
      RECT 42.455 7.12 44.045 7.29 ;
      RECT 43.875 5.915 44.045 7.29 ;
      RECT 42.395 7.025 42.685 7.255 ;
      RECT 43.82 5.915 44.11 6.145 ;
      RECT 43.82 5.945 44.28 6.115 ;
      RECT 42.825 1.965 43.175 2.315 ;
      RECT 42.655 2.025 43.175 2.195 ;
      RECT 42.85 6.655 43.175 6.98 ;
      RECT 42.825 6.655 43.175 6.885 ;
      RECT 42.655 6.685 43.175 6.855 ;
      RECT 40.445 2.7 40.785 3.05 ;
      RECT 40.535 2.395 40.705 3.05 ;
      RECT 42.05 2.365 42.37 2.685 ;
      RECT 42.02 2.365 42.37 2.595 ;
      RECT 40.535 2.395 42.37 2.565 ;
      RECT 42.05 6.28 42.37 6.605 ;
      RECT 42.02 6.285 42.37 6.515 ;
      RECT 41.85 6.315 42.37 6.485 ;
      RECT 41.005 2.705 41.345 3.055 ;
      RECT 41.005 2.765 41.485 2.935 ;
      RECT 41.005 5.86 41.345 6.21 ;
      RECT 41.005 5.945 41.485 6.115 ;
      RECT 39.155 1.89 39.475 2.15 ;
      RECT 38.72 1.905 39.01 2.135 ;
      RECT 38.72 1.95 39.475 2.09 ;
      RECT 39.155 3.57 39.475 3.83 ;
      RECT 38.72 3.585 39.01 3.815 ;
      RECT 38.72 3.63 39.475 3.77 ;
      RECT 38.48 3.025 38.77 3.255 ;
      RECT 38.48 3.07 39.055 3.21 ;
      RECT 38.915 2.93 39.175 3.07 ;
      RECT 38.96 2.745 39.055 3.21 ;
      RECT 39.045 2.735 39.365 3.055 ;
      RECT 37.115 2.93 38.215 3.07 ;
      RECT 36.92 2.73 37.24 2.99 ;
      RECT 38 2.745 38.29 2.975 ;
      RECT 36.92 2.745 37.33 2.99 ;
      RECT 37.295 1.89 37.615 2.15 ;
      RECT 37.76 1.905 38.05 2.135 ;
      RECT 37.295 1.95 38.05 2.09 ;
      RECT 34.595 3.155 36.775 3.295 ;
      RECT 36.635 2.165 36.775 3.295 ;
      RECT 34.595 3.07 35.89 3.295 ;
      RECT 35.6 3.025 35.89 3.295 ;
      RECT 34.595 2.79 34.93 3.295 ;
      RECT 34.64 2.745 34.93 3.295 ;
      RECT 37.52 2.465 37.81 2.695 ;
      RECT 36.635 2.37 37.735 2.51 ;
      RECT 36.56 2.165 36.85 2.415 ;
      RECT 36.545 3.57 36.865 3.83 ;
      RECT 36.545 3.585 37.06 3.815 ;
      RECT 35.12 2.465 35.41 2.695 ;
      RECT 35.27 2.07 35.41 2.695 ;
      RECT 35.27 2.07 35.575 2.21 ;
      RECT 36.065 1.89 36.385 2.15 ;
      RECT 35.345 1.89 35.665 2.15 ;
      RECT 35.84 1.905 36.385 2.135 ;
      RECT 35.345 1.95 36.385 2.09 ;
      RECT 34.985 3.57 35.305 3.83 ;
      RECT 34.88 3.585 35.305 3.815 ;
      RECT 32.96 3.025 33.25 3.255 ;
      RECT 32.96 3.025 33.415 3.21 ;
      RECT 33.275 2.55 33.415 3.21 ;
      RECT 33.395 1.95 33.535 2.69 ;
      RECT 34.265 1.89 34.585 2.15 ;
      RECT 33.44 1.905 33.73 2.135 ;
      RECT 33.395 1.95 34.585 2.09 ;
      RECT 34.145 2.45 34.465 2.71 ;
      RECT 33.68 2.465 33.97 2.695 ;
      RECT 33.68 2.51 34.465 2.65 ;
      RECT 33.905 3.01 34.225 3.27 ;
      RECT 33.905 3.025 34.45 3.255 ;
      RECT 33.44 3.585 33.73 3.815 ;
      RECT 32.555 3.465 33.655 3.605 ;
      RECT 32.48 3.305 32.77 3.535 ;
      RECT 31.76 2.745 32.05 2.975 ;
      RECT 31.835 2.37 31.975 2.975 ;
      RECT 31.835 2.37 32.455 2.51 ;
      RECT 32.315 1.95 32.455 2.51 ;
      RECT 32.075 1.95 32.455 2.21 ;
      RECT 32.345 1.89 32.665 2.15 ;
      RECT 32.96 1.905 33.25 2.135 ;
      RECT 32.075 1.95 33.25 2.09 ;
      RECT 29.92 2.365 30.21 2.595 ;
      RECT 29.98 0.885 30.15 2.595 ;
      RECT 29.955 1.095 30.295 1.445 ;
      RECT 29.92 0.885 30.21 1.115 ;
      RECT 29.92 7.765 30.21 7.995 ;
      RECT 29.98 6.285 30.15 7.995 ;
      RECT 29.92 6.285 30.21 6.515 ;
      RECT 29.51 2.735 29.84 2.965 ;
      RECT 29.51 2.765 30.01 2.935 ;
      RECT 29.51 2.395 29.7 2.965 ;
      RECT 28.93 2.365 29.22 2.595 ;
      RECT 28.93 2.395 29.7 2.565 ;
      RECT 28.99 0.885 29.16 2.595 ;
      RECT 28.93 0.885 29.22 1.115 ;
      RECT 28.93 7.765 29.22 7.995 ;
      RECT 28.99 6.285 29.16 7.995 ;
      RECT 28.93 6.285 29.22 6.515 ;
      RECT 28.93 6.325 29.78 6.485 ;
      RECT 29.61 5.915 29.78 6.485 ;
      RECT 28.93 6.32 29.32 6.485 ;
      RECT 29.55 5.915 29.84 6.145 ;
      RECT 29.55 5.945 30.01 6.115 ;
      RECT 28.56 2.735 28.85 2.965 ;
      RECT 28.56 2.765 29.02 2.935 ;
      RECT 28.62 1.655 28.785 2.965 ;
      RECT 27.135 1.625 27.425 1.855 ;
      RECT 27.135 1.655 28.785 1.825 ;
      RECT 27.195 0.885 27.365 1.855 ;
      RECT 27.135 0.885 27.425 1.115 ;
      RECT 27.135 7.765 27.425 7.995 ;
      RECT 27.195 7.025 27.365 7.995 ;
      RECT 27.195 7.12 28.785 7.29 ;
      RECT 28.615 5.915 28.785 7.29 ;
      RECT 27.135 7.025 27.425 7.255 ;
      RECT 28.56 5.915 28.85 6.145 ;
      RECT 28.56 5.945 29.02 6.115 ;
      RECT 27.565 1.965 27.915 2.315 ;
      RECT 27.395 2.025 27.915 2.195 ;
      RECT 27.59 6.655 27.915 6.98 ;
      RECT 27.565 6.655 27.915 6.885 ;
      RECT 27.395 6.685 27.915 6.855 ;
      RECT 25.185 2.7 25.525 3.05 ;
      RECT 25.275 2.395 25.445 3.05 ;
      RECT 26.79 2.365 27.11 2.685 ;
      RECT 26.76 2.365 27.11 2.595 ;
      RECT 25.275 2.395 27.11 2.565 ;
      RECT 26.79 6.28 27.11 6.605 ;
      RECT 26.76 6.285 27.11 6.515 ;
      RECT 26.59 6.315 27.11 6.485 ;
      RECT 25.745 2.705 26.085 3.055 ;
      RECT 25.745 2.765 26.225 2.935 ;
      RECT 25.745 5.86 26.085 6.21 ;
      RECT 25.745 5.945 26.225 6.115 ;
      RECT 23.895 1.89 24.215 2.15 ;
      RECT 23.46 1.905 23.75 2.135 ;
      RECT 23.46 1.95 24.215 2.09 ;
      RECT 23.895 3.57 24.215 3.83 ;
      RECT 23.46 3.585 23.75 3.815 ;
      RECT 23.46 3.63 24.215 3.77 ;
      RECT 23.22 3.025 23.51 3.255 ;
      RECT 23.22 3.07 23.795 3.21 ;
      RECT 23.655 2.93 23.915 3.07 ;
      RECT 23.7 2.745 23.795 3.21 ;
      RECT 23.785 2.735 24.105 3.055 ;
      RECT 21.855 2.93 22.955 3.07 ;
      RECT 21.66 2.73 21.98 2.99 ;
      RECT 22.74 2.745 23.03 2.975 ;
      RECT 21.66 2.745 22.07 2.99 ;
      RECT 22.035 1.89 22.355 2.15 ;
      RECT 22.5 1.905 22.79 2.135 ;
      RECT 22.035 1.95 22.79 2.09 ;
      RECT 19.335 3.155 21.515 3.295 ;
      RECT 21.375 2.165 21.515 3.295 ;
      RECT 19.335 3.07 20.63 3.295 ;
      RECT 20.34 3.025 20.63 3.295 ;
      RECT 19.335 2.79 19.67 3.295 ;
      RECT 19.38 2.745 19.67 3.295 ;
      RECT 22.26 2.465 22.55 2.695 ;
      RECT 21.375 2.37 22.475 2.51 ;
      RECT 21.3 2.165 21.59 2.415 ;
      RECT 21.285 3.57 21.605 3.83 ;
      RECT 21.285 3.585 21.8 3.815 ;
      RECT 19.86 2.465 20.15 2.695 ;
      RECT 20.01 2.07 20.15 2.695 ;
      RECT 20.01 2.07 20.315 2.21 ;
      RECT 20.805 1.89 21.125 2.15 ;
      RECT 20.085 1.89 20.405 2.15 ;
      RECT 20.58 1.905 21.125 2.135 ;
      RECT 20.085 1.95 21.125 2.09 ;
      RECT 19.725 3.57 20.045 3.83 ;
      RECT 19.62 3.585 20.045 3.815 ;
      RECT 17.7 3.025 17.99 3.255 ;
      RECT 17.7 3.025 18.155 3.21 ;
      RECT 18.015 2.55 18.155 3.21 ;
      RECT 18.135 1.95 18.275 2.69 ;
      RECT 19.005 1.89 19.325 2.15 ;
      RECT 18.18 1.905 18.47 2.135 ;
      RECT 18.135 1.95 19.325 2.09 ;
      RECT 18.885 2.45 19.205 2.71 ;
      RECT 18.42 2.465 18.71 2.695 ;
      RECT 18.42 2.51 19.205 2.65 ;
      RECT 18.645 3.01 18.965 3.27 ;
      RECT 18.645 3.025 19.19 3.255 ;
      RECT 18.18 3.585 18.47 3.815 ;
      RECT 17.295 3.465 18.395 3.605 ;
      RECT 17.22 3.305 17.51 3.535 ;
      RECT 16.5 2.745 16.79 2.975 ;
      RECT 16.575 2.37 16.715 2.975 ;
      RECT 16.575 2.37 17.195 2.51 ;
      RECT 17.055 1.95 17.195 2.51 ;
      RECT 16.815 1.95 17.195 2.21 ;
      RECT 17.085 1.89 17.405 2.15 ;
      RECT 17.7 1.905 17.99 2.135 ;
      RECT 16.815 1.95 17.99 2.09 ;
      RECT 14.66 2.365 14.95 2.595 ;
      RECT 14.72 0.885 14.89 2.595 ;
      RECT 14.7 1.1 15.04 1.45 ;
      RECT 14.66 0.885 14.95 1.115 ;
      RECT 14.66 7.765 14.95 7.995 ;
      RECT 14.72 6.285 14.89 7.995 ;
      RECT 14.66 6.285 14.95 6.515 ;
      RECT 14.25 2.735 14.58 2.965 ;
      RECT 14.25 2.765 14.75 2.935 ;
      RECT 14.25 2.395 14.44 2.965 ;
      RECT 13.67 2.365 13.96 2.595 ;
      RECT 13.67 2.395 14.44 2.565 ;
      RECT 13.73 0.885 13.9 2.595 ;
      RECT 13.67 0.885 13.96 1.115 ;
      RECT 13.67 7.765 13.96 7.995 ;
      RECT 13.73 6.285 13.9 7.995 ;
      RECT 13.67 6.285 13.96 6.515 ;
      RECT 13.67 6.325 14.52 6.485 ;
      RECT 14.35 5.915 14.52 6.485 ;
      RECT 13.67 6.32 14.06 6.485 ;
      RECT 14.29 5.915 14.58 6.145 ;
      RECT 14.29 5.945 14.75 6.115 ;
      RECT 13.3 2.735 13.59 2.965 ;
      RECT 13.3 2.765 13.76 2.935 ;
      RECT 13.36 1.655 13.525 2.965 ;
      RECT 11.875 1.625 12.165 1.855 ;
      RECT 11.875 1.655 13.525 1.825 ;
      RECT 11.935 0.885 12.105 1.855 ;
      RECT 11.875 0.885 12.165 1.115 ;
      RECT 11.875 7.765 12.165 7.995 ;
      RECT 11.935 7.025 12.105 7.995 ;
      RECT 11.935 7.12 13.525 7.29 ;
      RECT 13.355 5.915 13.525 7.29 ;
      RECT 11.875 7.025 12.165 7.255 ;
      RECT 13.3 5.915 13.59 6.145 ;
      RECT 13.3 5.945 13.76 6.115 ;
      RECT 12.305 1.965 12.655 2.315 ;
      RECT 12.135 2.025 12.655 2.195 ;
      RECT 12.33 6.655 12.655 6.98 ;
      RECT 12.305 6.655 12.655 6.885 ;
      RECT 12.135 6.685 12.655 6.855 ;
      RECT 9.925 2.7 10.265 3.05 ;
      RECT 10.015 2.395 10.185 3.05 ;
      RECT 11.53 2.365 11.85 2.685 ;
      RECT 11.5 2.365 11.85 2.595 ;
      RECT 10.015 2.395 11.85 2.565 ;
      RECT 11.53 6.28 11.85 6.605 ;
      RECT 11.5 6.285 11.85 6.515 ;
      RECT 11.33 6.315 11.85 6.485 ;
      RECT 10.485 2.705 10.825 3.055 ;
      RECT 10.485 2.765 10.965 2.935 ;
      RECT 10.485 5.86 10.825 6.21 ;
      RECT 10.485 5.945 10.965 6.115 ;
      RECT 8.635 1.89 8.955 2.15 ;
      RECT 8.2 1.905 8.49 2.135 ;
      RECT 8.2 1.95 8.955 2.09 ;
      RECT 8.635 3.57 8.955 3.83 ;
      RECT 8.2 3.585 8.49 3.815 ;
      RECT 8.2 3.63 8.955 3.77 ;
      RECT 7.96 3.025 8.25 3.255 ;
      RECT 7.96 3.07 8.535 3.21 ;
      RECT 8.395 2.93 8.655 3.07 ;
      RECT 8.44 2.745 8.535 3.21 ;
      RECT 8.525 2.735 8.845 3.055 ;
      RECT 6.595 2.93 7.695 3.07 ;
      RECT 6.4 2.73 6.72 2.99 ;
      RECT 7.48 2.745 7.77 2.975 ;
      RECT 6.4 2.745 6.81 2.99 ;
      RECT 6.775 1.89 7.095 2.15 ;
      RECT 7.24 1.905 7.53 2.135 ;
      RECT 6.775 1.95 7.53 2.09 ;
      RECT 4.075 3.155 6.255 3.295 ;
      RECT 6.115 2.165 6.255 3.295 ;
      RECT 4.075 3.07 5.37 3.295 ;
      RECT 5.08 3.025 5.37 3.295 ;
      RECT 4.075 2.79 4.41 3.295 ;
      RECT 4.12 2.745 4.41 3.295 ;
      RECT 7 2.465 7.29 2.695 ;
      RECT 6.115 2.37 7.215 2.51 ;
      RECT 6.04 2.165 6.33 2.415 ;
      RECT 6.025 3.57 6.345 3.83 ;
      RECT 6.025 3.585 6.54 3.815 ;
      RECT 4.6 2.465 4.89 2.695 ;
      RECT 4.75 2.07 4.89 2.695 ;
      RECT 4.75 2.07 5.055 2.21 ;
      RECT 5.545 1.89 5.865 2.15 ;
      RECT 4.825 1.89 5.145 2.15 ;
      RECT 5.32 1.905 5.865 2.135 ;
      RECT 4.825 1.95 5.865 2.09 ;
      RECT 4.465 3.57 4.785 3.83 ;
      RECT 4.36 3.585 4.785 3.815 ;
      RECT 2.44 3.025 2.73 3.255 ;
      RECT 2.44 3.025 2.895 3.21 ;
      RECT 2.755 2.55 2.895 3.21 ;
      RECT 2.875 1.95 3.015 2.69 ;
      RECT 3.745 1.89 4.065 2.15 ;
      RECT 2.92 1.905 3.21 2.135 ;
      RECT 2.875 1.95 4.065 2.09 ;
      RECT 3.625 2.45 3.945 2.71 ;
      RECT 3.16 2.465 3.45 2.695 ;
      RECT 3.16 2.51 3.945 2.65 ;
      RECT 3.385 3.01 3.705 3.27 ;
      RECT 3.385 3.025 3.93 3.255 ;
      RECT 2.92 3.585 3.21 3.815 ;
      RECT 2.035 3.465 3.135 3.605 ;
      RECT 1.96 3.305 2.25 3.535 ;
      RECT 1.24 2.745 1.53 2.975 ;
      RECT 1.315 2.37 1.455 2.975 ;
      RECT 1.315 2.37 1.935 2.51 ;
      RECT 1.795 1.95 1.935 2.51 ;
      RECT 1.555 1.95 1.935 2.21 ;
      RECT 1.825 1.89 2.145 2.15 ;
      RECT 2.44 1.905 2.73 2.135 ;
      RECT 1.555 1.95 2.73 2.09 ;
      RECT 0 8.575 76.3 8.88 ;
      RECT 68.985 2.45 69.305 2.71 ;
      RECT 67.815 3.29 68.135 3.55 ;
      RECT 66.585 2.73 66.905 2.99 ;
      RECT 66.105 2.45 66.425 2.71 ;
      RECT 65.25 1.89 65.65 2.15 ;
      RECT 64.905 3.57 65.225 3.83 ;
      RECT 63.225 2.45 63.545 2.71 ;
      RECT 62.745 2.73 63.065 2.99 ;
      RECT 62.055 1.89 62.375 2.15 ;
      RECT 62.055 3.29 62.375 3.55 ;
      RECT 53.725 2.45 54.045 2.71 ;
      RECT 52.555 3.29 52.875 3.55 ;
      RECT 51.325 2.73 51.645 2.99 ;
      RECT 50.845 2.45 51.165 2.71 ;
      RECT 49.99 1.89 50.39 2.15 ;
      RECT 49.645 3.57 49.965 3.83 ;
      RECT 47.965 2.45 48.285 2.71 ;
      RECT 47.485 2.73 47.805 2.99 ;
      RECT 46.795 1.89 47.115 2.15 ;
      RECT 46.795 3.29 47.115 3.55 ;
      RECT 38.465 2.45 38.785 2.71 ;
      RECT 37.295 3.29 37.615 3.55 ;
      RECT 36.065 2.73 36.385 2.99 ;
      RECT 35.585 2.45 35.905 2.71 ;
      RECT 34.73 1.89 35.13 2.15 ;
      RECT 34.385 3.57 34.705 3.83 ;
      RECT 32.705 2.45 33.025 2.71 ;
      RECT 32.225 2.73 32.545 2.99 ;
      RECT 31.535 1.89 31.855 2.15 ;
      RECT 31.535 3.29 31.855 3.55 ;
      RECT 23.205 2.45 23.525 2.71 ;
      RECT 22.035 3.29 22.355 3.55 ;
      RECT 20.805 2.73 21.125 2.99 ;
      RECT 20.325 2.45 20.645 2.71 ;
      RECT 19.47 1.89 19.87 2.15 ;
      RECT 19.125 3.57 19.445 3.83 ;
      RECT 17.445 2.45 17.765 2.71 ;
      RECT 16.965 2.73 17.285 2.99 ;
      RECT 16.275 1.89 16.595 2.15 ;
      RECT 16.275 3.29 16.595 3.55 ;
      RECT 7.945 2.45 8.265 2.71 ;
      RECT 6.775 3.29 7.095 3.55 ;
      RECT 5.545 2.73 5.865 2.99 ;
      RECT 5.065 2.45 5.385 2.71 ;
      RECT 4.21 1.89 4.61 2.15 ;
      RECT 3.865 3.57 4.185 3.83 ;
      RECT 2.185 2.45 2.505 2.71 ;
      RECT 1.705 2.73 2.025 2.99 ;
      RECT 1.015 1.89 1.335 2.15 ;
      RECT 1.015 3.29 1.335 3.55 ;
    LAYER mcon ;
      RECT 75.76 0.915 75.93 1.085 ;
      RECT 75.76 2.395 75.93 2.565 ;
      RECT 75.76 6.315 75.93 6.485 ;
      RECT 75.76 7.795 75.93 7.965 ;
      RECT 75.41 0.105 75.58 0.275 ;
      RECT 75.41 4.165 75.58 4.335 ;
      RECT 75.41 4.545 75.58 4.715 ;
      RECT 75.41 8.605 75.58 8.775 ;
      RECT 75.39 2.765 75.56 2.935 ;
      RECT 75.39 5.945 75.56 6.115 ;
      RECT 74.77 0.915 74.94 1.085 ;
      RECT 74.77 2.395 74.94 2.565 ;
      RECT 74.77 6.315 74.94 6.485 ;
      RECT 74.77 7.795 74.94 7.965 ;
      RECT 74.42 0.105 74.59 0.275 ;
      RECT 74.42 4.165 74.59 4.335 ;
      RECT 74.42 4.545 74.59 4.715 ;
      RECT 74.42 8.605 74.59 8.775 ;
      RECT 74.4 2.765 74.57 2.935 ;
      RECT 74.4 5.945 74.57 6.115 ;
      RECT 73.715 0.105 73.885 0.275 ;
      RECT 73.715 4.165 73.885 4.335 ;
      RECT 73.715 4.545 73.885 4.715 ;
      RECT 73.715 8.605 73.885 8.775 ;
      RECT 73.405 2.025 73.575 2.195 ;
      RECT 73.405 6.685 73.575 6.855 ;
      RECT 73.035 0.105 73.205 0.275 ;
      RECT 73.035 8.605 73.205 8.775 ;
      RECT 72.975 0.915 73.145 1.085 ;
      RECT 72.975 1.655 73.145 1.825 ;
      RECT 72.975 7.055 73.145 7.225 ;
      RECT 72.975 7.795 73.145 7.965 ;
      RECT 72.6 2.395 72.77 2.565 ;
      RECT 72.6 6.315 72.77 6.485 ;
      RECT 72.355 0.105 72.525 0.275 ;
      RECT 72.355 8.605 72.525 8.775 ;
      RECT 71.675 0.105 71.845 0.275 ;
      RECT 71.675 8.605 71.845 8.775 ;
      RECT 71.605 2.765 71.775 2.935 ;
      RECT 71.605 5.945 71.775 6.115 ;
      RECT 70.215 1.415 70.385 1.585 ;
      RECT 70.215 4.135 70.385 4.305 ;
      RECT 69.755 1.415 69.925 1.585 ;
      RECT 69.755 4.135 69.925 4.305 ;
      RECT 69.54 2.775 69.71 2.945 ;
      RECT 69.3 1.935 69.47 2.105 ;
      RECT 69.3 3.615 69.47 3.785 ;
      RECT 69.295 1.415 69.465 1.585 ;
      RECT 69.295 4.135 69.465 4.305 ;
      RECT 69.06 2.495 69.23 2.665 ;
      RECT 69.06 3.055 69.23 3.225 ;
      RECT 68.835 1.415 69.005 1.585 ;
      RECT 68.835 4.135 69.005 4.305 ;
      RECT 68.58 2.775 68.75 2.945 ;
      RECT 68.375 1.415 68.545 1.585 ;
      RECT 68.375 4.135 68.545 4.305 ;
      RECT 68.34 1.935 68.51 2.105 ;
      RECT 68.1 2.495 68.27 2.665 ;
      RECT 67.915 1.415 68.085 1.585 ;
      RECT 67.915 4.135 68.085 4.305 ;
      RECT 67.89 3.335 68.06 3.505 ;
      RECT 67.62 2.775 67.79 2.945 ;
      RECT 67.455 1.415 67.625 1.585 ;
      RECT 67.455 4.135 67.625 4.305 ;
      RECT 67.35 3.615 67.52 3.785 ;
      RECT 67.14 2.195 67.31 2.365 ;
      RECT 66.995 1.415 67.165 1.585 ;
      RECT 66.995 4.135 67.165 4.305 ;
      RECT 66.66 2.775 66.83 2.945 ;
      RECT 66.535 1.415 66.705 1.585 ;
      RECT 66.535 4.135 66.705 4.305 ;
      RECT 66.42 1.935 66.59 2.105 ;
      RECT 66.18 2.495 66.35 2.665 ;
      RECT 66.18 3.055 66.35 3.225 ;
      RECT 66.075 1.415 66.245 1.585 ;
      RECT 66.075 4.135 66.245 4.305 ;
      RECT 65.7 2.495 65.87 2.665 ;
      RECT 65.615 1.415 65.785 1.585 ;
      RECT 65.615 4.135 65.785 4.305 ;
      RECT 65.46 3.615 65.63 3.785 ;
      RECT 65.42 1.935 65.59 2.105 ;
      RECT 65.22 2.775 65.39 2.945 ;
      RECT 65.155 1.415 65.325 1.585 ;
      RECT 65.155 4.135 65.325 4.305 ;
      RECT 64.98 3.615 65.15 3.785 ;
      RECT 64.74 3.055 64.91 3.225 ;
      RECT 64.695 1.415 64.865 1.585 ;
      RECT 64.695 4.135 64.865 4.305 ;
      RECT 64.26 2.495 64.43 2.665 ;
      RECT 64.235 1.415 64.405 1.585 ;
      RECT 64.235 4.135 64.405 4.305 ;
      RECT 64.02 1.935 64.19 2.105 ;
      RECT 64.02 3.615 64.19 3.785 ;
      RECT 63.775 1.415 63.945 1.585 ;
      RECT 63.775 4.135 63.945 4.305 ;
      RECT 63.54 1.935 63.71 2.105 ;
      RECT 63.54 3.055 63.71 3.225 ;
      RECT 63.315 1.415 63.485 1.585 ;
      RECT 63.315 4.135 63.485 4.305 ;
      RECT 63.3 2.495 63.47 2.665 ;
      RECT 63.06 3.335 63.23 3.505 ;
      RECT 62.855 1.415 63.025 1.585 ;
      RECT 62.855 4.135 63.025 4.305 ;
      RECT 62.82 2.775 62.99 2.945 ;
      RECT 62.395 1.415 62.565 1.585 ;
      RECT 62.395 4.135 62.565 4.305 ;
      RECT 62.34 2.775 62.51 2.945 ;
      RECT 62.13 1.935 62.3 2.105 ;
      RECT 62.13 3.335 62.3 3.505 ;
      RECT 61.935 1.415 62.105 1.585 ;
      RECT 61.935 4.135 62.105 4.305 ;
      RECT 60.5 0.915 60.67 1.085 ;
      RECT 60.5 2.395 60.67 2.565 ;
      RECT 60.5 6.315 60.67 6.485 ;
      RECT 60.5 7.795 60.67 7.965 ;
      RECT 60.15 0.105 60.32 0.275 ;
      RECT 60.15 4.165 60.32 4.335 ;
      RECT 60.15 4.545 60.32 4.715 ;
      RECT 60.15 8.605 60.32 8.775 ;
      RECT 60.13 2.765 60.3 2.935 ;
      RECT 60.13 5.945 60.3 6.115 ;
      RECT 59.51 0.915 59.68 1.085 ;
      RECT 59.51 2.395 59.68 2.565 ;
      RECT 59.51 6.315 59.68 6.485 ;
      RECT 59.51 7.795 59.68 7.965 ;
      RECT 59.16 0.105 59.33 0.275 ;
      RECT 59.16 4.165 59.33 4.335 ;
      RECT 59.16 4.545 59.33 4.715 ;
      RECT 59.16 8.605 59.33 8.775 ;
      RECT 59.14 2.765 59.31 2.935 ;
      RECT 59.14 5.945 59.31 6.115 ;
      RECT 58.455 0.105 58.625 0.275 ;
      RECT 58.455 4.165 58.625 4.335 ;
      RECT 58.455 4.545 58.625 4.715 ;
      RECT 58.455 8.605 58.625 8.775 ;
      RECT 58.145 2.025 58.315 2.195 ;
      RECT 58.145 6.685 58.315 6.855 ;
      RECT 57.775 0.105 57.945 0.275 ;
      RECT 57.775 8.605 57.945 8.775 ;
      RECT 57.715 0.915 57.885 1.085 ;
      RECT 57.715 1.655 57.885 1.825 ;
      RECT 57.715 7.055 57.885 7.225 ;
      RECT 57.715 7.795 57.885 7.965 ;
      RECT 57.34 2.395 57.51 2.565 ;
      RECT 57.34 6.315 57.51 6.485 ;
      RECT 57.095 0.105 57.265 0.275 ;
      RECT 57.095 8.605 57.265 8.775 ;
      RECT 56.415 0.105 56.585 0.275 ;
      RECT 56.415 8.605 56.585 8.775 ;
      RECT 56.345 2.765 56.515 2.935 ;
      RECT 56.345 5.945 56.515 6.115 ;
      RECT 54.955 1.415 55.125 1.585 ;
      RECT 54.955 4.135 55.125 4.305 ;
      RECT 54.495 1.415 54.665 1.585 ;
      RECT 54.495 4.135 54.665 4.305 ;
      RECT 54.28 2.775 54.45 2.945 ;
      RECT 54.04 1.935 54.21 2.105 ;
      RECT 54.04 3.615 54.21 3.785 ;
      RECT 54.035 1.415 54.205 1.585 ;
      RECT 54.035 4.135 54.205 4.305 ;
      RECT 53.8 2.495 53.97 2.665 ;
      RECT 53.8 3.055 53.97 3.225 ;
      RECT 53.575 1.415 53.745 1.585 ;
      RECT 53.575 4.135 53.745 4.305 ;
      RECT 53.32 2.775 53.49 2.945 ;
      RECT 53.115 1.415 53.285 1.585 ;
      RECT 53.115 4.135 53.285 4.305 ;
      RECT 53.08 1.935 53.25 2.105 ;
      RECT 52.84 2.495 53.01 2.665 ;
      RECT 52.655 1.415 52.825 1.585 ;
      RECT 52.655 4.135 52.825 4.305 ;
      RECT 52.63 3.335 52.8 3.505 ;
      RECT 52.36 2.775 52.53 2.945 ;
      RECT 52.195 1.415 52.365 1.585 ;
      RECT 52.195 4.135 52.365 4.305 ;
      RECT 52.09 3.615 52.26 3.785 ;
      RECT 51.88 2.195 52.05 2.365 ;
      RECT 51.735 1.415 51.905 1.585 ;
      RECT 51.735 4.135 51.905 4.305 ;
      RECT 51.4 2.775 51.57 2.945 ;
      RECT 51.275 1.415 51.445 1.585 ;
      RECT 51.275 4.135 51.445 4.305 ;
      RECT 51.16 1.935 51.33 2.105 ;
      RECT 50.92 2.495 51.09 2.665 ;
      RECT 50.92 3.055 51.09 3.225 ;
      RECT 50.815 1.415 50.985 1.585 ;
      RECT 50.815 4.135 50.985 4.305 ;
      RECT 50.44 2.495 50.61 2.665 ;
      RECT 50.355 1.415 50.525 1.585 ;
      RECT 50.355 4.135 50.525 4.305 ;
      RECT 50.2 3.615 50.37 3.785 ;
      RECT 50.16 1.935 50.33 2.105 ;
      RECT 49.96 2.775 50.13 2.945 ;
      RECT 49.895 1.415 50.065 1.585 ;
      RECT 49.895 4.135 50.065 4.305 ;
      RECT 49.72 3.615 49.89 3.785 ;
      RECT 49.48 3.055 49.65 3.225 ;
      RECT 49.435 1.415 49.605 1.585 ;
      RECT 49.435 4.135 49.605 4.305 ;
      RECT 49 2.495 49.17 2.665 ;
      RECT 48.975 1.415 49.145 1.585 ;
      RECT 48.975 4.135 49.145 4.305 ;
      RECT 48.76 1.935 48.93 2.105 ;
      RECT 48.76 3.615 48.93 3.785 ;
      RECT 48.515 1.415 48.685 1.585 ;
      RECT 48.515 4.135 48.685 4.305 ;
      RECT 48.28 1.935 48.45 2.105 ;
      RECT 48.28 3.055 48.45 3.225 ;
      RECT 48.055 1.415 48.225 1.585 ;
      RECT 48.055 4.135 48.225 4.305 ;
      RECT 48.04 2.495 48.21 2.665 ;
      RECT 47.8 3.335 47.97 3.505 ;
      RECT 47.595 1.415 47.765 1.585 ;
      RECT 47.595 4.135 47.765 4.305 ;
      RECT 47.56 2.775 47.73 2.945 ;
      RECT 47.135 1.415 47.305 1.585 ;
      RECT 47.135 4.135 47.305 4.305 ;
      RECT 47.08 2.775 47.25 2.945 ;
      RECT 46.87 1.935 47.04 2.105 ;
      RECT 46.87 3.335 47.04 3.505 ;
      RECT 46.675 1.415 46.845 1.585 ;
      RECT 46.675 4.135 46.845 4.305 ;
      RECT 45.24 0.915 45.41 1.085 ;
      RECT 45.24 2.395 45.41 2.565 ;
      RECT 45.24 6.315 45.41 6.485 ;
      RECT 45.24 7.795 45.41 7.965 ;
      RECT 44.89 0.105 45.06 0.275 ;
      RECT 44.89 4.165 45.06 4.335 ;
      RECT 44.89 4.545 45.06 4.715 ;
      RECT 44.89 8.605 45.06 8.775 ;
      RECT 44.87 2.765 45.04 2.935 ;
      RECT 44.87 5.945 45.04 6.115 ;
      RECT 44.25 0.915 44.42 1.085 ;
      RECT 44.25 2.395 44.42 2.565 ;
      RECT 44.25 6.315 44.42 6.485 ;
      RECT 44.25 7.795 44.42 7.965 ;
      RECT 43.9 0.105 44.07 0.275 ;
      RECT 43.9 4.165 44.07 4.335 ;
      RECT 43.9 4.545 44.07 4.715 ;
      RECT 43.9 8.605 44.07 8.775 ;
      RECT 43.88 2.765 44.05 2.935 ;
      RECT 43.88 5.945 44.05 6.115 ;
      RECT 43.195 0.105 43.365 0.275 ;
      RECT 43.195 4.165 43.365 4.335 ;
      RECT 43.195 4.545 43.365 4.715 ;
      RECT 43.195 8.605 43.365 8.775 ;
      RECT 42.885 2.025 43.055 2.195 ;
      RECT 42.885 6.685 43.055 6.855 ;
      RECT 42.515 0.105 42.685 0.275 ;
      RECT 42.515 8.605 42.685 8.775 ;
      RECT 42.455 0.915 42.625 1.085 ;
      RECT 42.455 1.655 42.625 1.825 ;
      RECT 42.455 7.055 42.625 7.225 ;
      RECT 42.455 7.795 42.625 7.965 ;
      RECT 42.08 2.395 42.25 2.565 ;
      RECT 42.08 6.315 42.25 6.485 ;
      RECT 41.835 0.105 42.005 0.275 ;
      RECT 41.835 8.605 42.005 8.775 ;
      RECT 41.155 0.105 41.325 0.275 ;
      RECT 41.155 8.605 41.325 8.775 ;
      RECT 41.085 2.765 41.255 2.935 ;
      RECT 41.085 5.945 41.255 6.115 ;
      RECT 39.695 1.415 39.865 1.585 ;
      RECT 39.695 4.135 39.865 4.305 ;
      RECT 39.235 1.415 39.405 1.585 ;
      RECT 39.235 4.135 39.405 4.305 ;
      RECT 39.02 2.775 39.19 2.945 ;
      RECT 38.78 1.935 38.95 2.105 ;
      RECT 38.78 3.615 38.95 3.785 ;
      RECT 38.775 1.415 38.945 1.585 ;
      RECT 38.775 4.135 38.945 4.305 ;
      RECT 38.54 2.495 38.71 2.665 ;
      RECT 38.54 3.055 38.71 3.225 ;
      RECT 38.315 1.415 38.485 1.585 ;
      RECT 38.315 4.135 38.485 4.305 ;
      RECT 38.06 2.775 38.23 2.945 ;
      RECT 37.855 1.415 38.025 1.585 ;
      RECT 37.855 4.135 38.025 4.305 ;
      RECT 37.82 1.935 37.99 2.105 ;
      RECT 37.58 2.495 37.75 2.665 ;
      RECT 37.395 1.415 37.565 1.585 ;
      RECT 37.395 4.135 37.565 4.305 ;
      RECT 37.37 3.335 37.54 3.505 ;
      RECT 37.1 2.775 37.27 2.945 ;
      RECT 36.935 1.415 37.105 1.585 ;
      RECT 36.935 4.135 37.105 4.305 ;
      RECT 36.83 3.615 37 3.785 ;
      RECT 36.62 2.195 36.79 2.365 ;
      RECT 36.475 1.415 36.645 1.585 ;
      RECT 36.475 4.135 36.645 4.305 ;
      RECT 36.14 2.775 36.31 2.945 ;
      RECT 36.015 1.415 36.185 1.585 ;
      RECT 36.015 4.135 36.185 4.305 ;
      RECT 35.9 1.935 36.07 2.105 ;
      RECT 35.66 2.495 35.83 2.665 ;
      RECT 35.66 3.055 35.83 3.225 ;
      RECT 35.555 1.415 35.725 1.585 ;
      RECT 35.555 4.135 35.725 4.305 ;
      RECT 35.18 2.495 35.35 2.665 ;
      RECT 35.095 1.415 35.265 1.585 ;
      RECT 35.095 4.135 35.265 4.305 ;
      RECT 34.94 3.615 35.11 3.785 ;
      RECT 34.9 1.935 35.07 2.105 ;
      RECT 34.7 2.775 34.87 2.945 ;
      RECT 34.635 1.415 34.805 1.585 ;
      RECT 34.635 4.135 34.805 4.305 ;
      RECT 34.46 3.615 34.63 3.785 ;
      RECT 34.22 3.055 34.39 3.225 ;
      RECT 34.175 1.415 34.345 1.585 ;
      RECT 34.175 4.135 34.345 4.305 ;
      RECT 33.74 2.495 33.91 2.665 ;
      RECT 33.715 1.415 33.885 1.585 ;
      RECT 33.715 4.135 33.885 4.305 ;
      RECT 33.5 1.935 33.67 2.105 ;
      RECT 33.5 3.615 33.67 3.785 ;
      RECT 33.255 1.415 33.425 1.585 ;
      RECT 33.255 4.135 33.425 4.305 ;
      RECT 33.02 1.935 33.19 2.105 ;
      RECT 33.02 3.055 33.19 3.225 ;
      RECT 32.795 1.415 32.965 1.585 ;
      RECT 32.795 4.135 32.965 4.305 ;
      RECT 32.78 2.495 32.95 2.665 ;
      RECT 32.54 3.335 32.71 3.505 ;
      RECT 32.335 1.415 32.505 1.585 ;
      RECT 32.335 4.135 32.505 4.305 ;
      RECT 32.3 2.775 32.47 2.945 ;
      RECT 31.875 1.415 32.045 1.585 ;
      RECT 31.875 4.135 32.045 4.305 ;
      RECT 31.82 2.775 31.99 2.945 ;
      RECT 31.61 1.935 31.78 2.105 ;
      RECT 31.61 3.335 31.78 3.505 ;
      RECT 31.415 1.415 31.585 1.585 ;
      RECT 31.415 4.135 31.585 4.305 ;
      RECT 29.98 0.915 30.15 1.085 ;
      RECT 29.98 2.395 30.15 2.565 ;
      RECT 29.98 6.315 30.15 6.485 ;
      RECT 29.98 7.795 30.15 7.965 ;
      RECT 29.63 0.105 29.8 0.275 ;
      RECT 29.63 4.165 29.8 4.335 ;
      RECT 29.63 4.545 29.8 4.715 ;
      RECT 29.63 8.605 29.8 8.775 ;
      RECT 29.61 2.765 29.78 2.935 ;
      RECT 29.61 5.945 29.78 6.115 ;
      RECT 28.99 0.915 29.16 1.085 ;
      RECT 28.99 2.395 29.16 2.565 ;
      RECT 28.99 6.315 29.16 6.485 ;
      RECT 28.99 7.795 29.16 7.965 ;
      RECT 28.64 0.105 28.81 0.275 ;
      RECT 28.64 4.165 28.81 4.335 ;
      RECT 28.64 4.545 28.81 4.715 ;
      RECT 28.64 8.605 28.81 8.775 ;
      RECT 28.62 2.765 28.79 2.935 ;
      RECT 28.62 5.945 28.79 6.115 ;
      RECT 27.935 0.105 28.105 0.275 ;
      RECT 27.935 4.165 28.105 4.335 ;
      RECT 27.935 4.545 28.105 4.715 ;
      RECT 27.935 8.605 28.105 8.775 ;
      RECT 27.625 2.025 27.795 2.195 ;
      RECT 27.625 6.685 27.795 6.855 ;
      RECT 27.255 0.105 27.425 0.275 ;
      RECT 27.255 8.605 27.425 8.775 ;
      RECT 27.195 0.915 27.365 1.085 ;
      RECT 27.195 1.655 27.365 1.825 ;
      RECT 27.195 7.055 27.365 7.225 ;
      RECT 27.195 7.795 27.365 7.965 ;
      RECT 26.82 2.395 26.99 2.565 ;
      RECT 26.82 6.315 26.99 6.485 ;
      RECT 26.575 0.105 26.745 0.275 ;
      RECT 26.575 8.605 26.745 8.775 ;
      RECT 25.895 0.105 26.065 0.275 ;
      RECT 25.895 8.605 26.065 8.775 ;
      RECT 25.825 2.765 25.995 2.935 ;
      RECT 25.825 5.945 25.995 6.115 ;
      RECT 24.435 1.415 24.605 1.585 ;
      RECT 24.435 4.135 24.605 4.305 ;
      RECT 23.975 1.415 24.145 1.585 ;
      RECT 23.975 4.135 24.145 4.305 ;
      RECT 23.76 2.775 23.93 2.945 ;
      RECT 23.52 1.935 23.69 2.105 ;
      RECT 23.52 3.615 23.69 3.785 ;
      RECT 23.515 1.415 23.685 1.585 ;
      RECT 23.515 4.135 23.685 4.305 ;
      RECT 23.28 2.495 23.45 2.665 ;
      RECT 23.28 3.055 23.45 3.225 ;
      RECT 23.055 1.415 23.225 1.585 ;
      RECT 23.055 4.135 23.225 4.305 ;
      RECT 22.8 2.775 22.97 2.945 ;
      RECT 22.595 1.415 22.765 1.585 ;
      RECT 22.595 4.135 22.765 4.305 ;
      RECT 22.56 1.935 22.73 2.105 ;
      RECT 22.32 2.495 22.49 2.665 ;
      RECT 22.135 1.415 22.305 1.585 ;
      RECT 22.135 4.135 22.305 4.305 ;
      RECT 22.11 3.335 22.28 3.505 ;
      RECT 21.84 2.775 22.01 2.945 ;
      RECT 21.675 1.415 21.845 1.585 ;
      RECT 21.675 4.135 21.845 4.305 ;
      RECT 21.57 3.615 21.74 3.785 ;
      RECT 21.36 2.195 21.53 2.365 ;
      RECT 21.215 1.415 21.385 1.585 ;
      RECT 21.215 4.135 21.385 4.305 ;
      RECT 20.88 2.775 21.05 2.945 ;
      RECT 20.755 1.415 20.925 1.585 ;
      RECT 20.755 4.135 20.925 4.305 ;
      RECT 20.64 1.935 20.81 2.105 ;
      RECT 20.4 2.495 20.57 2.665 ;
      RECT 20.4 3.055 20.57 3.225 ;
      RECT 20.295 1.415 20.465 1.585 ;
      RECT 20.295 4.135 20.465 4.305 ;
      RECT 19.92 2.495 20.09 2.665 ;
      RECT 19.835 1.415 20.005 1.585 ;
      RECT 19.835 4.135 20.005 4.305 ;
      RECT 19.68 3.615 19.85 3.785 ;
      RECT 19.64 1.935 19.81 2.105 ;
      RECT 19.44 2.775 19.61 2.945 ;
      RECT 19.375 1.415 19.545 1.585 ;
      RECT 19.375 4.135 19.545 4.305 ;
      RECT 19.2 3.615 19.37 3.785 ;
      RECT 18.96 3.055 19.13 3.225 ;
      RECT 18.915 1.415 19.085 1.585 ;
      RECT 18.915 4.135 19.085 4.305 ;
      RECT 18.48 2.495 18.65 2.665 ;
      RECT 18.455 1.415 18.625 1.585 ;
      RECT 18.455 4.135 18.625 4.305 ;
      RECT 18.24 1.935 18.41 2.105 ;
      RECT 18.24 3.615 18.41 3.785 ;
      RECT 17.995 1.415 18.165 1.585 ;
      RECT 17.995 4.135 18.165 4.305 ;
      RECT 17.76 1.935 17.93 2.105 ;
      RECT 17.76 3.055 17.93 3.225 ;
      RECT 17.535 1.415 17.705 1.585 ;
      RECT 17.535 4.135 17.705 4.305 ;
      RECT 17.52 2.495 17.69 2.665 ;
      RECT 17.28 3.335 17.45 3.505 ;
      RECT 17.075 1.415 17.245 1.585 ;
      RECT 17.075 4.135 17.245 4.305 ;
      RECT 17.04 2.775 17.21 2.945 ;
      RECT 16.615 1.415 16.785 1.585 ;
      RECT 16.615 4.135 16.785 4.305 ;
      RECT 16.56 2.775 16.73 2.945 ;
      RECT 16.35 1.935 16.52 2.105 ;
      RECT 16.35 3.335 16.52 3.505 ;
      RECT 16.155 1.415 16.325 1.585 ;
      RECT 16.155 4.135 16.325 4.305 ;
      RECT 14.72 0.915 14.89 1.085 ;
      RECT 14.72 2.395 14.89 2.565 ;
      RECT 14.72 6.315 14.89 6.485 ;
      RECT 14.72 7.795 14.89 7.965 ;
      RECT 14.37 0.105 14.54 0.275 ;
      RECT 14.37 4.165 14.54 4.335 ;
      RECT 14.37 4.545 14.54 4.715 ;
      RECT 14.37 8.605 14.54 8.775 ;
      RECT 14.35 2.765 14.52 2.935 ;
      RECT 14.35 5.945 14.52 6.115 ;
      RECT 13.73 0.915 13.9 1.085 ;
      RECT 13.73 2.395 13.9 2.565 ;
      RECT 13.73 6.315 13.9 6.485 ;
      RECT 13.73 7.795 13.9 7.965 ;
      RECT 13.38 0.105 13.55 0.275 ;
      RECT 13.38 4.165 13.55 4.335 ;
      RECT 13.38 4.545 13.55 4.715 ;
      RECT 13.38 8.605 13.55 8.775 ;
      RECT 13.36 2.765 13.53 2.935 ;
      RECT 13.36 5.945 13.53 6.115 ;
      RECT 12.675 0.105 12.845 0.275 ;
      RECT 12.675 4.165 12.845 4.335 ;
      RECT 12.675 4.545 12.845 4.715 ;
      RECT 12.675 8.605 12.845 8.775 ;
      RECT 12.365 2.025 12.535 2.195 ;
      RECT 12.365 6.685 12.535 6.855 ;
      RECT 11.995 0.105 12.165 0.275 ;
      RECT 11.995 8.605 12.165 8.775 ;
      RECT 11.935 0.915 12.105 1.085 ;
      RECT 11.935 1.655 12.105 1.825 ;
      RECT 11.935 7.055 12.105 7.225 ;
      RECT 11.935 7.795 12.105 7.965 ;
      RECT 11.56 2.395 11.73 2.565 ;
      RECT 11.56 6.315 11.73 6.485 ;
      RECT 11.315 0.105 11.485 0.275 ;
      RECT 11.315 8.605 11.485 8.775 ;
      RECT 10.635 0.105 10.805 0.275 ;
      RECT 10.635 8.605 10.805 8.775 ;
      RECT 10.565 2.765 10.735 2.935 ;
      RECT 10.565 5.945 10.735 6.115 ;
      RECT 9.175 1.415 9.345 1.585 ;
      RECT 9.175 4.135 9.345 4.305 ;
      RECT 8.715 1.415 8.885 1.585 ;
      RECT 8.715 4.135 8.885 4.305 ;
      RECT 8.5 2.775 8.67 2.945 ;
      RECT 8.26 1.935 8.43 2.105 ;
      RECT 8.26 3.615 8.43 3.785 ;
      RECT 8.255 1.415 8.425 1.585 ;
      RECT 8.255 4.135 8.425 4.305 ;
      RECT 8.02 2.495 8.19 2.665 ;
      RECT 8.02 3.055 8.19 3.225 ;
      RECT 7.795 1.415 7.965 1.585 ;
      RECT 7.795 4.135 7.965 4.305 ;
      RECT 7.54 2.775 7.71 2.945 ;
      RECT 7.335 1.415 7.505 1.585 ;
      RECT 7.335 4.135 7.505 4.305 ;
      RECT 7.3 1.935 7.47 2.105 ;
      RECT 7.06 2.495 7.23 2.665 ;
      RECT 6.875 1.415 7.045 1.585 ;
      RECT 6.875 4.135 7.045 4.305 ;
      RECT 6.85 3.335 7.02 3.505 ;
      RECT 6.58 2.775 6.75 2.945 ;
      RECT 6.415 1.415 6.585 1.585 ;
      RECT 6.415 4.135 6.585 4.305 ;
      RECT 6.31 3.615 6.48 3.785 ;
      RECT 6.1 2.195 6.27 2.365 ;
      RECT 5.955 1.415 6.125 1.585 ;
      RECT 5.955 4.135 6.125 4.305 ;
      RECT 5.62 2.775 5.79 2.945 ;
      RECT 5.495 1.415 5.665 1.585 ;
      RECT 5.495 4.135 5.665 4.305 ;
      RECT 5.38 1.935 5.55 2.105 ;
      RECT 5.14 2.495 5.31 2.665 ;
      RECT 5.14 3.055 5.31 3.225 ;
      RECT 5.035 1.415 5.205 1.585 ;
      RECT 5.035 4.135 5.205 4.305 ;
      RECT 4.66 2.495 4.83 2.665 ;
      RECT 4.575 1.415 4.745 1.585 ;
      RECT 4.575 4.135 4.745 4.305 ;
      RECT 4.42 3.615 4.59 3.785 ;
      RECT 4.38 1.935 4.55 2.105 ;
      RECT 4.18 2.775 4.35 2.945 ;
      RECT 4.115 1.415 4.285 1.585 ;
      RECT 4.115 4.135 4.285 4.305 ;
      RECT 3.94 3.615 4.11 3.785 ;
      RECT 3.7 3.055 3.87 3.225 ;
      RECT 3.655 1.415 3.825 1.585 ;
      RECT 3.655 4.135 3.825 4.305 ;
      RECT 3.22 2.495 3.39 2.665 ;
      RECT 3.195 1.415 3.365 1.585 ;
      RECT 3.195 4.135 3.365 4.305 ;
      RECT 2.98 1.935 3.15 2.105 ;
      RECT 2.98 3.615 3.15 3.785 ;
      RECT 2.735 1.415 2.905 1.585 ;
      RECT 2.735 4.135 2.905 4.305 ;
      RECT 2.5 1.935 2.67 2.105 ;
      RECT 2.5 3.055 2.67 3.225 ;
      RECT 2.275 1.415 2.445 1.585 ;
      RECT 2.275 4.135 2.445 4.305 ;
      RECT 2.26 2.495 2.43 2.665 ;
      RECT 2.02 3.335 2.19 3.505 ;
      RECT 1.815 1.415 1.985 1.585 ;
      RECT 1.815 4.135 1.985 4.305 ;
      RECT 1.78 2.775 1.95 2.945 ;
      RECT 1.355 1.415 1.525 1.585 ;
      RECT 1.355 4.135 1.525 4.305 ;
      RECT 1.3 2.775 1.47 2.945 ;
      RECT 1.09 1.935 1.26 2.105 ;
      RECT 1.09 3.335 1.26 3.505 ;
      RECT 0.895 1.415 1.065 1.585 ;
      RECT 0.895 4.135 1.065 4.305 ;
    LAYER li ;
      RECT 69.76 0 69.93 2.085 ;
      RECT 68.82 0 68.99 2.085 ;
      RECT 67.86 0 68.03 2.085 ;
      RECT 65.94 0 66.11 2.085 ;
      RECT 64.98 0 65.15 2.085 ;
      RECT 63.06 0 63.23 2.085 ;
      RECT 54.5 0 54.67 2.085 ;
      RECT 53.56 0 53.73 2.085 ;
      RECT 52.6 0 52.77 2.085 ;
      RECT 50.68 0 50.85 2.085 ;
      RECT 49.72 0 49.89 2.085 ;
      RECT 47.8 0 47.97 2.085 ;
      RECT 39.24 0 39.41 2.085 ;
      RECT 38.3 0 38.47 2.085 ;
      RECT 37.34 0 37.51 2.085 ;
      RECT 35.42 0 35.59 2.085 ;
      RECT 34.46 0 34.63 2.085 ;
      RECT 32.54 0 32.71 2.085 ;
      RECT 23.98 0 24.15 2.085 ;
      RECT 23.04 0 23.21 2.085 ;
      RECT 22.08 0 22.25 2.085 ;
      RECT 20.16 0 20.33 2.085 ;
      RECT 19.2 0 19.37 2.085 ;
      RECT 17.28 0 17.45 2.085 ;
      RECT 8.72 0 8.89 2.085 ;
      RECT 7.78 0 7.95 2.085 ;
      RECT 6.82 0 6.99 2.085 ;
      RECT 4.9 0 5.07 2.085 ;
      RECT 3.94 0 4.11 2.085 ;
      RECT 2.02 0 2.19 2.085 ;
      RECT 66.815 0 67.01 1.595 ;
      RECT 63.06 0 63.335 1.595 ;
      RECT 51.555 0 51.75 1.595 ;
      RECT 47.8 0 48.075 1.595 ;
      RECT 36.295 0 36.49 1.595 ;
      RECT 32.54 0 32.815 1.595 ;
      RECT 21.035 0 21.23 1.595 ;
      RECT 17.28 0 17.555 1.595 ;
      RECT 5.775 0 5.97 1.595 ;
      RECT 2.02 0 2.295 1.595 ;
      RECT 61.79 0 70.53 1.585 ;
      RECT 46.53 0 55.27 1.585 ;
      RECT 31.27 0 40.01 1.585 ;
      RECT 16.01 0 24.75 1.585 ;
      RECT 0.75 0 9.49 1.585 ;
      RECT 75.33 0 75.5 0.935 ;
      RECT 74.34 0 74.51 0.935 ;
      RECT 71.595 0 71.765 0.935 ;
      RECT 60.07 0 60.24 0.935 ;
      RECT 59.08 0 59.25 0.935 ;
      RECT 56.335 0 56.505 0.935 ;
      RECT 44.81 0 44.98 0.935 ;
      RECT 43.82 0 43.99 0.935 ;
      RECT 41.075 0 41.245 0.935 ;
      RECT 29.55 0 29.72 0.935 ;
      RECT 28.56 0 28.73 0.935 ;
      RECT 25.815 0 25.985 0.935 ;
      RECT 14.29 0 14.46 0.935 ;
      RECT 13.3 0 13.47 0.935 ;
      RECT 10.555 0 10.725 0.935 ;
      RECT 0 0 76.3 0.305 ;
      RECT 75.33 3.405 75.5 5.475 ;
      RECT 74.34 3.405 74.51 5.475 ;
      RECT 71.595 3.405 71.765 5.475 ;
      RECT 60.07 3.405 60.24 5.475 ;
      RECT 59.08 3.405 59.25 5.475 ;
      RECT 56.335 3.405 56.505 5.475 ;
      RECT 44.81 3.405 44.98 5.475 ;
      RECT 43.82 3.405 43.99 5.475 ;
      RECT 41.075 3.405 41.245 5.475 ;
      RECT 29.55 3.405 29.72 5.475 ;
      RECT 28.56 3.405 28.73 5.475 ;
      RECT 25.815 3.405 25.985 5.475 ;
      RECT 14.29 3.405 14.46 5.475 ;
      RECT 13.3 3.405 13.47 5.475 ;
      RECT 10.555 3.405 10.725 5.475 ;
      RECT 0 4.14 76.3 4.745 ;
      RECT 61.79 4.135 76.3 4.745 ;
      RECT 46.53 4.135 61.04 4.745 ;
      RECT 31.27 4.135 45.78 4.745 ;
      RECT 16.01 4.135 30.52 4.745 ;
      RECT 0.75 4.135 15.26 4.745 ;
      RECT 68.82 3.635 68.99 4.745 ;
      RECT 66.9 3.635 67.07 4.745 ;
      RECT 65.96 3.635 66.13 4.745 ;
      RECT 64.5 3.635 64.67 4.745 ;
      RECT 62.58 3.635 62.75 4.745 ;
      RECT 53.56 3.635 53.73 4.745 ;
      RECT 51.64 3.635 51.81 4.745 ;
      RECT 50.7 3.635 50.87 4.745 ;
      RECT 49.24 3.635 49.41 4.745 ;
      RECT 47.32 3.635 47.49 4.745 ;
      RECT 38.3 3.635 38.47 4.745 ;
      RECT 36.38 3.635 36.55 4.745 ;
      RECT 35.44 3.635 35.61 4.745 ;
      RECT 33.98 3.635 34.15 4.745 ;
      RECT 32.06 3.635 32.23 4.745 ;
      RECT 23.04 3.635 23.21 4.745 ;
      RECT 21.12 3.635 21.29 4.745 ;
      RECT 20.18 3.635 20.35 4.745 ;
      RECT 18.72 3.635 18.89 4.745 ;
      RECT 16.8 3.635 16.97 4.745 ;
      RECT 7.78 3.635 7.95 4.745 ;
      RECT 5.86 3.635 6.03 4.745 ;
      RECT 4.92 3.635 5.09 4.745 ;
      RECT 3.46 3.635 3.63 4.745 ;
      RECT 1.54 3.635 1.71 4.745 ;
      RECT 0 8.575 76.3 8.88 ;
      RECT 75.33 7.945 75.5 8.88 ;
      RECT 74.34 7.945 74.51 8.88 ;
      RECT 71.595 7.945 71.765 8.88 ;
      RECT 60.07 7.945 60.24 8.88 ;
      RECT 59.08 7.945 59.25 8.88 ;
      RECT 56.335 7.945 56.505 8.88 ;
      RECT 44.81 7.945 44.98 8.88 ;
      RECT 43.82 7.945 43.99 8.88 ;
      RECT 41.075 7.945 41.245 8.88 ;
      RECT 29.55 7.945 29.72 8.88 ;
      RECT 28.56 7.945 28.73 8.88 ;
      RECT 25.815 7.945 25.985 8.88 ;
      RECT 14.29 7.945 14.46 8.88 ;
      RECT 13.3 7.945 13.47 8.88 ;
      RECT 10.555 7.945 10.725 8.88 ;
      RECT 75.39 1.74 75.56 2.935 ;
      RECT 75.39 1.74 75.855 1.91 ;
      RECT 75.39 6.97 75.855 7.14 ;
      RECT 75.39 5.945 75.56 7.14 ;
      RECT 74.4 1.74 74.57 2.935 ;
      RECT 74.4 1.74 74.865 1.91 ;
      RECT 74.4 6.97 74.865 7.14 ;
      RECT 74.4 5.945 74.57 7.14 ;
      RECT 72.545 2.635 72.715 3.865 ;
      RECT 72.6 0.855 72.77 2.805 ;
      RECT 72.545 0.575 72.715 1.025 ;
      RECT 72.545 7.855 72.715 8.305 ;
      RECT 72.6 6.075 72.77 8.025 ;
      RECT 72.545 5.015 72.715 6.245 ;
      RECT 72.025 0.575 72.195 3.865 ;
      RECT 72.025 2.075 72.43 2.405 ;
      RECT 72.025 1.235 72.43 1.565 ;
      RECT 72.025 5.015 72.195 8.305 ;
      RECT 72.025 7.315 72.43 7.645 ;
      RECT 72.025 6.475 72.43 6.805 ;
      RECT 69.3 3.615 69.815 3.785 ;
      RECT 69.645 3.225 69.815 3.785 ;
      RECT 69.75 3.145 69.92 3.475 ;
      RECT 69.54 2.535 69.815 2.945 ;
      RECT 69.42 2.535 69.815 2.745 ;
      RECT 67.89 3.145 68.06 3.505 ;
      RECT 67.89 3.225 69.23 3.395 ;
      RECT 69.06 3.055 69.23 3.395 ;
      RECT 67.62 2.575 67.79 2.945 ;
      RECT 67.14 2.575 67.79 2.845 ;
      RECT 67.06 2.575 67.87 2.745 ;
      RECT 66.42 1.815 66.59 2.105 ;
      RECT 66.42 1.815 67.66 1.985 ;
      RECT 67.14 2.155 67.31 2.365 ;
      RECT 66.78 2.155 67.31 2.325 ;
      RECT 66.18 3.225 66.67 3.395 ;
      RECT 66.18 3.055 66.35 3.395 ;
      RECT 65.46 3.225 65.63 3.785 ;
      RECT 65.35 3.225 65.68 3.395 ;
      RECT 65.42 1.835 65.59 2.105 ;
      RECT 65.46 1.755 65.63 2.085 ;
      RECT 65.325 1.835 65.63 2.055 ;
      RECT 63.9 3.225 64.19 3.785 ;
      RECT 64.02 3.145 64.19 3.785 ;
      RECT 63.66 2.575 64.03 2.745 ;
      RECT 63.66 1.935 63.83 2.745 ;
      RECT 63.54 1.935 63.83 2.105 ;
      RECT 60.13 1.74 60.3 2.935 ;
      RECT 60.13 1.74 60.595 1.91 ;
      RECT 60.13 6.97 60.595 7.14 ;
      RECT 60.13 5.945 60.3 7.14 ;
      RECT 59.14 1.74 59.31 2.935 ;
      RECT 59.14 1.74 59.605 1.91 ;
      RECT 59.14 6.97 59.605 7.14 ;
      RECT 59.14 5.945 59.31 7.14 ;
      RECT 57.285 2.635 57.455 3.865 ;
      RECT 57.34 0.855 57.51 2.805 ;
      RECT 57.285 0.575 57.455 1.025 ;
      RECT 57.285 7.855 57.455 8.305 ;
      RECT 57.34 6.075 57.51 8.025 ;
      RECT 57.285 5.015 57.455 6.245 ;
      RECT 56.765 0.575 56.935 3.865 ;
      RECT 56.765 2.075 57.17 2.405 ;
      RECT 56.765 1.235 57.17 1.565 ;
      RECT 56.765 5.015 56.935 8.305 ;
      RECT 56.765 7.315 57.17 7.645 ;
      RECT 56.765 6.475 57.17 6.805 ;
      RECT 54.04 3.615 54.555 3.785 ;
      RECT 54.385 3.225 54.555 3.785 ;
      RECT 54.49 3.145 54.66 3.475 ;
      RECT 54.28 2.535 54.555 2.945 ;
      RECT 54.16 2.535 54.555 2.745 ;
      RECT 52.63 3.145 52.8 3.505 ;
      RECT 52.63 3.225 53.97 3.395 ;
      RECT 53.8 3.055 53.97 3.395 ;
      RECT 52.36 2.575 52.53 2.945 ;
      RECT 51.88 2.575 52.53 2.845 ;
      RECT 51.8 2.575 52.61 2.745 ;
      RECT 51.16 1.815 51.33 2.105 ;
      RECT 51.16 1.815 52.4 1.985 ;
      RECT 51.88 2.155 52.05 2.365 ;
      RECT 51.52 2.155 52.05 2.325 ;
      RECT 50.92 3.225 51.41 3.395 ;
      RECT 50.92 3.055 51.09 3.395 ;
      RECT 50.2 3.225 50.37 3.785 ;
      RECT 50.09 3.225 50.42 3.395 ;
      RECT 50.16 1.835 50.33 2.105 ;
      RECT 50.2 1.755 50.37 2.085 ;
      RECT 50.065 1.835 50.37 2.055 ;
      RECT 48.64 3.225 48.93 3.785 ;
      RECT 48.76 3.145 48.93 3.785 ;
      RECT 48.4 2.575 48.77 2.745 ;
      RECT 48.4 1.935 48.57 2.745 ;
      RECT 48.28 1.935 48.57 2.105 ;
      RECT 44.87 1.74 45.04 2.935 ;
      RECT 44.87 1.74 45.335 1.91 ;
      RECT 44.87 6.97 45.335 7.14 ;
      RECT 44.87 5.945 45.04 7.14 ;
      RECT 43.88 1.74 44.05 2.935 ;
      RECT 43.88 1.74 44.345 1.91 ;
      RECT 43.88 6.97 44.345 7.14 ;
      RECT 43.88 5.945 44.05 7.14 ;
      RECT 42.025 2.635 42.195 3.865 ;
      RECT 42.08 0.855 42.25 2.805 ;
      RECT 42.025 0.575 42.195 1.025 ;
      RECT 42.025 7.855 42.195 8.305 ;
      RECT 42.08 6.075 42.25 8.025 ;
      RECT 42.025 5.015 42.195 6.245 ;
      RECT 41.505 0.575 41.675 3.865 ;
      RECT 41.505 2.075 41.91 2.405 ;
      RECT 41.505 1.235 41.91 1.565 ;
      RECT 41.505 5.015 41.675 8.305 ;
      RECT 41.505 7.315 41.91 7.645 ;
      RECT 41.505 6.475 41.91 6.805 ;
      RECT 38.78 3.615 39.295 3.785 ;
      RECT 39.125 3.225 39.295 3.785 ;
      RECT 39.23 3.145 39.4 3.475 ;
      RECT 39.02 2.535 39.295 2.945 ;
      RECT 38.9 2.535 39.295 2.745 ;
      RECT 37.37 3.145 37.54 3.505 ;
      RECT 37.37 3.225 38.71 3.395 ;
      RECT 38.54 3.055 38.71 3.395 ;
      RECT 37.1 2.575 37.27 2.945 ;
      RECT 36.62 2.575 37.27 2.845 ;
      RECT 36.54 2.575 37.35 2.745 ;
      RECT 35.9 1.815 36.07 2.105 ;
      RECT 35.9 1.815 37.14 1.985 ;
      RECT 36.62 2.155 36.79 2.365 ;
      RECT 36.26 2.155 36.79 2.325 ;
      RECT 35.66 3.225 36.15 3.395 ;
      RECT 35.66 3.055 35.83 3.395 ;
      RECT 34.94 3.225 35.11 3.785 ;
      RECT 34.83 3.225 35.16 3.395 ;
      RECT 34.9 1.835 35.07 2.105 ;
      RECT 34.94 1.755 35.11 2.085 ;
      RECT 34.805 1.835 35.11 2.055 ;
      RECT 33.38 3.225 33.67 3.785 ;
      RECT 33.5 3.145 33.67 3.785 ;
      RECT 33.14 2.575 33.51 2.745 ;
      RECT 33.14 1.935 33.31 2.745 ;
      RECT 33.02 1.935 33.31 2.105 ;
      RECT 29.61 1.74 29.78 2.935 ;
      RECT 29.61 1.74 30.075 1.91 ;
      RECT 29.61 6.97 30.075 7.14 ;
      RECT 29.61 5.945 29.78 7.14 ;
      RECT 28.62 1.74 28.79 2.935 ;
      RECT 28.62 1.74 29.085 1.91 ;
      RECT 28.62 6.97 29.085 7.14 ;
      RECT 28.62 5.945 28.79 7.14 ;
      RECT 26.765 2.635 26.935 3.865 ;
      RECT 26.82 0.855 26.99 2.805 ;
      RECT 26.765 0.575 26.935 1.025 ;
      RECT 26.765 7.855 26.935 8.305 ;
      RECT 26.82 6.075 26.99 8.025 ;
      RECT 26.765 5.015 26.935 6.245 ;
      RECT 26.245 0.575 26.415 3.865 ;
      RECT 26.245 2.075 26.65 2.405 ;
      RECT 26.245 1.235 26.65 1.565 ;
      RECT 26.245 5.015 26.415 8.305 ;
      RECT 26.245 7.315 26.65 7.645 ;
      RECT 26.245 6.475 26.65 6.805 ;
      RECT 23.52 3.615 24.035 3.785 ;
      RECT 23.865 3.225 24.035 3.785 ;
      RECT 23.97 3.145 24.14 3.475 ;
      RECT 23.76 2.535 24.035 2.945 ;
      RECT 23.64 2.535 24.035 2.745 ;
      RECT 22.11 3.145 22.28 3.505 ;
      RECT 22.11 3.225 23.45 3.395 ;
      RECT 23.28 3.055 23.45 3.395 ;
      RECT 21.84 2.575 22.01 2.945 ;
      RECT 21.36 2.575 22.01 2.845 ;
      RECT 21.28 2.575 22.09 2.745 ;
      RECT 20.64 1.815 20.81 2.105 ;
      RECT 20.64 1.815 21.88 1.985 ;
      RECT 21.36 2.155 21.53 2.365 ;
      RECT 21 2.155 21.53 2.325 ;
      RECT 20.4 3.225 20.89 3.395 ;
      RECT 20.4 3.055 20.57 3.395 ;
      RECT 19.68 3.225 19.85 3.785 ;
      RECT 19.57 3.225 19.9 3.395 ;
      RECT 19.64 1.835 19.81 2.105 ;
      RECT 19.68 1.755 19.85 2.085 ;
      RECT 19.545 1.835 19.85 2.055 ;
      RECT 18.12 3.225 18.41 3.785 ;
      RECT 18.24 3.145 18.41 3.785 ;
      RECT 17.88 2.575 18.25 2.745 ;
      RECT 17.88 1.935 18.05 2.745 ;
      RECT 17.76 1.935 18.05 2.105 ;
      RECT 14.35 1.74 14.52 2.935 ;
      RECT 14.35 1.74 14.815 1.91 ;
      RECT 14.35 6.97 14.815 7.14 ;
      RECT 14.35 5.945 14.52 7.14 ;
      RECT 13.36 1.74 13.53 2.935 ;
      RECT 13.36 1.74 13.825 1.91 ;
      RECT 13.36 6.97 13.825 7.14 ;
      RECT 13.36 5.945 13.53 7.14 ;
      RECT 11.505 2.635 11.675 3.865 ;
      RECT 11.56 0.855 11.73 2.805 ;
      RECT 11.505 0.575 11.675 1.025 ;
      RECT 11.505 7.855 11.675 8.305 ;
      RECT 11.56 6.075 11.73 8.025 ;
      RECT 11.505 5.015 11.675 6.245 ;
      RECT 10.985 0.575 11.155 3.865 ;
      RECT 10.985 2.075 11.39 2.405 ;
      RECT 10.985 1.235 11.39 1.565 ;
      RECT 10.985 5.015 11.155 8.305 ;
      RECT 10.985 7.315 11.39 7.645 ;
      RECT 10.985 6.475 11.39 6.805 ;
      RECT 8.26 3.615 8.775 3.785 ;
      RECT 8.605 3.225 8.775 3.785 ;
      RECT 8.71 3.145 8.88 3.475 ;
      RECT 8.5 2.535 8.775 2.945 ;
      RECT 8.38 2.535 8.775 2.745 ;
      RECT 6.85 3.145 7.02 3.505 ;
      RECT 6.85 3.225 8.19 3.395 ;
      RECT 8.02 3.055 8.19 3.395 ;
      RECT 6.58 2.575 6.75 2.945 ;
      RECT 6.1 2.575 6.75 2.845 ;
      RECT 6.02 2.575 6.83 2.745 ;
      RECT 5.38 1.815 5.55 2.105 ;
      RECT 5.38 1.815 6.62 1.985 ;
      RECT 6.1 2.155 6.27 2.365 ;
      RECT 5.74 2.155 6.27 2.325 ;
      RECT 5.14 3.225 5.63 3.395 ;
      RECT 5.14 3.055 5.31 3.395 ;
      RECT 4.42 3.225 4.59 3.785 ;
      RECT 4.31 3.225 4.64 3.395 ;
      RECT 4.38 1.835 4.55 2.105 ;
      RECT 4.42 1.755 4.59 2.085 ;
      RECT 4.285 1.835 4.59 2.055 ;
      RECT 2.86 3.225 3.15 3.785 ;
      RECT 2.98 3.145 3.15 3.785 ;
      RECT 2.62 2.575 2.99 2.745 ;
      RECT 2.62 1.935 2.79 2.745 ;
      RECT 2.5 1.935 2.79 2.105 ;
      RECT 75.76 0.575 75.93 1.085 ;
      RECT 75.76 2.395 75.93 3.865 ;
      RECT 75.76 5.015 75.93 6.485 ;
      RECT 75.76 7.795 75.93 8.305 ;
      RECT 74.77 0.575 74.94 1.085 ;
      RECT 74.77 2.395 74.94 3.865 ;
      RECT 74.77 5.015 74.94 6.485 ;
      RECT 74.77 7.795 74.94 8.305 ;
      RECT 73.405 0.575 73.575 3.865 ;
      RECT 73.405 5.015 73.575 8.305 ;
      RECT 72.975 0.575 73.145 1.085 ;
      RECT 72.975 1.655 73.145 3.865 ;
      RECT 72.975 5.015 73.145 7.225 ;
      RECT 72.975 7.795 73.145 8.305 ;
      RECT 71.605 1.66 71.775 2.935 ;
      RECT 71.605 5.945 71.775 7.22 ;
      RECT 69.3 1.755 69.47 2.105 ;
      RECT 69.06 2.495 69.23 2.825 ;
      RECT 68.58 2.495 68.75 2.945 ;
      RECT 68.34 1.755 68.51 2.105 ;
      RECT 68.1 2.495 68.27 2.825 ;
      RECT 67.35 3.485 67.52 3.815 ;
      RECT 66.66 2.495 66.83 2.945 ;
      RECT 66.18 2.495 66.35 2.825 ;
      RECT 65.7 2.495 65.87 2.825 ;
      RECT 65.22 2.495 65.39 2.945 ;
      RECT 64.98 3.485 65.15 3.815 ;
      RECT 64.74 2.495 64.91 3.225 ;
      RECT 64.26 2.495 64.43 2.825 ;
      RECT 64.02 1.755 64.19 2.105 ;
      RECT 63.54 3.055 63.71 3.475 ;
      RECT 63.3 2.495 63.47 2.825 ;
      RECT 63.06 3.145 63.23 3.505 ;
      RECT 62.82 2.495 62.99 2.945 ;
      RECT 62.34 2.495 62.51 2.945 ;
      RECT 62.13 1.755 62.3 2.105 ;
      RECT 62.13 3.145 62.3 3.505 ;
      RECT 60.5 0.575 60.67 1.085 ;
      RECT 60.5 2.395 60.67 3.865 ;
      RECT 60.5 5.015 60.67 6.485 ;
      RECT 60.5 7.795 60.67 8.305 ;
      RECT 59.51 0.575 59.68 1.085 ;
      RECT 59.51 2.395 59.68 3.865 ;
      RECT 59.51 5.015 59.68 6.485 ;
      RECT 59.51 7.795 59.68 8.305 ;
      RECT 58.145 0.575 58.315 3.865 ;
      RECT 58.145 5.015 58.315 8.305 ;
      RECT 57.715 0.575 57.885 1.085 ;
      RECT 57.715 1.655 57.885 3.865 ;
      RECT 57.715 5.015 57.885 7.225 ;
      RECT 57.715 7.795 57.885 8.305 ;
      RECT 56.345 1.66 56.515 2.935 ;
      RECT 56.345 5.945 56.515 7.22 ;
      RECT 54.04 1.755 54.21 2.105 ;
      RECT 53.8 2.495 53.97 2.825 ;
      RECT 53.32 2.495 53.49 2.945 ;
      RECT 53.08 1.755 53.25 2.105 ;
      RECT 52.84 2.495 53.01 2.825 ;
      RECT 52.09 3.485 52.26 3.815 ;
      RECT 51.4 2.495 51.57 2.945 ;
      RECT 50.92 2.495 51.09 2.825 ;
      RECT 50.44 2.495 50.61 2.825 ;
      RECT 49.96 2.495 50.13 2.945 ;
      RECT 49.72 3.485 49.89 3.815 ;
      RECT 49.48 2.495 49.65 3.225 ;
      RECT 49 2.495 49.17 2.825 ;
      RECT 48.76 1.755 48.93 2.105 ;
      RECT 48.28 3.055 48.45 3.475 ;
      RECT 48.04 2.495 48.21 2.825 ;
      RECT 47.8 3.145 47.97 3.505 ;
      RECT 47.56 2.495 47.73 2.945 ;
      RECT 47.08 2.495 47.25 2.945 ;
      RECT 46.87 1.755 47.04 2.105 ;
      RECT 46.87 3.145 47.04 3.505 ;
      RECT 45.24 0.575 45.41 1.085 ;
      RECT 45.24 2.395 45.41 3.865 ;
      RECT 45.24 5.015 45.41 6.485 ;
      RECT 45.24 7.795 45.41 8.305 ;
      RECT 44.25 0.575 44.42 1.085 ;
      RECT 44.25 2.395 44.42 3.865 ;
      RECT 44.25 5.015 44.42 6.485 ;
      RECT 44.25 7.795 44.42 8.305 ;
      RECT 42.885 0.575 43.055 3.865 ;
      RECT 42.885 5.015 43.055 8.305 ;
      RECT 42.455 0.575 42.625 1.085 ;
      RECT 42.455 1.655 42.625 3.865 ;
      RECT 42.455 5.015 42.625 7.225 ;
      RECT 42.455 7.795 42.625 8.305 ;
      RECT 41.085 1.66 41.255 2.935 ;
      RECT 41.085 5.945 41.255 7.22 ;
      RECT 38.78 1.755 38.95 2.105 ;
      RECT 38.54 2.495 38.71 2.825 ;
      RECT 38.06 2.495 38.23 2.945 ;
      RECT 37.82 1.755 37.99 2.105 ;
      RECT 37.58 2.495 37.75 2.825 ;
      RECT 36.83 3.485 37 3.815 ;
      RECT 36.14 2.495 36.31 2.945 ;
      RECT 35.66 2.495 35.83 2.825 ;
      RECT 35.18 2.495 35.35 2.825 ;
      RECT 34.7 2.495 34.87 2.945 ;
      RECT 34.46 3.485 34.63 3.815 ;
      RECT 34.22 2.495 34.39 3.225 ;
      RECT 33.74 2.495 33.91 2.825 ;
      RECT 33.5 1.755 33.67 2.105 ;
      RECT 33.02 3.055 33.19 3.475 ;
      RECT 32.78 2.495 32.95 2.825 ;
      RECT 32.54 3.145 32.71 3.505 ;
      RECT 32.3 2.495 32.47 2.945 ;
      RECT 31.82 2.495 31.99 2.945 ;
      RECT 31.61 1.755 31.78 2.105 ;
      RECT 31.61 3.145 31.78 3.505 ;
      RECT 29.98 0.575 30.15 1.085 ;
      RECT 29.98 2.395 30.15 3.865 ;
      RECT 29.98 5.015 30.15 6.485 ;
      RECT 29.98 7.795 30.15 8.305 ;
      RECT 28.99 0.575 29.16 1.085 ;
      RECT 28.99 2.395 29.16 3.865 ;
      RECT 28.99 5.015 29.16 6.485 ;
      RECT 28.99 7.795 29.16 8.305 ;
      RECT 27.625 0.575 27.795 3.865 ;
      RECT 27.625 5.015 27.795 8.305 ;
      RECT 27.195 0.575 27.365 1.085 ;
      RECT 27.195 1.655 27.365 3.865 ;
      RECT 27.195 5.015 27.365 7.225 ;
      RECT 27.195 7.795 27.365 8.305 ;
      RECT 25.825 1.66 25.995 2.935 ;
      RECT 25.825 5.945 25.995 7.22 ;
      RECT 23.52 1.755 23.69 2.105 ;
      RECT 23.28 2.495 23.45 2.825 ;
      RECT 22.8 2.495 22.97 2.945 ;
      RECT 22.56 1.755 22.73 2.105 ;
      RECT 22.32 2.495 22.49 2.825 ;
      RECT 21.57 3.485 21.74 3.815 ;
      RECT 20.88 2.495 21.05 2.945 ;
      RECT 20.4 2.495 20.57 2.825 ;
      RECT 19.92 2.495 20.09 2.825 ;
      RECT 19.44 2.495 19.61 2.945 ;
      RECT 19.2 3.485 19.37 3.815 ;
      RECT 18.96 2.495 19.13 3.225 ;
      RECT 18.48 2.495 18.65 2.825 ;
      RECT 18.24 1.755 18.41 2.105 ;
      RECT 17.76 3.055 17.93 3.475 ;
      RECT 17.52 2.495 17.69 2.825 ;
      RECT 17.28 3.145 17.45 3.505 ;
      RECT 17.04 2.495 17.21 2.945 ;
      RECT 16.56 2.495 16.73 2.945 ;
      RECT 16.35 1.755 16.52 2.105 ;
      RECT 16.35 3.145 16.52 3.505 ;
      RECT 14.72 0.575 14.89 1.085 ;
      RECT 14.72 2.395 14.89 3.865 ;
      RECT 14.72 5.015 14.89 6.485 ;
      RECT 14.72 7.795 14.89 8.305 ;
      RECT 13.73 0.575 13.9 1.085 ;
      RECT 13.73 2.395 13.9 3.865 ;
      RECT 13.73 5.015 13.9 6.485 ;
      RECT 13.73 7.795 13.9 8.305 ;
      RECT 12.365 0.575 12.535 3.865 ;
      RECT 12.365 5.015 12.535 8.305 ;
      RECT 11.935 0.575 12.105 1.085 ;
      RECT 11.935 1.655 12.105 3.865 ;
      RECT 11.935 5.015 12.105 7.225 ;
      RECT 11.935 7.795 12.105 8.305 ;
      RECT 10.565 1.66 10.735 2.935 ;
      RECT 10.565 5.945 10.735 7.22 ;
      RECT 8.26 1.755 8.43 2.105 ;
      RECT 8.02 2.495 8.19 2.825 ;
      RECT 7.54 2.495 7.71 2.945 ;
      RECT 7.3 1.755 7.47 2.105 ;
      RECT 7.06 2.495 7.23 2.825 ;
      RECT 6.31 3.485 6.48 3.815 ;
      RECT 5.62 2.495 5.79 2.945 ;
      RECT 5.14 2.495 5.31 2.825 ;
      RECT 4.66 2.495 4.83 2.825 ;
      RECT 4.18 2.495 4.35 2.945 ;
      RECT 3.94 3.485 4.11 3.815 ;
      RECT 3.7 2.495 3.87 3.225 ;
      RECT 3.22 2.495 3.39 2.825 ;
      RECT 2.98 1.755 3.15 2.105 ;
      RECT 2.5 3.055 2.67 3.475 ;
      RECT 2.26 2.495 2.43 2.825 ;
      RECT 2.02 3.145 2.19 3.505 ;
      RECT 1.78 2.495 1.95 2.945 ;
      RECT 1.3 2.495 1.47 2.945 ;
      RECT 1.09 1.755 1.26 2.105 ;
      RECT 1.09 3.145 1.26 3.505 ;
  END
END sky130_osu_ring_oscillator_mpr2xa_8

MACRO sky130_osu_ring_oscillator_mpr2ya_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ya_8 0 0 ;
  SIZE 76.3 BY 8.88 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT 64.9 1.855 65.23 2.585 ;
      RECT 64.93 1.04 65.24 1.985 ;
      RECT 64.905 1.04 65.28 1.41 ;
      RECT 49.64 1.855 49.97 2.585 ;
      RECT 49.67 1.04 49.98 1.985 ;
      RECT 49.645 1.04 50.02 1.41 ;
      RECT 34.38 1.855 34.71 2.585 ;
      RECT 34.41 1.04 34.72 1.985 ;
      RECT 34.385 1.04 34.76 1.41 ;
      RECT 19.12 1.855 19.45 2.585 ;
      RECT 19.15 1.04 19.46 1.985 ;
      RECT 19.125 1.04 19.5 1.41 ;
      RECT 3.86 1.855 4.19 2.585 ;
      RECT 3.89 1.04 4.2 1.985 ;
      RECT 3.865 1.04 4.24 1.41 ;
      RECT 69.34 2.015 69.67 2.745 ;
      RECT 68.14 2.88 68.47 3.61 ;
      RECT 67.3 1.855 68.03 2.185 ;
      RECT 65.86 1.855 66.59 2.185 ;
      RECT 66.22 2.76 66.55 3.49 ;
      RECT 63.7 2.015 64.03 2.745 ;
      RECT 62.98 2.015 63.31 2.745 ;
      RECT 54.08 2.015 54.41 2.745 ;
      RECT 52.88 2.88 53.21 3.61 ;
      RECT 52.04 1.855 52.77 2.185 ;
      RECT 50.6 1.855 51.33 2.185 ;
      RECT 50.96 2.76 51.29 3.49 ;
      RECT 48.44 2.015 48.77 2.745 ;
      RECT 47.72 2.015 48.05 2.745 ;
      RECT 38.82 2.015 39.15 2.745 ;
      RECT 37.62 2.88 37.95 3.61 ;
      RECT 36.78 1.855 37.51 2.185 ;
      RECT 35.34 1.855 36.07 2.185 ;
      RECT 35.7 2.76 36.03 3.49 ;
      RECT 33.18 2.015 33.51 2.745 ;
      RECT 32.46 2.015 32.79 2.745 ;
      RECT 23.56 2.015 23.89 2.745 ;
      RECT 22.36 2.88 22.69 3.61 ;
      RECT 21.52 1.855 22.25 2.185 ;
      RECT 20.08 1.855 20.81 2.185 ;
      RECT 20.44 2.76 20.77 3.49 ;
      RECT 17.92 2.015 18.25 2.745 ;
      RECT 17.2 2.015 17.53 2.745 ;
      RECT 8.3 2.015 8.63 2.745 ;
      RECT 7.1 2.88 7.43 3.61 ;
      RECT 6.26 1.855 6.99 2.185 ;
      RECT 4.82 1.855 5.55 2.185 ;
      RECT 5.18 2.76 5.51 3.49 ;
      RECT 2.66 2.015 2.99 2.745 ;
      RECT 1.94 2.015 2.27 2.745 ;
    LAYER via2 ;
      RECT 69.405 2.48 69.605 2.68 ;
      RECT 68.205 3.04 68.405 3.24 ;
      RECT 67.365 1.92 67.565 2.12 ;
      RECT 66.285 2.825 66.485 3.025 ;
      RECT 65.925 1.92 66.125 2.12 ;
      RECT 64.995 1.125 65.195 1.325 ;
      RECT 64.965 1.92 65.165 2.12 ;
      RECT 63.765 2.48 63.965 2.68 ;
      RECT 63.045 2.48 63.245 2.68 ;
      RECT 54.145 2.48 54.345 2.68 ;
      RECT 52.945 3.04 53.145 3.24 ;
      RECT 52.105 1.92 52.305 2.12 ;
      RECT 51.025 2.825 51.225 3.025 ;
      RECT 50.665 1.92 50.865 2.12 ;
      RECT 49.735 1.125 49.935 1.325 ;
      RECT 49.705 1.92 49.905 2.12 ;
      RECT 48.505 2.48 48.705 2.68 ;
      RECT 47.785 2.48 47.985 2.68 ;
      RECT 38.885 2.48 39.085 2.68 ;
      RECT 37.685 3.04 37.885 3.24 ;
      RECT 36.845 1.92 37.045 2.12 ;
      RECT 35.765 2.825 35.965 3.025 ;
      RECT 35.405 1.92 35.605 2.12 ;
      RECT 34.475 1.125 34.675 1.325 ;
      RECT 34.445 1.92 34.645 2.12 ;
      RECT 33.245 2.48 33.445 2.68 ;
      RECT 32.525 2.48 32.725 2.68 ;
      RECT 23.625 2.48 23.825 2.68 ;
      RECT 22.425 3.04 22.625 3.24 ;
      RECT 21.585 1.92 21.785 2.12 ;
      RECT 20.505 2.825 20.705 3.025 ;
      RECT 20.145 1.92 20.345 2.12 ;
      RECT 19.215 1.125 19.415 1.325 ;
      RECT 19.185 1.92 19.385 2.12 ;
      RECT 17.985 2.48 18.185 2.68 ;
      RECT 17.265 2.48 17.465 2.68 ;
      RECT 8.365 2.48 8.565 2.68 ;
      RECT 7.165 3.04 7.365 3.24 ;
      RECT 6.325 1.92 6.525 2.12 ;
      RECT 5.245 2.825 5.445 3.025 ;
      RECT 4.885 1.92 5.085 2.12 ;
      RECT 3.955 1.125 4.155 1.325 ;
      RECT 3.925 1.92 4.125 2.12 ;
      RECT 2.725 2.48 2.925 2.68 ;
      RECT 2.005 2.48 2.205 2.68 ;
    LAYER met2 ;
      RECT 11.53 6.28 11.85 6.605 ;
      RECT 11.56 5.695 11.73 6.605 ;
      RECT 11.56 5.695 11.735 6.045 ;
      RECT 11.56 5.695 12.535 5.87 ;
      RECT 12.36 1.965 12.535 5.87 ;
      RECT 2.685 2.44 2.965 2.72 ;
      RECT 2.685 2.44 2.985 2.615 ;
      RECT 2.775 2.33 3.035 2.59 ;
      RECT 2.74 2.425 3.035 2.59 ;
      RECT 2.875 0.73 3.03 2.59 ;
      RECT 12.305 1.965 12.655 2.315 ;
      RECT 9.895 2.025 12.655 2.195 ;
      RECT 9.895 0.73 10.065 2.195 ;
      RECT 9.9 0.195 10.065 2.195 ;
      RECT 75.73 1.095 76.07 1.445 ;
      RECT 75.765 0.195 75.93 1.445 ;
      RECT 2.875 0.73 10.065 0.9 ;
      RECT 9.9 0.195 75.93 0.36 ;
      RECT 72.57 6.28 72.89 6.605 ;
      RECT 72.6 5.695 72.77 6.605 ;
      RECT 72.6 5.695 72.775 6.045 ;
      RECT 72.6 5.695 73.575 5.87 ;
      RECT 73.4 1.965 73.575 5.87 ;
      RECT 63.725 2.44 64.005 2.72 ;
      RECT 63.725 2.44 64.025 2.615 ;
      RECT 63.815 2.33 64.075 2.59 ;
      RECT 63.78 2.425 64.075 2.59 ;
      RECT 63.915 0.73 64.07 2.59 ;
      RECT 73.345 1.965 73.695 2.315 ;
      RECT 70.935 2.025 73.695 2.195 ;
      RECT 70.935 0.73 71.105 2.195 ;
      RECT 60.47 1.095 60.81 1.445 ;
      RECT 60.47 1.26 64.07 1.435 ;
      RECT 63.915 0.73 71.105 0.9 ;
      RECT 73.37 6.655 73.695 6.98 ;
      RECT 72.255 6.745 73.695 6.915 ;
      RECT 72.255 2.395 72.415 6.915 ;
      RECT 72.57 2.365 72.89 2.685 ;
      RECT 72.255 2.395 72.89 2.565 ;
      RECT 71.52 5.86 71.86 6.21 ;
      RECT 71.6 2.705 71.775 6.21 ;
      RECT 71.525 2.705 71.865 3.055 ;
      RECT 70.965 2.705 71.305 3.055 ;
      RECT 70.265 2.77 71.305 2.97 ;
      RECT 70.265 2.765 70.575 2.97 ;
      RECT 70.265 1.04 70.47 2.97 ;
      RECT 71.055 2.7 71.225 3.055 ;
      RECT 64.905 1.04 65.28 1.41 ;
      RECT 64.905 1.04 70.47 1.245 ;
      RECT 69.365 2.44 69.645 2.72 ;
      RECT 69.36 2.44 69.645 2.673 ;
      RECT 69.34 2.44 69.645 2.65 ;
      RECT 69.33 2.44 69.645 2.63 ;
      RECT 69.32 2.44 69.645 2.615 ;
      RECT 69.295 2.44 69.645 2.588 ;
      RECT 69.285 2.44 69.645 2.563 ;
      RECT 69.24 2.295 69.52 2.555 ;
      RECT 69.24 2.39 69.62 2.555 ;
      RECT 69.24 2.335 69.565 2.555 ;
      RECT 69.24 2.327 69.56 2.555 ;
      RECT 69.24 2.317 69.555 2.555 ;
      RECT 69.24 2.305 69.55 2.555 ;
      RECT 68.165 3 68.445 3.28 ;
      RECT 68.165 3 68.48 3.26 ;
      RECT 68.2 2.42 68.25 2.68 ;
      RECT 67.99 2.42 67.995 2.68 ;
      RECT 67.185 1.975 67.215 2.235 ;
      RECT 66.955 1.975 67.03 2.235 ;
      RECT 68.175 2.37 68.2 2.68 ;
      RECT 68.17 2.327 68.175 2.68 ;
      RECT 68.165 2.31 68.17 2.68 ;
      RECT 68.16 2.297 68.165 2.68 ;
      RECT 68.085 2.18 68.16 2.68 ;
      RECT 68.04 1.997 68.085 2.68 ;
      RECT 68.035 1.925 68.04 2.68 ;
      RECT 68.02 1.9 68.035 2.68 ;
      RECT 67.995 1.862 68.02 2.68 ;
      RECT 67.985 1.842 67.995 2.402 ;
      RECT 67.97 1.834 67.985 2.357 ;
      RECT 67.965 1.826 67.97 2.328 ;
      RECT 67.96 1.823 67.965 2.308 ;
      RECT 67.955 1.82 67.96 2.288 ;
      RECT 67.95 1.817 67.955 2.268 ;
      RECT 67.92 1.806 67.95 2.205 ;
      RECT 67.9 1.791 67.92 2.12 ;
      RECT 67.895 1.783 67.9 2.083 ;
      RECT 67.885 1.777 67.895 2.05 ;
      RECT 67.87 1.769 67.885 2.01 ;
      RECT 67.865 1.762 67.87 1.97 ;
      RECT 67.86 1.759 67.865 1.948 ;
      RECT 67.855 1.756 67.86 1.935 ;
      RECT 67.85 1.755 67.855 1.925 ;
      RECT 67.835 1.749 67.85 1.915 ;
      RECT 67.81 1.736 67.835 1.9 ;
      RECT 67.76 1.711 67.81 1.871 ;
      RECT 67.745 1.69 67.76 1.846 ;
      RECT 67.735 1.683 67.745 1.835 ;
      RECT 67.68 1.664 67.735 1.808 ;
      RECT 67.655 1.642 67.68 1.781 ;
      RECT 67.65 1.635 67.655 1.776 ;
      RECT 67.635 1.635 67.65 1.774 ;
      RECT 67.61 1.627 67.635 1.77 ;
      RECT 67.595 1.625 67.61 1.766 ;
      RECT 67.565 1.625 67.595 1.763 ;
      RECT 67.555 1.625 67.565 1.758 ;
      RECT 67.51 1.625 67.555 1.756 ;
      RECT 67.481 1.625 67.51 1.757 ;
      RECT 67.395 1.625 67.481 1.759 ;
      RECT 67.381 1.626 67.395 1.761 ;
      RECT 67.295 1.627 67.381 1.763 ;
      RECT 67.28 1.628 67.295 1.773 ;
      RECT 67.275 1.629 67.28 1.782 ;
      RECT 67.255 1.632 67.275 1.792 ;
      RECT 67.24 1.64 67.255 1.807 ;
      RECT 67.22 1.658 67.24 1.822 ;
      RECT 67.21 1.67 67.22 1.845 ;
      RECT 67.2 1.679 67.21 1.875 ;
      RECT 67.185 1.691 67.2 1.92 ;
      RECT 67.13 1.724 67.185 2.235 ;
      RECT 67.125 1.752 67.13 2.235 ;
      RECT 67.105 1.767 67.125 2.235 ;
      RECT 67.07 1.827 67.105 2.235 ;
      RECT 67.068 1.877 67.07 2.235 ;
      RECT 67.065 1.885 67.068 2.235 ;
      RECT 67.055 1.9 67.065 2.235 ;
      RECT 67.05 1.912 67.055 2.235 ;
      RECT 67.04 1.937 67.05 2.235 ;
      RECT 67.03 1.965 67.04 2.235 ;
      RECT 64.935 3.47 64.985 3.73 ;
      RECT 67.845 3.02 67.905 3.28 ;
      RECT 67.83 3.02 67.845 3.29 ;
      RECT 67.811 3.02 67.83 3.323 ;
      RECT 67.725 3.02 67.811 3.448 ;
      RECT 67.645 3.02 67.725 3.63 ;
      RECT 67.64 3.257 67.645 3.715 ;
      RECT 67.615 3.327 67.64 3.743 ;
      RECT 67.61 3.397 67.615 3.77 ;
      RECT 67.59 3.469 67.61 3.792 ;
      RECT 67.585 3.536 67.59 3.815 ;
      RECT 67.575 3.565 67.585 3.83 ;
      RECT 67.565 3.587 67.575 3.847 ;
      RECT 67.56 3.597 67.565 3.858 ;
      RECT 67.555 3.605 67.56 3.866 ;
      RECT 67.545 3.613 67.555 3.878 ;
      RECT 67.54 3.625 67.545 3.888 ;
      RECT 67.535 3.633 67.54 3.893 ;
      RECT 67.515 3.651 67.535 3.903 ;
      RECT 67.51 3.668 67.515 3.91 ;
      RECT 67.505 3.676 67.51 3.911 ;
      RECT 67.5 3.687 67.505 3.913 ;
      RECT 67.46 3.725 67.5 3.923 ;
      RECT 67.455 3.76 67.46 3.934 ;
      RECT 67.45 3.765 67.455 3.937 ;
      RECT 67.425 3.775 67.45 3.944 ;
      RECT 67.415 3.789 67.425 3.953 ;
      RECT 67.395 3.801 67.415 3.956 ;
      RECT 67.345 3.82 67.395 3.96 ;
      RECT 67.3 3.835 67.345 3.965 ;
      RECT 67.235 3.838 67.3 3.971 ;
      RECT 67.22 3.836 67.235 3.978 ;
      RECT 67.19 3.835 67.22 3.978 ;
      RECT 67.151 3.834 67.19 3.974 ;
      RECT 67.065 3.831 67.151 3.97 ;
      RECT 67.048 3.829 67.065 3.967 ;
      RECT 66.962 3.827 67.048 3.964 ;
      RECT 66.876 3.824 66.962 3.958 ;
      RECT 66.79 3.82 66.876 3.953 ;
      RECT 66.712 3.817 66.79 3.949 ;
      RECT 66.626 3.814 66.712 3.947 ;
      RECT 66.54 3.811 66.626 3.944 ;
      RECT 66.482 3.809 66.54 3.941 ;
      RECT 66.396 3.806 66.482 3.939 ;
      RECT 66.31 3.802 66.396 3.937 ;
      RECT 66.224 3.799 66.31 3.934 ;
      RECT 66.138 3.795 66.224 3.932 ;
      RECT 66.052 3.791 66.138 3.929 ;
      RECT 65.966 3.788 66.052 3.927 ;
      RECT 65.88 3.784 65.966 3.924 ;
      RECT 65.794 3.781 65.88 3.922 ;
      RECT 65.708 3.777 65.794 3.919 ;
      RECT 65.622 3.774 65.708 3.917 ;
      RECT 65.536 3.77 65.622 3.914 ;
      RECT 65.45 3.767 65.536 3.912 ;
      RECT 65.44 3.765 65.45 3.908 ;
      RECT 65.435 3.765 65.44 3.906 ;
      RECT 65.395 3.76 65.435 3.9 ;
      RECT 65.381 3.751 65.395 3.893 ;
      RECT 65.295 3.721 65.381 3.878 ;
      RECT 65.275 3.687 65.295 3.863 ;
      RECT 65.205 3.656 65.275 3.85 ;
      RECT 65.2 3.631 65.205 3.839 ;
      RECT 65.195 3.625 65.2 3.837 ;
      RECT 65.126 3.47 65.195 3.825 ;
      RECT 65.04 3.47 65.126 3.799 ;
      RECT 65.015 3.47 65.04 3.778 ;
      RECT 65.01 3.47 65.015 3.768 ;
      RECT 65.005 3.47 65.01 3.76 ;
      RECT 64.985 3.47 65.005 3.743 ;
      RECT 67.405 2.04 67.665 2.3 ;
      RECT 67.39 2.04 67.665 2.203 ;
      RECT 67.36 2.04 67.665 2.178 ;
      RECT 67.325 1.88 67.605 2.16 ;
      RECT 67.295 3.37 67.355 3.63 ;
      RECT 66.32 2.06 66.375 2.32 ;
      RECT 67.255 3.327 67.295 3.63 ;
      RECT 67.226 3.248 67.255 3.63 ;
      RECT 67.14 3.12 67.226 3.63 ;
      RECT 67.12 3 67.14 3.63 ;
      RECT 67.095 2.951 67.12 3.63 ;
      RECT 67.09 2.916 67.095 3.48 ;
      RECT 67.06 2.876 67.09 3.418 ;
      RECT 67.035 2.813 67.06 3.333 ;
      RECT 67.025 2.775 67.035 3.27 ;
      RECT 67.01 2.75 67.025 3.231 ;
      RECT 66.967 2.708 67.01 3.137 ;
      RECT 66.965 2.681 66.967 3.064 ;
      RECT 66.96 2.676 66.965 3.055 ;
      RECT 66.955 2.669 66.96 3.03 ;
      RECT 66.95 2.663 66.955 3.015 ;
      RECT 66.945 2.657 66.95 3.003 ;
      RECT 66.935 2.648 66.945 2.985 ;
      RECT 66.93 2.639 66.935 2.963 ;
      RECT 66.905 2.62 66.93 2.913 ;
      RECT 66.9 2.601 66.905 2.863 ;
      RECT 66.885 2.587 66.9 2.823 ;
      RECT 66.88 2.573 66.885 2.79 ;
      RECT 66.875 2.566 66.88 2.783 ;
      RECT 66.86 2.553 66.875 2.775 ;
      RECT 66.815 2.515 66.86 2.748 ;
      RECT 66.785 2.468 66.815 2.713 ;
      RECT 66.765 2.437 66.785 2.69 ;
      RECT 66.685 2.37 66.765 2.643 ;
      RECT 66.655 2.3 66.685 2.59 ;
      RECT 66.65 2.277 66.655 2.573 ;
      RECT 66.62 2.255 66.65 2.558 ;
      RECT 66.59 2.214 66.62 2.53 ;
      RECT 66.585 2.189 66.59 2.515 ;
      RECT 66.58 2.183 66.585 2.508 ;
      RECT 66.57 2.06 66.58 2.5 ;
      RECT 66.56 2.06 66.57 2.493 ;
      RECT 66.555 2.06 66.56 2.485 ;
      RECT 66.535 2.06 66.555 2.473 ;
      RECT 66.485 2.06 66.535 2.443 ;
      RECT 66.43 2.06 66.485 2.393 ;
      RECT 66.4 2.06 66.43 2.353 ;
      RECT 66.375 2.06 66.4 2.33 ;
      RECT 66.245 2.785 66.525 3.065 ;
      RECT 66.21 2.7 66.47 2.96 ;
      RECT 66.21 2.782 66.48 2.96 ;
      RECT 64.41 2.155 64.415 2.64 ;
      RECT 64.3 2.34 64.305 2.64 ;
      RECT 64.21 2.38 64.275 2.64 ;
      RECT 65.885 1.88 65.975 2.51 ;
      RECT 65.85 1.93 65.855 2.51 ;
      RECT 65.795 1.955 65.805 2.51 ;
      RECT 65.75 1.955 65.76 2.51 ;
      RECT 66.12 1.88 66.165 2.16 ;
      RECT 64.97 1.61 65.17 1.75 ;
      RECT 66.086 1.88 66.12 2.172 ;
      RECT 66 1.88 66.086 2.212 ;
      RECT 65.985 1.88 66 2.253 ;
      RECT 65.98 1.88 65.985 2.273 ;
      RECT 65.975 1.88 65.98 2.293 ;
      RECT 65.855 1.922 65.885 2.51 ;
      RECT 65.805 1.942 65.85 2.51 ;
      RECT 65.79 1.957 65.795 2.51 ;
      RECT 65.76 1.957 65.79 2.51 ;
      RECT 65.715 1.942 65.75 2.51 ;
      RECT 65.71 1.93 65.715 2.29 ;
      RECT 65.705 1.927 65.71 2.27 ;
      RECT 65.69 1.917 65.705 2.223 ;
      RECT 65.685 1.91 65.69 2.186 ;
      RECT 65.68 1.907 65.685 2.169 ;
      RECT 65.665 1.897 65.68 2.125 ;
      RECT 65.66 1.888 65.665 2.085 ;
      RECT 65.655 1.884 65.66 2.07 ;
      RECT 65.645 1.878 65.655 2.053 ;
      RECT 65.605 1.859 65.645 2.028 ;
      RECT 65.6 1.841 65.605 2.008 ;
      RECT 65.59 1.835 65.6 2.003 ;
      RECT 65.56 1.819 65.59 1.99 ;
      RECT 65.545 1.801 65.56 1.973 ;
      RECT 65.53 1.789 65.545 1.96 ;
      RECT 65.525 1.781 65.53 1.953 ;
      RECT 65.495 1.767 65.525 1.94 ;
      RECT 65.49 1.752 65.495 1.928 ;
      RECT 65.48 1.746 65.49 1.92 ;
      RECT 65.46 1.734 65.48 1.908 ;
      RECT 65.45 1.722 65.46 1.895 ;
      RECT 65.42 1.706 65.45 1.88 ;
      RECT 65.4 1.686 65.42 1.863 ;
      RECT 65.395 1.676 65.4 1.853 ;
      RECT 65.37 1.664 65.395 1.84 ;
      RECT 65.365 1.652 65.37 1.828 ;
      RECT 65.36 1.647 65.365 1.824 ;
      RECT 65.345 1.64 65.36 1.816 ;
      RECT 65.335 1.627 65.345 1.806 ;
      RECT 65.33 1.625 65.335 1.8 ;
      RECT 65.305 1.618 65.33 1.789 ;
      RECT 65.3 1.611 65.305 1.778 ;
      RECT 65.275 1.61 65.3 1.765 ;
      RECT 65.256 1.61 65.275 1.755 ;
      RECT 65.17 1.61 65.256 1.752 ;
      RECT 64.94 1.61 64.97 1.755 ;
      RECT 64.9 1.617 64.94 1.768 ;
      RECT 64.875 1.627 64.9 1.781 ;
      RECT 64.86 1.636 64.875 1.791 ;
      RECT 64.83 1.641 64.86 1.81 ;
      RECT 64.825 1.647 64.83 1.828 ;
      RECT 64.805 1.657 64.825 1.843 ;
      RECT 64.795 1.67 64.805 1.863 ;
      RECT 64.78 1.682 64.795 1.88 ;
      RECT 64.775 1.692 64.78 1.89 ;
      RECT 64.77 1.697 64.775 1.895 ;
      RECT 64.76 1.705 64.77 1.908 ;
      RECT 64.71 1.737 64.76 1.945 ;
      RECT 64.695 1.772 64.71 1.986 ;
      RECT 64.69 1.782 64.695 2.001 ;
      RECT 64.685 1.787 64.69 2.008 ;
      RECT 64.66 1.803 64.685 2.028 ;
      RECT 64.645 1.824 64.66 2.053 ;
      RECT 64.62 1.845 64.645 2.078 ;
      RECT 64.61 1.864 64.62 2.101 ;
      RECT 64.585 1.882 64.61 2.124 ;
      RECT 64.57 1.902 64.585 2.148 ;
      RECT 64.565 1.912 64.57 2.16 ;
      RECT 64.55 1.924 64.565 2.18 ;
      RECT 64.54 1.939 64.55 2.22 ;
      RECT 64.535 1.947 64.54 2.248 ;
      RECT 64.525 1.957 64.535 2.268 ;
      RECT 64.52 1.97 64.525 2.293 ;
      RECT 64.515 1.983 64.52 2.313 ;
      RECT 64.51 1.989 64.515 2.335 ;
      RECT 64.5 1.998 64.51 2.355 ;
      RECT 64.495 2.018 64.5 2.378 ;
      RECT 64.49 2.024 64.495 2.398 ;
      RECT 64.485 2.031 64.49 2.42 ;
      RECT 64.48 2.042 64.485 2.433 ;
      RECT 64.47 2.052 64.48 2.458 ;
      RECT 64.45 2.077 64.47 2.64 ;
      RECT 64.42 2.117 64.45 2.64 ;
      RECT 64.415 2.147 64.42 2.64 ;
      RECT 64.39 2.175 64.41 2.64 ;
      RECT 64.36 2.22 64.39 2.64 ;
      RECT 64.355 2.247 64.36 2.64 ;
      RECT 64.335 2.265 64.355 2.64 ;
      RECT 64.325 2.29 64.335 2.64 ;
      RECT 64.32 2.302 64.325 2.64 ;
      RECT 64.305 2.325 64.32 2.64 ;
      RECT 64.285 2.352 64.3 2.64 ;
      RECT 64.275 2.375 64.285 2.64 ;
      RECT 66.065 3.26 66.145 3.52 ;
      RECT 65.3 2.48 65.37 2.74 ;
      RECT 66.031 3.227 66.065 3.52 ;
      RECT 65.945 3.13 66.031 3.52 ;
      RECT 65.925 3.042 65.945 3.52 ;
      RECT 65.915 3.012 65.925 3.52 ;
      RECT 65.905 2.992 65.915 3.52 ;
      RECT 65.885 2.979 65.905 3.52 ;
      RECT 65.87 2.969 65.885 3.348 ;
      RECT 65.865 2.962 65.87 3.303 ;
      RECT 65.855 2.956 65.865 3.293 ;
      RECT 65.845 2.948 65.855 3.275 ;
      RECT 65.84 2.942 65.845 3.263 ;
      RECT 65.83 2.937 65.84 3.25 ;
      RECT 65.81 2.927 65.83 3.223 ;
      RECT 65.77 2.906 65.81 3.175 ;
      RECT 65.755 2.887 65.77 3.133 ;
      RECT 65.73 2.873 65.755 3.103 ;
      RECT 65.72 2.861 65.73 3.07 ;
      RECT 65.715 2.856 65.72 3.06 ;
      RECT 65.685 2.842 65.715 3.04 ;
      RECT 65.675 2.826 65.685 3.013 ;
      RECT 65.67 2.821 65.675 3.003 ;
      RECT 65.645 2.812 65.67 2.983 ;
      RECT 65.635 2.8 65.645 2.963 ;
      RECT 65.565 2.768 65.635 2.938 ;
      RECT 65.56 2.737 65.565 2.915 ;
      RECT 65.511 2.48 65.56 2.898 ;
      RECT 65.425 2.48 65.511 2.857 ;
      RECT 65.37 2.48 65.425 2.785 ;
      RECT 65.46 3.265 65.62 3.525 ;
      RECT 64.985 1.88 65.035 2.565 ;
      RECT 64.775 2.305 64.81 2.565 ;
      RECT 65.09 1.88 65.095 2.34 ;
      RECT 65.18 1.88 65.205 2.16 ;
      RECT 65.455 3.262 65.46 3.525 ;
      RECT 65.42 3.25 65.455 3.525 ;
      RECT 65.36 3.223 65.42 3.525 ;
      RECT 65.355 3.206 65.36 3.379 ;
      RECT 65.35 3.203 65.355 3.366 ;
      RECT 65.33 3.196 65.35 3.353 ;
      RECT 65.295 3.179 65.33 3.335 ;
      RECT 65.255 3.158 65.295 3.315 ;
      RECT 65.25 3.146 65.255 3.303 ;
      RECT 65.21 3.132 65.25 3.289 ;
      RECT 65.19 3.115 65.21 3.271 ;
      RECT 65.18 3.107 65.19 3.263 ;
      RECT 65.165 1.88 65.18 2.178 ;
      RECT 65.15 3.097 65.18 3.25 ;
      RECT 65.135 1.88 65.165 2.223 ;
      RECT 65.14 3.087 65.15 3.237 ;
      RECT 65.11 3.072 65.14 3.224 ;
      RECT 65.095 1.88 65.135 2.29 ;
      RECT 65.095 3.04 65.11 3.21 ;
      RECT 65.09 3.012 65.095 3.204 ;
      RECT 65.085 1.88 65.09 2.345 ;
      RECT 65.075 2.982 65.09 3.198 ;
      RECT 65.08 1.88 65.085 2.358 ;
      RECT 65.07 1.88 65.08 2.378 ;
      RECT 65.035 2.895 65.075 3.183 ;
      RECT 65.035 1.88 65.07 2.418 ;
      RECT 65.03 2.827 65.035 3.171 ;
      RECT 65.015 2.782 65.03 3.166 ;
      RECT 65.01 2.72 65.015 3.161 ;
      RECT 64.985 2.627 65.01 3.154 ;
      RECT 64.98 1.88 64.985 3.146 ;
      RECT 64.965 1.88 64.98 3.133 ;
      RECT 64.945 1.88 64.965 3.09 ;
      RECT 64.935 1.88 64.945 3.04 ;
      RECT 64.93 1.88 64.935 3.013 ;
      RECT 64.925 1.88 64.93 2.991 ;
      RECT 64.92 2.106 64.925 2.974 ;
      RECT 64.915 2.128 64.92 2.952 ;
      RECT 64.91 2.17 64.915 2.935 ;
      RECT 64.88 2.22 64.91 2.879 ;
      RECT 64.875 2.247 64.88 2.821 ;
      RECT 64.86 2.265 64.875 2.785 ;
      RECT 64.855 2.283 64.86 2.749 ;
      RECT 64.849 2.29 64.855 2.73 ;
      RECT 64.845 2.297 64.849 2.713 ;
      RECT 64.84 2.302 64.845 2.682 ;
      RECT 64.83 2.305 64.84 2.657 ;
      RECT 64.82 2.305 64.83 2.623 ;
      RECT 64.815 2.305 64.82 2.6 ;
      RECT 64.81 2.305 64.815 2.58 ;
      RECT 63.43 3.47 63.69 3.73 ;
      RECT 63.45 3.397 63.63 3.73 ;
      RECT 63.45 3.14 63.625 3.73 ;
      RECT 63.45 2.932 63.615 3.73 ;
      RECT 63.455 2.85 63.615 3.73 ;
      RECT 63.455 2.615 63.605 3.73 ;
      RECT 63.455 2.462 63.6 3.73 ;
      RECT 63.46 2.447 63.6 3.73 ;
      RECT 63.51 2.162 63.6 3.73 ;
      RECT 63.465 2.397 63.6 3.73 ;
      RECT 63.495 2.215 63.6 3.73 ;
      RECT 63.48 2.327 63.6 3.73 ;
      RECT 63.485 2.285 63.6 3.73 ;
      RECT 63.48 2.327 63.615 2.39 ;
      RECT 63.515 1.915 63.62 2.335 ;
      RECT 63.515 1.915 63.635 2.318 ;
      RECT 63.515 1.915 63.67 2.28 ;
      RECT 63.51 2.162 63.72 2.213 ;
      RECT 63.515 1.915 63.775 2.175 ;
      RECT 62.775 2.62 63.035 2.88 ;
      RECT 62.775 2.62 63.045 2.838 ;
      RECT 62.775 2.62 63.131 2.809 ;
      RECT 62.775 2.62 63.2 2.761 ;
      RECT 62.775 2.62 63.235 2.73 ;
      RECT 63.005 2.44 63.285 2.72 ;
      RECT 62.84 2.605 63.285 2.72 ;
      RECT 62.93 2.482 63.035 2.88 ;
      RECT 62.86 2.545 63.285 2.72 ;
      RECT 57.31 6.28 57.63 6.605 ;
      RECT 57.34 5.695 57.51 6.605 ;
      RECT 57.34 5.695 57.515 6.045 ;
      RECT 57.34 5.695 58.315 5.87 ;
      RECT 58.14 1.965 58.315 5.87 ;
      RECT 48.465 2.44 48.745 2.72 ;
      RECT 48.465 2.44 48.765 2.615 ;
      RECT 48.555 2.33 48.815 2.59 ;
      RECT 48.52 2.425 48.815 2.59 ;
      RECT 48.655 0.73 48.81 2.59 ;
      RECT 58.085 1.965 58.435 2.315 ;
      RECT 55.675 2.025 58.435 2.195 ;
      RECT 55.675 0.73 55.845 2.195 ;
      RECT 45.21 1.095 45.55 1.445 ;
      RECT 45.21 1.26 48.81 1.435 ;
      RECT 48.655 0.73 55.845 0.9 ;
      RECT 58.11 6.655 58.435 6.98 ;
      RECT 56.995 6.745 58.435 6.915 ;
      RECT 56.995 2.395 57.155 6.915 ;
      RECT 57.31 2.365 57.63 2.685 ;
      RECT 56.995 2.395 57.63 2.565 ;
      RECT 56.26 5.86 56.6 6.21 ;
      RECT 56.34 2.705 56.515 6.21 ;
      RECT 56.265 2.705 56.605 3.055 ;
      RECT 55.705 2.705 56.045 3.055 ;
      RECT 55.005 2.77 56.045 2.97 ;
      RECT 55.005 2.765 55.315 2.97 ;
      RECT 55.005 1.04 55.21 2.97 ;
      RECT 55.795 2.7 55.965 3.055 ;
      RECT 49.645 1.04 50.02 1.41 ;
      RECT 49.645 1.04 55.21 1.245 ;
      RECT 54.105 2.44 54.385 2.72 ;
      RECT 54.1 2.44 54.385 2.673 ;
      RECT 54.08 2.44 54.385 2.65 ;
      RECT 54.07 2.44 54.385 2.63 ;
      RECT 54.06 2.44 54.385 2.615 ;
      RECT 54.035 2.44 54.385 2.588 ;
      RECT 54.025 2.44 54.385 2.563 ;
      RECT 53.98 2.295 54.26 2.555 ;
      RECT 53.98 2.39 54.36 2.555 ;
      RECT 53.98 2.335 54.305 2.555 ;
      RECT 53.98 2.327 54.3 2.555 ;
      RECT 53.98 2.317 54.295 2.555 ;
      RECT 53.98 2.305 54.29 2.555 ;
      RECT 52.905 3 53.185 3.28 ;
      RECT 52.905 3 53.22 3.26 ;
      RECT 52.94 2.42 52.99 2.68 ;
      RECT 52.73 2.42 52.735 2.68 ;
      RECT 51.925 1.975 51.955 2.235 ;
      RECT 51.695 1.975 51.77 2.235 ;
      RECT 52.915 2.37 52.94 2.68 ;
      RECT 52.91 2.327 52.915 2.68 ;
      RECT 52.905 2.31 52.91 2.68 ;
      RECT 52.9 2.297 52.905 2.68 ;
      RECT 52.825 2.18 52.9 2.68 ;
      RECT 52.78 1.997 52.825 2.68 ;
      RECT 52.775 1.925 52.78 2.68 ;
      RECT 52.76 1.9 52.775 2.68 ;
      RECT 52.735 1.862 52.76 2.68 ;
      RECT 52.725 1.842 52.735 2.402 ;
      RECT 52.71 1.834 52.725 2.357 ;
      RECT 52.705 1.826 52.71 2.328 ;
      RECT 52.7 1.823 52.705 2.308 ;
      RECT 52.695 1.82 52.7 2.288 ;
      RECT 52.69 1.817 52.695 2.268 ;
      RECT 52.66 1.806 52.69 2.205 ;
      RECT 52.64 1.791 52.66 2.12 ;
      RECT 52.635 1.783 52.64 2.083 ;
      RECT 52.625 1.777 52.635 2.05 ;
      RECT 52.61 1.769 52.625 2.01 ;
      RECT 52.605 1.762 52.61 1.97 ;
      RECT 52.6 1.759 52.605 1.948 ;
      RECT 52.595 1.756 52.6 1.935 ;
      RECT 52.59 1.755 52.595 1.925 ;
      RECT 52.575 1.749 52.59 1.915 ;
      RECT 52.55 1.736 52.575 1.9 ;
      RECT 52.5 1.711 52.55 1.871 ;
      RECT 52.485 1.69 52.5 1.846 ;
      RECT 52.475 1.683 52.485 1.835 ;
      RECT 52.42 1.664 52.475 1.808 ;
      RECT 52.395 1.642 52.42 1.781 ;
      RECT 52.39 1.635 52.395 1.776 ;
      RECT 52.375 1.635 52.39 1.774 ;
      RECT 52.35 1.627 52.375 1.77 ;
      RECT 52.335 1.625 52.35 1.766 ;
      RECT 52.305 1.625 52.335 1.763 ;
      RECT 52.295 1.625 52.305 1.758 ;
      RECT 52.25 1.625 52.295 1.756 ;
      RECT 52.221 1.625 52.25 1.757 ;
      RECT 52.135 1.625 52.221 1.759 ;
      RECT 52.121 1.626 52.135 1.761 ;
      RECT 52.035 1.627 52.121 1.763 ;
      RECT 52.02 1.628 52.035 1.773 ;
      RECT 52.015 1.629 52.02 1.782 ;
      RECT 51.995 1.632 52.015 1.792 ;
      RECT 51.98 1.64 51.995 1.807 ;
      RECT 51.96 1.658 51.98 1.822 ;
      RECT 51.95 1.67 51.96 1.845 ;
      RECT 51.94 1.679 51.95 1.875 ;
      RECT 51.925 1.691 51.94 1.92 ;
      RECT 51.87 1.724 51.925 2.235 ;
      RECT 51.865 1.752 51.87 2.235 ;
      RECT 51.845 1.767 51.865 2.235 ;
      RECT 51.81 1.827 51.845 2.235 ;
      RECT 51.808 1.877 51.81 2.235 ;
      RECT 51.805 1.885 51.808 2.235 ;
      RECT 51.795 1.9 51.805 2.235 ;
      RECT 51.79 1.912 51.795 2.235 ;
      RECT 51.78 1.937 51.79 2.235 ;
      RECT 51.77 1.965 51.78 2.235 ;
      RECT 49.675 3.47 49.725 3.73 ;
      RECT 52.585 3.02 52.645 3.28 ;
      RECT 52.57 3.02 52.585 3.29 ;
      RECT 52.551 3.02 52.57 3.323 ;
      RECT 52.465 3.02 52.551 3.448 ;
      RECT 52.385 3.02 52.465 3.63 ;
      RECT 52.38 3.257 52.385 3.715 ;
      RECT 52.355 3.327 52.38 3.743 ;
      RECT 52.35 3.397 52.355 3.77 ;
      RECT 52.33 3.469 52.35 3.792 ;
      RECT 52.325 3.536 52.33 3.815 ;
      RECT 52.315 3.565 52.325 3.83 ;
      RECT 52.305 3.587 52.315 3.847 ;
      RECT 52.3 3.597 52.305 3.858 ;
      RECT 52.295 3.605 52.3 3.866 ;
      RECT 52.285 3.613 52.295 3.878 ;
      RECT 52.28 3.625 52.285 3.888 ;
      RECT 52.275 3.633 52.28 3.893 ;
      RECT 52.255 3.651 52.275 3.903 ;
      RECT 52.25 3.668 52.255 3.91 ;
      RECT 52.245 3.676 52.25 3.911 ;
      RECT 52.24 3.687 52.245 3.913 ;
      RECT 52.2 3.725 52.24 3.923 ;
      RECT 52.195 3.76 52.2 3.934 ;
      RECT 52.19 3.765 52.195 3.937 ;
      RECT 52.165 3.775 52.19 3.944 ;
      RECT 52.155 3.789 52.165 3.953 ;
      RECT 52.135 3.801 52.155 3.956 ;
      RECT 52.085 3.82 52.135 3.96 ;
      RECT 52.04 3.835 52.085 3.965 ;
      RECT 51.975 3.838 52.04 3.971 ;
      RECT 51.96 3.836 51.975 3.978 ;
      RECT 51.93 3.835 51.96 3.978 ;
      RECT 51.891 3.834 51.93 3.974 ;
      RECT 51.805 3.831 51.891 3.97 ;
      RECT 51.788 3.829 51.805 3.967 ;
      RECT 51.702 3.827 51.788 3.964 ;
      RECT 51.616 3.824 51.702 3.958 ;
      RECT 51.53 3.82 51.616 3.953 ;
      RECT 51.452 3.817 51.53 3.949 ;
      RECT 51.366 3.814 51.452 3.947 ;
      RECT 51.28 3.811 51.366 3.944 ;
      RECT 51.222 3.809 51.28 3.941 ;
      RECT 51.136 3.806 51.222 3.939 ;
      RECT 51.05 3.802 51.136 3.937 ;
      RECT 50.964 3.799 51.05 3.934 ;
      RECT 50.878 3.795 50.964 3.932 ;
      RECT 50.792 3.791 50.878 3.929 ;
      RECT 50.706 3.788 50.792 3.927 ;
      RECT 50.62 3.784 50.706 3.924 ;
      RECT 50.534 3.781 50.62 3.922 ;
      RECT 50.448 3.777 50.534 3.919 ;
      RECT 50.362 3.774 50.448 3.917 ;
      RECT 50.276 3.77 50.362 3.914 ;
      RECT 50.19 3.767 50.276 3.912 ;
      RECT 50.18 3.765 50.19 3.908 ;
      RECT 50.175 3.765 50.18 3.906 ;
      RECT 50.135 3.76 50.175 3.9 ;
      RECT 50.121 3.751 50.135 3.893 ;
      RECT 50.035 3.721 50.121 3.878 ;
      RECT 50.015 3.687 50.035 3.863 ;
      RECT 49.945 3.656 50.015 3.85 ;
      RECT 49.94 3.631 49.945 3.839 ;
      RECT 49.935 3.625 49.94 3.837 ;
      RECT 49.866 3.47 49.935 3.825 ;
      RECT 49.78 3.47 49.866 3.799 ;
      RECT 49.755 3.47 49.78 3.778 ;
      RECT 49.75 3.47 49.755 3.768 ;
      RECT 49.745 3.47 49.75 3.76 ;
      RECT 49.725 3.47 49.745 3.743 ;
      RECT 52.145 2.04 52.405 2.3 ;
      RECT 52.13 2.04 52.405 2.203 ;
      RECT 52.1 2.04 52.405 2.178 ;
      RECT 52.065 1.88 52.345 2.16 ;
      RECT 52.035 3.37 52.095 3.63 ;
      RECT 51.06 2.06 51.115 2.32 ;
      RECT 51.995 3.327 52.035 3.63 ;
      RECT 51.966 3.248 51.995 3.63 ;
      RECT 51.88 3.12 51.966 3.63 ;
      RECT 51.86 3 51.88 3.63 ;
      RECT 51.835 2.951 51.86 3.63 ;
      RECT 51.83 2.916 51.835 3.48 ;
      RECT 51.8 2.876 51.83 3.418 ;
      RECT 51.775 2.813 51.8 3.333 ;
      RECT 51.765 2.775 51.775 3.27 ;
      RECT 51.75 2.75 51.765 3.231 ;
      RECT 51.707 2.708 51.75 3.137 ;
      RECT 51.705 2.681 51.707 3.064 ;
      RECT 51.7 2.676 51.705 3.055 ;
      RECT 51.695 2.669 51.7 3.03 ;
      RECT 51.69 2.663 51.695 3.015 ;
      RECT 51.685 2.657 51.69 3.003 ;
      RECT 51.675 2.648 51.685 2.985 ;
      RECT 51.67 2.639 51.675 2.963 ;
      RECT 51.645 2.62 51.67 2.913 ;
      RECT 51.64 2.601 51.645 2.863 ;
      RECT 51.625 2.587 51.64 2.823 ;
      RECT 51.62 2.573 51.625 2.79 ;
      RECT 51.615 2.566 51.62 2.783 ;
      RECT 51.6 2.553 51.615 2.775 ;
      RECT 51.555 2.515 51.6 2.748 ;
      RECT 51.525 2.468 51.555 2.713 ;
      RECT 51.505 2.437 51.525 2.69 ;
      RECT 51.425 2.37 51.505 2.643 ;
      RECT 51.395 2.3 51.425 2.59 ;
      RECT 51.39 2.277 51.395 2.573 ;
      RECT 51.36 2.255 51.39 2.558 ;
      RECT 51.33 2.214 51.36 2.53 ;
      RECT 51.325 2.189 51.33 2.515 ;
      RECT 51.32 2.183 51.325 2.508 ;
      RECT 51.31 2.06 51.32 2.5 ;
      RECT 51.3 2.06 51.31 2.493 ;
      RECT 51.295 2.06 51.3 2.485 ;
      RECT 51.275 2.06 51.295 2.473 ;
      RECT 51.225 2.06 51.275 2.443 ;
      RECT 51.17 2.06 51.225 2.393 ;
      RECT 51.14 2.06 51.17 2.353 ;
      RECT 51.115 2.06 51.14 2.33 ;
      RECT 50.985 2.785 51.265 3.065 ;
      RECT 50.95 2.7 51.21 2.96 ;
      RECT 50.95 2.782 51.22 2.96 ;
      RECT 49.15 2.155 49.155 2.64 ;
      RECT 49.04 2.34 49.045 2.64 ;
      RECT 48.95 2.38 49.015 2.64 ;
      RECT 50.625 1.88 50.715 2.51 ;
      RECT 50.59 1.93 50.595 2.51 ;
      RECT 50.535 1.955 50.545 2.51 ;
      RECT 50.49 1.955 50.5 2.51 ;
      RECT 50.86 1.88 50.905 2.16 ;
      RECT 49.71 1.61 49.91 1.75 ;
      RECT 50.826 1.88 50.86 2.172 ;
      RECT 50.74 1.88 50.826 2.212 ;
      RECT 50.725 1.88 50.74 2.253 ;
      RECT 50.72 1.88 50.725 2.273 ;
      RECT 50.715 1.88 50.72 2.293 ;
      RECT 50.595 1.922 50.625 2.51 ;
      RECT 50.545 1.942 50.59 2.51 ;
      RECT 50.53 1.957 50.535 2.51 ;
      RECT 50.5 1.957 50.53 2.51 ;
      RECT 50.455 1.942 50.49 2.51 ;
      RECT 50.45 1.93 50.455 2.29 ;
      RECT 50.445 1.927 50.45 2.27 ;
      RECT 50.43 1.917 50.445 2.223 ;
      RECT 50.425 1.91 50.43 2.186 ;
      RECT 50.42 1.907 50.425 2.169 ;
      RECT 50.405 1.897 50.42 2.125 ;
      RECT 50.4 1.888 50.405 2.085 ;
      RECT 50.395 1.884 50.4 2.07 ;
      RECT 50.385 1.878 50.395 2.053 ;
      RECT 50.345 1.859 50.385 2.028 ;
      RECT 50.34 1.841 50.345 2.008 ;
      RECT 50.33 1.835 50.34 2.003 ;
      RECT 50.3 1.819 50.33 1.99 ;
      RECT 50.285 1.801 50.3 1.973 ;
      RECT 50.27 1.789 50.285 1.96 ;
      RECT 50.265 1.781 50.27 1.953 ;
      RECT 50.235 1.767 50.265 1.94 ;
      RECT 50.23 1.752 50.235 1.928 ;
      RECT 50.22 1.746 50.23 1.92 ;
      RECT 50.2 1.734 50.22 1.908 ;
      RECT 50.19 1.722 50.2 1.895 ;
      RECT 50.16 1.706 50.19 1.88 ;
      RECT 50.14 1.686 50.16 1.863 ;
      RECT 50.135 1.676 50.14 1.853 ;
      RECT 50.11 1.664 50.135 1.84 ;
      RECT 50.105 1.652 50.11 1.828 ;
      RECT 50.1 1.647 50.105 1.824 ;
      RECT 50.085 1.64 50.1 1.816 ;
      RECT 50.075 1.627 50.085 1.806 ;
      RECT 50.07 1.625 50.075 1.8 ;
      RECT 50.045 1.618 50.07 1.789 ;
      RECT 50.04 1.611 50.045 1.778 ;
      RECT 50.015 1.61 50.04 1.765 ;
      RECT 49.996 1.61 50.015 1.755 ;
      RECT 49.91 1.61 49.996 1.752 ;
      RECT 49.68 1.61 49.71 1.755 ;
      RECT 49.64 1.617 49.68 1.768 ;
      RECT 49.615 1.627 49.64 1.781 ;
      RECT 49.6 1.636 49.615 1.791 ;
      RECT 49.57 1.641 49.6 1.81 ;
      RECT 49.565 1.647 49.57 1.828 ;
      RECT 49.545 1.657 49.565 1.843 ;
      RECT 49.535 1.67 49.545 1.863 ;
      RECT 49.52 1.682 49.535 1.88 ;
      RECT 49.515 1.692 49.52 1.89 ;
      RECT 49.51 1.697 49.515 1.895 ;
      RECT 49.5 1.705 49.51 1.908 ;
      RECT 49.45 1.737 49.5 1.945 ;
      RECT 49.435 1.772 49.45 1.986 ;
      RECT 49.43 1.782 49.435 2.001 ;
      RECT 49.425 1.787 49.43 2.008 ;
      RECT 49.4 1.803 49.425 2.028 ;
      RECT 49.385 1.824 49.4 2.053 ;
      RECT 49.36 1.845 49.385 2.078 ;
      RECT 49.35 1.864 49.36 2.101 ;
      RECT 49.325 1.882 49.35 2.124 ;
      RECT 49.31 1.902 49.325 2.148 ;
      RECT 49.305 1.912 49.31 2.16 ;
      RECT 49.29 1.924 49.305 2.18 ;
      RECT 49.28 1.939 49.29 2.22 ;
      RECT 49.275 1.947 49.28 2.248 ;
      RECT 49.265 1.957 49.275 2.268 ;
      RECT 49.26 1.97 49.265 2.293 ;
      RECT 49.255 1.983 49.26 2.313 ;
      RECT 49.25 1.989 49.255 2.335 ;
      RECT 49.24 1.998 49.25 2.355 ;
      RECT 49.235 2.018 49.24 2.378 ;
      RECT 49.23 2.024 49.235 2.398 ;
      RECT 49.225 2.031 49.23 2.42 ;
      RECT 49.22 2.042 49.225 2.433 ;
      RECT 49.21 2.052 49.22 2.458 ;
      RECT 49.19 2.077 49.21 2.64 ;
      RECT 49.16 2.117 49.19 2.64 ;
      RECT 49.155 2.147 49.16 2.64 ;
      RECT 49.13 2.175 49.15 2.64 ;
      RECT 49.1 2.22 49.13 2.64 ;
      RECT 49.095 2.247 49.1 2.64 ;
      RECT 49.075 2.265 49.095 2.64 ;
      RECT 49.065 2.29 49.075 2.64 ;
      RECT 49.06 2.302 49.065 2.64 ;
      RECT 49.045 2.325 49.06 2.64 ;
      RECT 49.025 2.352 49.04 2.64 ;
      RECT 49.015 2.375 49.025 2.64 ;
      RECT 50.805 3.26 50.885 3.52 ;
      RECT 50.04 2.48 50.11 2.74 ;
      RECT 50.771 3.227 50.805 3.52 ;
      RECT 50.685 3.13 50.771 3.52 ;
      RECT 50.665 3.042 50.685 3.52 ;
      RECT 50.655 3.012 50.665 3.52 ;
      RECT 50.645 2.992 50.655 3.52 ;
      RECT 50.625 2.979 50.645 3.52 ;
      RECT 50.61 2.969 50.625 3.348 ;
      RECT 50.605 2.962 50.61 3.303 ;
      RECT 50.595 2.956 50.605 3.293 ;
      RECT 50.585 2.948 50.595 3.275 ;
      RECT 50.58 2.942 50.585 3.263 ;
      RECT 50.57 2.937 50.58 3.25 ;
      RECT 50.55 2.927 50.57 3.223 ;
      RECT 50.51 2.906 50.55 3.175 ;
      RECT 50.495 2.887 50.51 3.133 ;
      RECT 50.47 2.873 50.495 3.103 ;
      RECT 50.46 2.861 50.47 3.07 ;
      RECT 50.455 2.856 50.46 3.06 ;
      RECT 50.425 2.842 50.455 3.04 ;
      RECT 50.415 2.826 50.425 3.013 ;
      RECT 50.41 2.821 50.415 3.003 ;
      RECT 50.385 2.812 50.41 2.983 ;
      RECT 50.375 2.8 50.385 2.963 ;
      RECT 50.305 2.768 50.375 2.938 ;
      RECT 50.3 2.737 50.305 2.915 ;
      RECT 50.251 2.48 50.3 2.898 ;
      RECT 50.165 2.48 50.251 2.857 ;
      RECT 50.11 2.48 50.165 2.785 ;
      RECT 50.2 3.265 50.36 3.525 ;
      RECT 49.725 1.88 49.775 2.565 ;
      RECT 49.515 2.305 49.55 2.565 ;
      RECT 49.83 1.88 49.835 2.34 ;
      RECT 49.92 1.88 49.945 2.16 ;
      RECT 50.195 3.262 50.2 3.525 ;
      RECT 50.16 3.25 50.195 3.525 ;
      RECT 50.1 3.223 50.16 3.525 ;
      RECT 50.095 3.206 50.1 3.379 ;
      RECT 50.09 3.203 50.095 3.366 ;
      RECT 50.07 3.196 50.09 3.353 ;
      RECT 50.035 3.179 50.07 3.335 ;
      RECT 49.995 3.158 50.035 3.315 ;
      RECT 49.99 3.146 49.995 3.303 ;
      RECT 49.95 3.132 49.99 3.289 ;
      RECT 49.93 3.115 49.95 3.271 ;
      RECT 49.92 3.107 49.93 3.263 ;
      RECT 49.905 1.88 49.92 2.178 ;
      RECT 49.89 3.097 49.92 3.25 ;
      RECT 49.875 1.88 49.905 2.223 ;
      RECT 49.88 3.087 49.89 3.237 ;
      RECT 49.85 3.072 49.88 3.224 ;
      RECT 49.835 1.88 49.875 2.29 ;
      RECT 49.835 3.04 49.85 3.21 ;
      RECT 49.83 3.012 49.835 3.204 ;
      RECT 49.825 1.88 49.83 2.345 ;
      RECT 49.815 2.982 49.83 3.198 ;
      RECT 49.82 1.88 49.825 2.358 ;
      RECT 49.81 1.88 49.82 2.378 ;
      RECT 49.775 2.895 49.815 3.183 ;
      RECT 49.775 1.88 49.81 2.418 ;
      RECT 49.77 2.827 49.775 3.171 ;
      RECT 49.755 2.782 49.77 3.166 ;
      RECT 49.75 2.72 49.755 3.161 ;
      RECT 49.725 2.627 49.75 3.154 ;
      RECT 49.72 1.88 49.725 3.146 ;
      RECT 49.705 1.88 49.72 3.133 ;
      RECT 49.685 1.88 49.705 3.09 ;
      RECT 49.675 1.88 49.685 3.04 ;
      RECT 49.67 1.88 49.675 3.013 ;
      RECT 49.665 1.88 49.67 2.991 ;
      RECT 49.66 2.106 49.665 2.974 ;
      RECT 49.655 2.128 49.66 2.952 ;
      RECT 49.65 2.17 49.655 2.935 ;
      RECT 49.62 2.22 49.65 2.879 ;
      RECT 49.615 2.247 49.62 2.821 ;
      RECT 49.6 2.265 49.615 2.785 ;
      RECT 49.595 2.283 49.6 2.749 ;
      RECT 49.589 2.29 49.595 2.73 ;
      RECT 49.585 2.297 49.589 2.713 ;
      RECT 49.58 2.302 49.585 2.682 ;
      RECT 49.57 2.305 49.58 2.657 ;
      RECT 49.56 2.305 49.57 2.623 ;
      RECT 49.555 2.305 49.56 2.6 ;
      RECT 49.55 2.305 49.555 2.58 ;
      RECT 48.17 3.47 48.43 3.73 ;
      RECT 48.19 3.397 48.37 3.73 ;
      RECT 48.19 3.14 48.365 3.73 ;
      RECT 48.19 2.932 48.355 3.73 ;
      RECT 48.195 2.85 48.355 3.73 ;
      RECT 48.195 2.615 48.345 3.73 ;
      RECT 48.195 2.462 48.34 3.73 ;
      RECT 48.2 2.447 48.34 3.73 ;
      RECT 48.25 2.162 48.34 3.73 ;
      RECT 48.205 2.397 48.34 3.73 ;
      RECT 48.235 2.215 48.34 3.73 ;
      RECT 48.22 2.327 48.34 3.73 ;
      RECT 48.225 2.285 48.34 3.73 ;
      RECT 48.22 2.327 48.355 2.39 ;
      RECT 48.255 1.915 48.36 2.335 ;
      RECT 48.255 1.915 48.375 2.318 ;
      RECT 48.255 1.915 48.41 2.28 ;
      RECT 48.25 2.162 48.46 2.213 ;
      RECT 48.255 1.915 48.515 2.175 ;
      RECT 47.515 2.62 47.775 2.88 ;
      RECT 47.515 2.62 47.785 2.838 ;
      RECT 47.515 2.62 47.871 2.809 ;
      RECT 47.515 2.62 47.94 2.761 ;
      RECT 47.515 2.62 47.975 2.73 ;
      RECT 47.745 2.44 48.025 2.72 ;
      RECT 47.58 2.605 48.025 2.72 ;
      RECT 47.67 2.482 47.775 2.88 ;
      RECT 47.6 2.545 48.025 2.72 ;
      RECT 42.05 6.28 42.37 6.605 ;
      RECT 42.08 5.695 42.25 6.605 ;
      RECT 42.08 5.695 42.255 6.045 ;
      RECT 42.08 5.695 43.055 5.87 ;
      RECT 42.88 1.965 43.055 5.87 ;
      RECT 33.205 2.44 33.485 2.72 ;
      RECT 33.205 2.44 33.505 2.615 ;
      RECT 33.295 2.33 33.555 2.59 ;
      RECT 33.26 2.425 33.555 2.59 ;
      RECT 33.395 0.73 33.55 2.59 ;
      RECT 42.825 1.965 43.175 2.315 ;
      RECT 40.415 2.025 43.175 2.195 ;
      RECT 40.415 0.73 40.585 2.195 ;
      RECT 29.95 1.095 30.29 1.445 ;
      RECT 29.95 1.26 33.55 1.435 ;
      RECT 33.395 0.73 40.585 0.9 ;
      RECT 42.85 6.655 43.175 6.98 ;
      RECT 41.735 6.745 43.175 6.915 ;
      RECT 41.735 2.395 41.895 6.915 ;
      RECT 42.05 2.365 42.37 2.685 ;
      RECT 41.735 2.395 42.37 2.565 ;
      RECT 41 5.86 41.34 6.21 ;
      RECT 41.08 2.705 41.255 6.21 ;
      RECT 41.005 2.705 41.345 3.055 ;
      RECT 40.445 2.705 40.785 3.055 ;
      RECT 39.745 2.77 40.785 2.97 ;
      RECT 39.745 2.765 40.055 2.97 ;
      RECT 39.745 1.04 39.95 2.97 ;
      RECT 40.535 2.7 40.705 3.055 ;
      RECT 34.385 1.04 34.76 1.41 ;
      RECT 34.385 1.04 39.95 1.245 ;
      RECT 38.845 2.44 39.125 2.72 ;
      RECT 38.84 2.44 39.125 2.673 ;
      RECT 38.82 2.44 39.125 2.65 ;
      RECT 38.81 2.44 39.125 2.63 ;
      RECT 38.8 2.44 39.125 2.615 ;
      RECT 38.775 2.44 39.125 2.588 ;
      RECT 38.765 2.44 39.125 2.563 ;
      RECT 38.72 2.295 39 2.555 ;
      RECT 38.72 2.39 39.1 2.555 ;
      RECT 38.72 2.335 39.045 2.555 ;
      RECT 38.72 2.327 39.04 2.555 ;
      RECT 38.72 2.317 39.035 2.555 ;
      RECT 38.72 2.305 39.03 2.555 ;
      RECT 37.645 3 37.925 3.28 ;
      RECT 37.645 3 37.96 3.26 ;
      RECT 37.68 2.42 37.73 2.68 ;
      RECT 37.47 2.42 37.475 2.68 ;
      RECT 36.665 1.975 36.695 2.235 ;
      RECT 36.435 1.975 36.51 2.235 ;
      RECT 37.655 2.37 37.68 2.68 ;
      RECT 37.65 2.327 37.655 2.68 ;
      RECT 37.645 2.31 37.65 2.68 ;
      RECT 37.64 2.297 37.645 2.68 ;
      RECT 37.565 2.18 37.64 2.68 ;
      RECT 37.52 1.997 37.565 2.68 ;
      RECT 37.515 1.925 37.52 2.68 ;
      RECT 37.5 1.9 37.515 2.68 ;
      RECT 37.475 1.862 37.5 2.68 ;
      RECT 37.465 1.842 37.475 2.402 ;
      RECT 37.45 1.834 37.465 2.357 ;
      RECT 37.445 1.826 37.45 2.328 ;
      RECT 37.44 1.823 37.445 2.308 ;
      RECT 37.435 1.82 37.44 2.288 ;
      RECT 37.43 1.817 37.435 2.268 ;
      RECT 37.4 1.806 37.43 2.205 ;
      RECT 37.38 1.791 37.4 2.12 ;
      RECT 37.375 1.783 37.38 2.083 ;
      RECT 37.365 1.777 37.375 2.05 ;
      RECT 37.35 1.769 37.365 2.01 ;
      RECT 37.345 1.762 37.35 1.97 ;
      RECT 37.34 1.759 37.345 1.948 ;
      RECT 37.335 1.756 37.34 1.935 ;
      RECT 37.33 1.755 37.335 1.925 ;
      RECT 37.315 1.749 37.33 1.915 ;
      RECT 37.29 1.736 37.315 1.9 ;
      RECT 37.24 1.711 37.29 1.871 ;
      RECT 37.225 1.69 37.24 1.846 ;
      RECT 37.215 1.683 37.225 1.835 ;
      RECT 37.16 1.664 37.215 1.808 ;
      RECT 37.135 1.642 37.16 1.781 ;
      RECT 37.13 1.635 37.135 1.776 ;
      RECT 37.115 1.635 37.13 1.774 ;
      RECT 37.09 1.627 37.115 1.77 ;
      RECT 37.075 1.625 37.09 1.766 ;
      RECT 37.045 1.625 37.075 1.763 ;
      RECT 37.035 1.625 37.045 1.758 ;
      RECT 36.99 1.625 37.035 1.756 ;
      RECT 36.961 1.625 36.99 1.757 ;
      RECT 36.875 1.625 36.961 1.759 ;
      RECT 36.861 1.626 36.875 1.761 ;
      RECT 36.775 1.627 36.861 1.763 ;
      RECT 36.76 1.628 36.775 1.773 ;
      RECT 36.755 1.629 36.76 1.782 ;
      RECT 36.735 1.632 36.755 1.792 ;
      RECT 36.72 1.64 36.735 1.807 ;
      RECT 36.7 1.658 36.72 1.822 ;
      RECT 36.69 1.67 36.7 1.845 ;
      RECT 36.68 1.679 36.69 1.875 ;
      RECT 36.665 1.691 36.68 1.92 ;
      RECT 36.61 1.724 36.665 2.235 ;
      RECT 36.605 1.752 36.61 2.235 ;
      RECT 36.585 1.767 36.605 2.235 ;
      RECT 36.55 1.827 36.585 2.235 ;
      RECT 36.548 1.877 36.55 2.235 ;
      RECT 36.545 1.885 36.548 2.235 ;
      RECT 36.535 1.9 36.545 2.235 ;
      RECT 36.53 1.912 36.535 2.235 ;
      RECT 36.52 1.937 36.53 2.235 ;
      RECT 36.51 1.965 36.52 2.235 ;
      RECT 34.415 3.47 34.465 3.73 ;
      RECT 37.325 3.02 37.385 3.28 ;
      RECT 37.31 3.02 37.325 3.29 ;
      RECT 37.291 3.02 37.31 3.323 ;
      RECT 37.205 3.02 37.291 3.448 ;
      RECT 37.125 3.02 37.205 3.63 ;
      RECT 37.12 3.257 37.125 3.715 ;
      RECT 37.095 3.327 37.12 3.743 ;
      RECT 37.09 3.397 37.095 3.77 ;
      RECT 37.07 3.469 37.09 3.792 ;
      RECT 37.065 3.536 37.07 3.815 ;
      RECT 37.055 3.565 37.065 3.83 ;
      RECT 37.045 3.587 37.055 3.847 ;
      RECT 37.04 3.597 37.045 3.858 ;
      RECT 37.035 3.605 37.04 3.866 ;
      RECT 37.025 3.613 37.035 3.878 ;
      RECT 37.02 3.625 37.025 3.888 ;
      RECT 37.015 3.633 37.02 3.893 ;
      RECT 36.995 3.651 37.015 3.903 ;
      RECT 36.99 3.668 36.995 3.91 ;
      RECT 36.985 3.676 36.99 3.911 ;
      RECT 36.98 3.687 36.985 3.913 ;
      RECT 36.94 3.725 36.98 3.923 ;
      RECT 36.935 3.76 36.94 3.934 ;
      RECT 36.93 3.765 36.935 3.937 ;
      RECT 36.905 3.775 36.93 3.944 ;
      RECT 36.895 3.789 36.905 3.953 ;
      RECT 36.875 3.801 36.895 3.956 ;
      RECT 36.825 3.82 36.875 3.96 ;
      RECT 36.78 3.835 36.825 3.965 ;
      RECT 36.715 3.838 36.78 3.971 ;
      RECT 36.7 3.836 36.715 3.978 ;
      RECT 36.67 3.835 36.7 3.978 ;
      RECT 36.631 3.834 36.67 3.974 ;
      RECT 36.545 3.831 36.631 3.97 ;
      RECT 36.528 3.829 36.545 3.967 ;
      RECT 36.442 3.827 36.528 3.964 ;
      RECT 36.356 3.824 36.442 3.958 ;
      RECT 36.27 3.82 36.356 3.953 ;
      RECT 36.192 3.817 36.27 3.949 ;
      RECT 36.106 3.814 36.192 3.947 ;
      RECT 36.02 3.811 36.106 3.944 ;
      RECT 35.962 3.809 36.02 3.941 ;
      RECT 35.876 3.806 35.962 3.939 ;
      RECT 35.79 3.802 35.876 3.937 ;
      RECT 35.704 3.799 35.79 3.934 ;
      RECT 35.618 3.795 35.704 3.932 ;
      RECT 35.532 3.791 35.618 3.929 ;
      RECT 35.446 3.788 35.532 3.927 ;
      RECT 35.36 3.784 35.446 3.924 ;
      RECT 35.274 3.781 35.36 3.922 ;
      RECT 35.188 3.777 35.274 3.919 ;
      RECT 35.102 3.774 35.188 3.917 ;
      RECT 35.016 3.77 35.102 3.914 ;
      RECT 34.93 3.767 35.016 3.912 ;
      RECT 34.92 3.765 34.93 3.908 ;
      RECT 34.915 3.765 34.92 3.906 ;
      RECT 34.875 3.76 34.915 3.9 ;
      RECT 34.861 3.751 34.875 3.893 ;
      RECT 34.775 3.721 34.861 3.878 ;
      RECT 34.755 3.687 34.775 3.863 ;
      RECT 34.685 3.656 34.755 3.85 ;
      RECT 34.68 3.631 34.685 3.839 ;
      RECT 34.675 3.625 34.68 3.837 ;
      RECT 34.606 3.47 34.675 3.825 ;
      RECT 34.52 3.47 34.606 3.799 ;
      RECT 34.495 3.47 34.52 3.778 ;
      RECT 34.49 3.47 34.495 3.768 ;
      RECT 34.485 3.47 34.49 3.76 ;
      RECT 34.465 3.47 34.485 3.743 ;
      RECT 36.885 2.04 37.145 2.3 ;
      RECT 36.87 2.04 37.145 2.203 ;
      RECT 36.84 2.04 37.145 2.178 ;
      RECT 36.805 1.88 37.085 2.16 ;
      RECT 36.775 3.37 36.835 3.63 ;
      RECT 35.8 2.06 35.855 2.32 ;
      RECT 36.735 3.327 36.775 3.63 ;
      RECT 36.706 3.248 36.735 3.63 ;
      RECT 36.62 3.12 36.706 3.63 ;
      RECT 36.6 3 36.62 3.63 ;
      RECT 36.575 2.951 36.6 3.63 ;
      RECT 36.57 2.916 36.575 3.48 ;
      RECT 36.54 2.876 36.57 3.418 ;
      RECT 36.515 2.813 36.54 3.333 ;
      RECT 36.505 2.775 36.515 3.27 ;
      RECT 36.49 2.75 36.505 3.231 ;
      RECT 36.447 2.708 36.49 3.137 ;
      RECT 36.445 2.681 36.447 3.064 ;
      RECT 36.44 2.676 36.445 3.055 ;
      RECT 36.435 2.669 36.44 3.03 ;
      RECT 36.43 2.663 36.435 3.015 ;
      RECT 36.425 2.657 36.43 3.003 ;
      RECT 36.415 2.648 36.425 2.985 ;
      RECT 36.41 2.639 36.415 2.963 ;
      RECT 36.385 2.62 36.41 2.913 ;
      RECT 36.38 2.601 36.385 2.863 ;
      RECT 36.365 2.587 36.38 2.823 ;
      RECT 36.36 2.573 36.365 2.79 ;
      RECT 36.355 2.566 36.36 2.783 ;
      RECT 36.34 2.553 36.355 2.775 ;
      RECT 36.295 2.515 36.34 2.748 ;
      RECT 36.265 2.468 36.295 2.713 ;
      RECT 36.245 2.437 36.265 2.69 ;
      RECT 36.165 2.37 36.245 2.643 ;
      RECT 36.135 2.3 36.165 2.59 ;
      RECT 36.13 2.277 36.135 2.573 ;
      RECT 36.1 2.255 36.13 2.558 ;
      RECT 36.07 2.214 36.1 2.53 ;
      RECT 36.065 2.189 36.07 2.515 ;
      RECT 36.06 2.183 36.065 2.508 ;
      RECT 36.05 2.06 36.06 2.5 ;
      RECT 36.04 2.06 36.05 2.493 ;
      RECT 36.035 2.06 36.04 2.485 ;
      RECT 36.015 2.06 36.035 2.473 ;
      RECT 35.965 2.06 36.015 2.443 ;
      RECT 35.91 2.06 35.965 2.393 ;
      RECT 35.88 2.06 35.91 2.353 ;
      RECT 35.855 2.06 35.88 2.33 ;
      RECT 35.725 2.785 36.005 3.065 ;
      RECT 35.69 2.7 35.95 2.96 ;
      RECT 35.69 2.782 35.96 2.96 ;
      RECT 33.89 2.155 33.895 2.64 ;
      RECT 33.78 2.34 33.785 2.64 ;
      RECT 33.69 2.38 33.755 2.64 ;
      RECT 35.365 1.88 35.455 2.51 ;
      RECT 35.33 1.93 35.335 2.51 ;
      RECT 35.275 1.955 35.285 2.51 ;
      RECT 35.23 1.955 35.24 2.51 ;
      RECT 35.6 1.88 35.645 2.16 ;
      RECT 34.45 1.61 34.65 1.75 ;
      RECT 35.566 1.88 35.6 2.172 ;
      RECT 35.48 1.88 35.566 2.212 ;
      RECT 35.465 1.88 35.48 2.253 ;
      RECT 35.46 1.88 35.465 2.273 ;
      RECT 35.455 1.88 35.46 2.293 ;
      RECT 35.335 1.922 35.365 2.51 ;
      RECT 35.285 1.942 35.33 2.51 ;
      RECT 35.27 1.957 35.275 2.51 ;
      RECT 35.24 1.957 35.27 2.51 ;
      RECT 35.195 1.942 35.23 2.51 ;
      RECT 35.19 1.93 35.195 2.29 ;
      RECT 35.185 1.927 35.19 2.27 ;
      RECT 35.17 1.917 35.185 2.223 ;
      RECT 35.165 1.91 35.17 2.186 ;
      RECT 35.16 1.907 35.165 2.169 ;
      RECT 35.145 1.897 35.16 2.125 ;
      RECT 35.14 1.888 35.145 2.085 ;
      RECT 35.135 1.884 35.14 2.07 ;
      RECT 35.125 1.878 35.135 2.053 ;
      RECT 35.085 1.859 35.125 2.028 ;
      RECT 35.08 1.841 35.085 2.008 ;
      RECT 35.07 1.835 35.08 2.003 ;
      RECT 35.04 1.819 35.07 1.99 ;
      RECT 35.025 1.801 35.04 1.973 ;
      RECT 35.01 1.789 35.025 1.96 ;
      RECT 35.005 1.781 35.01 1.953 ;
      RECT 34.975 1.767 35.005 1.94 ;
      RECT 34.97 1.752 34.975 1.928 ;
      RECT 34.96 1.746 34.97 1.92 ;
      RECT 34.94 1.734 34.96 1.908 ;
      RECT 34.93 1.722 34.94 1.895 ;
      RECT 34.9 1.706 34.93 1.88 ;
      RECT 34.88 1.686 34.9 1.863 ;
      RECT 34.875 1.676 34.88 1.853 ;
      RECT 34.85 1.664 34.875 1.84 ;
      RECT 34.845 1.652 34.85 1.828 ;
      RECT 34.84 1.647 34.845 1.824 ;
      RECT 34.825 1.64 34.84 1.816 ;
      RECT 34.815 1.627 34.825 1.806 ;
      RECT 34.81 1.625 34.815 1.8 ;
      RECT 34.785 1.618 34.81 1.789 ;
      RECT 34.78 1.611 34.785 1.778 ;
      RECT 34.755 1.61 34.78 1.765 ;
      RECT 34.736 1.61 34.755 1.755 ;
      RECT 34.65 1.61 34.736 1.752 ;
      RECT 34.42 1.61 34.45 1.755 ;
      RECT 34.38 1.617 34.42 1.768 ;
      RECT 34.355 1.627 34.38 1.781 ;
      RECT 34.34 1.636 34.355 1.791 ;
      RECT 34.31 1.641 34.34 1.81 ;
      RECT 34.305 1.647 34.31 1.828 ;
      RECT 34.285 1.657 34.305 1.843 ;
      RECT 34.275 1.67 34.285 1.863 ;
      RECT 34.26 1.682 34.275 1.88 ;
      RECT 34.255 1.692 34.26 1.89 ;
      RECT 34.25 1.697 34.255 1.895 ;
      RECT 34.24 1.705 34.25 1.908 ;
      RECT 34.19 1.737 34.24 1.945 ;
      RECT 34.175 1.772 34.19 1.986 ;
      RECT 34.17 1.782 34.175 2.001 ;
      RECT 34.165 1.787 34.17 2.008 ;
      RECT 34.14 1.803 34.165 2.028 ;
      RECT 34.125 1.824 34.14 2.053 ;
      RECT 34.1 1.845 34.125 2.078 ;
      RECT 34.09 1.864 34.1 2.101 ;
      RECT 34.065 1.882 34.09 2.124 ;
      RECT 34.05 1.902 34.065 2.148 ;
      RECT 34.045 1.912 34.05 2.16 ;
      RECT 34.03 1.924 34.045 2.18 ;
      RECT 34.02 1.939 34.03 2.22 ;
      RECT 34.015 1.947 34.02 2.248 ;
      RECT 34.005 1.957 34.015 2.268 ;
      RECT 34 1.97 34.005 2.293 ;
      RECT 33.995 1.983 34 2.313 ;
      RECT 33.99 1.989 33.995 2.335 ;
      RECT 33.98 1.998 33.99 2.355 ;
      RECT 33.975 2.018 33.98 2.378 ;
      RECT 33.97 2.024 33.975 2.398 ;
      RECT 33.965 2.031 33.97 2.42 ;
      RECT 33.96 2.042 33.965 2.433 ;
      RECT 33.95 2.052 33.96 2.458 ;
      RECT 33.93 2.077 33.95 2.64 ;
      RECT 33.9 2.117 33.93 2.64 ;
      RECT 33.895 2.147 33.9 2.64 ;
      RECT 33.87 2.175 33.89 2.64 ;
      RECT 33.84 2.22 33.87 2.64 ;
      RECT 33.835 2.247 33.84 2.64 ;
      RECT 33.815 2.265 33.835 2.64 ;
      RECT 33.805 2.29 33.815 2.64 ;
      RECT 33.8 2.302 33.805 2.64 ;
      RECT 33.785 2.325 33.8 2.64 ;
      RECT 33.765 2.352 33.78 2.64 ;
      RECT 33.755 2.375 33.765 2.64 ;
      RECT 35.545 3.26 35.625 3.52 ;
      RECT 34.78 2.48 34.85 2.74 ;
      RECT 35.511 3.227 35.545 3.52 ;
      RECT 35.425 3.13 35.511 3.52 ;
      RECT 35.405 3.042 35.425 3.52 ;
      RECT 35.395 3.012 35.405 3.52 ;
      RECT 35.385 2.992 35.395 3.52 ;
      RECT 35.365 2.979 35.385 3.52 ;
      RECT 35.35 2.969 35.365 3.348 ;
      RECT 35.345 2.962 35.35 3.303 ;
      RECT 35.335 2.956 35.345 3.293 ;
      RECT 35.325 2.948 35.335 3.275 ;
      RECT 35.32 2.942 35.325 3.263 ;
      RECT 35.31 2.937 35.32 3.25 ;
      RECT 35.29 2.927 35.31 3.223 ;
      RECT 35.25 2.906 35.29 3.175 ;
      RECT 35.235 2.887 35.25 3.133 ;
      RECT 35.21 2.873 35.235 3.103 ;
      RECT 35.2 2.861 35.21 3.07 ;
      RECT 35.195 2.856 35.2 3.06 ;
      RECT 35.165 2.842 35.195 3.04 ;
      RECT 35.155 2.826 35.165 3.013 ;
      RECT 35.15 2.821 35.155 3.003 ;
      RECT 35.125 2.812 35.15 2.983 ;
      RECT 35.115 2.8 35.125 2.963 ;
      RECT 35.045 2.768 35.115 2.938 ;
      RECT 35.04 2.737 35.045 2.915 ;
      RECT 34.991 2.48 35.04 2.898 ;
      RECT 34.905 2.48 34.991 2.857 ;
      RECT 34.85 2.48 34.905 2.785 ;
      RECT 34.94 3.265 35.1 3.525 ;
      RECT 34.465 1.88 34.515 2.565 ;
      RECT 34.255 2.305 34.29 2.565 ;
      RECT 34.57 1.88 34.575 2.34 ;
      RECT 34.66 1.88 34.685 2.16 ;
      RECT 34.935 3.262 34.94 3.525 ;
      RECT 34.9 3.25 34.935 3.525 ;
      RECT 34.84 3.223 34.9 3.525 ;
      RECT 34.835 3.206 34.84 3.379 ;
      RECT 34.83 3.203 34.835 3.366 ;
      RECT 34.81 3.196 34.83 3.353 ;
      RECT 34.775 3.179 34.81 3.335 ;
      RECT 34.735 3.158 34.775 3.315 ;
      RECT 34.73 3.146 34.735 3.303 ;
      RECT 34.69 3.132 34.73 3.289 ;
      RECT 34.67 3.115 34.69 3.271 ;
      RECT 34.66 3.107 34.67 3.263 ;
      RECT 34.645 1.88 34.66 2.178 ;
      RECT 34.63 3.097 34.66 3.25 ;
      RECT 34.615 1.88 34.645 2.223 ;
      RECT 34.62 3.087 34.63 3.237 ;
      RECT 34.59 3.072 34.62 3.224 ;
      RECT 34.575 1.88 34.615 2.29 ;
      RECT 34.575 3.04 34.59 3.21 ;
      RECT 34.57 3.012 34.575 3.204 ;
      RECT 34.565 1.88 34.57 2.345 ;
      RECT 34.555 2.982 34.57 3.198 ;
      RECT 34.56 1.88 34.565 2.358 ;
      RECT 34.55 1.88 34.56 2.378 ;
      RECT 34.515 2.895 34.555 3.183 ;
      RECT 34.515 1.88 34.55 2.418 ;
      RECT 34.51 2.827 34.515 3.171 ;
      RECT 34.495 2.782 34.51 3.166 ;
      RECT 34.49 2.72 34.495 3.161 ;
      RECT 34.465 2.627 34.49 3.154 ;
      RECT 34.46 1.88 34.465 3.146 ;
      RECT 34.445 1.88 34.46 3.133 ;
      RECT 34.425 1.88 34.445 3.09 ;
      RECT 34.415 1.88 34.425 3.04 ;
      RECT 34.41 1.88 34.415 3.013 ;
      RECT 34.405 1.88 34.41 2.991 ;
      RECT 34.4 2.106 34.405 2.974 ;
      RECT 34.395 2.128 34.4 2.952 ;
      RECT 34.39 2.17 34.395 2.935 ;
      RECT 34.36 2.22 34.39 2.879 ;
      RECT 34.355 2.247 34.36 2.821 ;
      RECT 34.34 2.265 34.355 2.785 ;
      RECT 34.335 2.283 34.34 2.749 ;
      RECT 34.329 2.29 34.335 2.73 ;
      RECT 34.325 2.297 34.329 2.713 ;
      RECT 34.32 2.302 34.325 2.682 ;
      RECT 34.31 2.305 34.32 2.657 ;
      RECT 34.3 2.305 34.31 2.623 ;
      RECT 34.295 2.305 34.3 2.6 ;
      RECT 34.29 2.305 34.295 2.58 ;
      RECT 32.91 3.47 33.17 3.73 ;
      RECT 32.93 3.397 33.11 3.73 ;
      RECT 32.93 3.14 33.105 3.73 ;
      RECT 32.93 2.932 33.095 3.73 ;
      RECT 32.935 2.85 33.095 3.73 ;
      RECT 32.935 2.615 33.085 3.73 ;
      RECT 32.935 2.462 33.08 3.73 ;
      RECT 32.94 2.447 33.08 3.73 ;
      RECT 32.99 2.162 33.08 3.73 ;
      RECT 32.945 2.397 33.08 3.73 ;
      RECT 32.975 2.215 33.08 3.73 ;
      RECT 32.96 2.327 33.08 3.73 ;
      RECT 32.965 2.285 33.08 3.73 ;
      RECT 32.96 2.327 33.095 2.39 ;
      RECT 32.995 1.915 33.1 2.335 ;
      RECT 32.995 1.915 33.115 2.318 ;
      RECT 32.995 1.915 33.15 2.28 ;
      RECT 32.99 2.162 33.2 2.213 ;
      RECT 32.995 1.915 33.255 2.175 ;
      RECT 32.255 2.62 32.515 2.88 ;
      RECT 32.255 2.62 32.525 2.838 ;
      RECT 32.255 2.62 32.611 2.809 ;
      RECT 32.255 2.62 32.68 2.761 ;
      RECT 32.255 2.62 32.715 2.73 ;
      RECT 32.485 2.44 32.765 2.72 ;
      RECT 32.32 2.605 32.765 2.72 ;
      RECT 32.41 2.482 32.515 2.88 ;
      RECT 32.34 2.545 32.765 2.72 ;
      RECT 26.79 6.28 27.11 6.605 ;
      RECT 26.82 5.695 26.99 6.605 ;
      RECT 26.82 5.695 26.995 6.045 ;
      RECT 26.82 5.695 27.795 5.87 ;
      RECT 27.62 1.965 27.795 5.87 ;
      RECT 17.945 2.44 18.225 2.72 ;
      RECT 17.945 2.44 18.245 2.615 ;
      RECT 18.035 2.33 18.295 2.59 ;
      RECT 18 2.425 18.295 2.59 ;
      RECT 18.135 0.73 18.29 2.59 ;
      RECT 27.565 1.965 27.915 2.315 ;
      RECT 25.155 2.025 27.915 2.195 ;
      RECT 25.155 0.73 25.325 2.195 ;
      RECT 14.69 1.095 15.03 1.445 ;
      RECT 14.69 1.26 18.29 1.42 ;
      RECT 18.135 0.73 25.325 0.9 ;
      RECT 27.59 6.655 27.915 6.98 ;
      RECT 26.475 6.745 27.915 6.915 ;
      RECT 26.475 2.395 26.635 6.915 ;
      RECT 26.79 2.365 27.11 2.685 ;
      RECT 26.475 2.395 27.11 2.565 ;
      RECT 25.74 5.86 26.08 6.21 ;
      RECT 25.82 2.705 25.995 6.21 ;
      RECT 25.745 2.705 26.085 3.055 ;
      RECT 25.185 2.705 25.525 3.055 ;
      RECT 24.485 2.77 25.525 2.97 ;
      RECT 24.485 2.765 24.795 2.97 ;
      RECT 24.485 1.04 24.69 2.97 ;
      RECT 25.275 2.7 25.445 3.055 ;
      RECT 19.125 1.04 19.5 1.41 ;
      RECT 19.125 1.04 24.69 1.245 ;
      RECT 23.585 2.44 23.865 2.72 ;
      RECT 23.58 2.44 23.865 2.673 ;
      RECT 23.56 2.44 23.865 2.65 ;
      RECT 23.55 2.44 23.865 2.63 ;
      RECT 23.54 2.44 23.865 2.615 ;
      RECT 23.515 2.44 23.865 2.588 ;
      RECT 23.505 2.44 23.865 2.563 ;
      RECT 23.46 2.295 23.74 2.555 ;
      RECT 23.46 2.39 23.84 2.555 ;
      RECT 23.46 2.335 23.785 2.555 ;
      RECT 23.46 2.327 23.78 2.555 ;
      RECT 23.46 2.317 23.775 2.555 ;
      RECT 23.46 2.305 23.77 2.555 ;
      RECT 22.385 3 22.665 3.28 ;
      RECT 22.385 3 22.7 3.26 ;
      RECT 22.42 2.42 22.47 2.68 ;
      RECT 22.21 2.42 22.215 2.68 ;
      RECT 21.405 1.975 21.435 2.235 ;
      RECT 21.175 1.975 21.25 2.235 ;
      RECT 22.395 2.37 22.42 2.68 ;
      RECT 22.39 2.327 22.395 2.68 ;
      RECT 22.385 2.31 22.39 2.68 ;
      RECT 22.38 2.297 22.385 2.68 ;
      RECT 22.305 2.18 22.38 2.68 ;
      RECT 22.26 1.997 22.305 2.68 ;
      RECT 22.255 1.925 22.26 2.68 ;
      RECT 22.24 1.9 22.255 2.68 ;
      RECT 22.215 1.862 22.24 2.68 ;
      RECT 22.205 1.842 22.215 2.402 ;
      RECT 22.19 1.834 22.205 2.357 ;
      RECT 22.185 1.826 22.19 2.328 ;
      RECT 22.18 1.823 22.185 2.308 ;
      RECT 22.175 1.82 22.18 2.288 ;
      RECT 22.17 1.817 22.175 2.268 ;
      RECT 22.14 1.806 22.17 2.205 ;
      RECT 22.12 1.791 22.14 2.12 ;
      RECT 22.115 1.783 22.12 2.083 ;
      RECT 22.105 1.777 22.115 2.05 ;
      RECT 22.09 1.769 22.105 2.01 ;
      RECT 22.085 1.762 22.09 1.97 ;
      RECT 22.08 1.759 22.085 1.948 ;
      RECT 22.075 1.756 22.08 1.935 ;
      RECT 22.07 1.755 22.075 1.925 ;
      RECT 22.055 1.749 22.07 1.915 ;
      RECT 22.03 1.736 22.055 1.9 ;
      RECT 21.98 1.711 22.03 1.871 ;
      RECT 21.965 1.69 21.98 1.846 ;
      RECT 21.955 1.683 21.965 1.835 ;
      RECT 21.9 1.664 21.955 1.808 ;
      RECT 21.875 1.642 21.9 1.781 ;
      RECT 21.87 1.635 21.875 1.776 ;
      RECT 21.855 1.635 21.87 1.774 ;
      RECT 21.83 1.627 21.855 1.77 ;
      RECT 21.815 1.625 21.83 1.766 ;
      RECT 21.785 1.625 21.815 1.763 ;
      RECT 21.775 1.625 21.785 1.758 ;
      RECT 21.73 1.625 21.775 1.756 ;
      RECT 21.701 1.625 21.73 1.757 ;
      RECT 21.615 1.625 21.701 1.759 ;
      RECT 21.601 1.626 21.615 1.761 ;
      RECT 21.515 1.627 21.601 1.763 ;
      RECT 21.5 1.628 21.515 1.773 ;
      RECT 21.495 1.629 21.5 1.782 ;
      RECT 21.475 1.632 21.495 1.792 ;
      RECT 21.46 1.64 21.475 1.807 ;
      RECT 21.44 1.658 21.46 1.822 ;
      RECT 21.43 1.67 21.44 1.845 ;
      RECT 21.42 1.679 21.43 1.875 ;
      RECT 21.405 1.691 21.42 1.92 ;
      RECT 21.35 1.724 21.405 2.235 ;
      RECT 21.345 1.752 21.35 2.235 ;
      RECT 21.325 1.767 21.345 2.235 ;
      RECT 21.29 1.827 21.325 2.235 ;
      RECT 21.288 1.877 21.29 2.235 ;
      RECT 21.285 1.885 21.288 2.235 ;
      RECT 21.275 1.9 21.285 2.235 ;
      RECT 21.27 1.912 21.275 2.235 ;
      RECT 21.26 1.937 21.27 2.235 ;
      RECT 21.25 1.965 21.26 2.235 ;
      RECT 19.155 3.47 19.205 3.73 ;
      RECT 22.065 3.02 22.125 3.28 ;
      RECT 22.05 3.02 22.065 3.29 ;
      RECT 22.031 3.02 22.05 3.323 ;
      RECT 21.945 3.02 22.031 3.448 ;
      RECT 21.865 3.02 21.945 3.63 ;
      RECT 21.86 3.257 21.865 3.715 ;
      RECT 21.835 3.327 21.86 3.743 ;
      RECT 21.83 3.397 21.835 3.77 ;
      RECT 21.81 3.469 21.83 3.792 ;
      RECT 21.805 3.536 21.81 3.815 ;
      RECT 21.795 3.565 21.805 3.83 ;
      RECT 21.785 3.587 21.795 3.847 ;
      RECT 21.78 3.597 21.785 3.858 ;
      RECT 21.775 3.605 21.78 3.866 ;
      RECT 21.765 3.613 21.775 3.878 ;
      RECT 21.76 3.625 21.765 3.888 ;
      RECT 21.755 3.633 21.76 3.893 ;
      RECT 21.735 3.651 21.755 3.903 ;
      RECT 21.73 3.668 21.735 3.91 ;
      RECT 21.725 3.676 21.73 3.911 ;
      RECT 21.72 3.687 21.725 3.913 ;
      RECT 21.68 3.725 21.72 3.923 ;
      RECT 21.675 3.76 21.68 3.934 ;
      RECT 21.67 3.765 21.675 3.937 ;
      RECT 21.645 3.775 21.67 3.944 ;
      RECT 21.635 3.789 21.645 3.953 ;
      RECT 21.615 3.801 21.635 3.956 ;
      RECT 21.565 3.82 21.615 3.96 ;
      RECT 21.52 3.835 21.565 3.965 ;
      RECT 21.455 3.838 21.52 3.971 ;
      RECT 21.44 3.836 21.455 3.978 ;
      RECT 21.41 3.835 21.44 3.978 ;
      RECT 21.371 3.834 21.41 3.974 ;
      RECT 21.285 3.831 21.371 3.97 ;
      RECT 21.268 3.829 21.285 3.967 ;
      RECT 21.182 3.827 21.268 3.964 ;
      RECT 21.096 3.824 21.182 3.958 ;
      RECT 21.01 3.82 21.096 3.953 ;
      RECT 20.932 3.817 21.01 3.949 ;
      RECT 20.846 3.814 20.932 3.947 ;
      RECT 20.76 3.811 20.846 3.944 ;
      RECT 20.702 3.809 20.76 3.941 ;
      RECT 20.616 3.806 20.702 3.939 ;
      RECT 20.53 3.802 20.616 3.937 ;
      RECT 20.444 3.799 20.53 3.934 ;
      RECT 20.358 3.795 20.444 3.932 ;
      RECT 20.272 3.791 20.358 3.929 ;
      RECT 20.186 3.788 20.272 3.927 ;
      RECT 20.1 3.784 20.186 3.924 ;
      RECT 20.014 3.781 20.1 3.922 ;
      RECT 19.928 3.777 20.014 3.919 ;
      RECT 19.842 3.774 19.928 3.917 ;
      RECT 19.756 3.77 19.842 3.914 ;
      RECT 19.67 3.767 19.756 3.912 ;
      RECT 19.66 3.765 19.67 3.908 ;
      RECT 19.655 3.765 19.66 3.906 ;
      RECT 19.615 3.76 19.655 3.9 ;
      RECT 19.601 3.751 19.615 3.893 ;
      RECT 19.515 3.721 19.601 3.878 ;
      RECT 19.495 3.687 19.515 3.863 ;
      RECT 19.425 3.656 19.495 3.85 ;
      RECT 19.42 3.631 19.425 3.839 ;
      RECT 19.415 3.625 19.42 3.837 ;
      RECT 19.346 3.47 19.415 3.825 ;
      RECT 19.26 3.47 19.346 3.799 ;
      RECT 19.235 3.47 19.26 3.778 ;
      RECT 19.23 3.47 19.235 3.768 ;
      RECT 19.225 3.47 19.23 3.76 ;
      RECT 19.205 3.47 19.225 3.743 ;
      RECT 21.625 2.04 21.885 2.3 ;
      RECT 21.61 2.04 21.885 2.203 ;
      RECT 21.58 2.04 21.885 2.178 ;
      RECT 21.545 1.88 21.825 2.16 ;
      RECT 21.515 3.37 21.575 3.63 ;
      RECT 20.54 2.06 20.595 2.32 ;
      RECT 21.475 3.327 21.515 3.63 ;
      RECT 21.446 3.248 21.475 3.63 ;
      RECT 21.36 3.12 21.446 3.63 ;
      RECT 21.34 3 21.36 3.63 ;
      RECT 21.315 2.951 21.34 3.63 ;
      RECT 21.31 2.916 21.315 3.48 ;
      RECT 21.28 2.876 21.31 3.418 ;
      RECT 21.255 2.813 21.28 3.333 ;
      RECT 21.245 2.775 21.255 3.27 ;
      RECT 21.23 2.75 21.245 3.231 ;
      RECT 21.187 2.708 21.23 3.137 ;
      RECT 21.185 2.681 21.187 3.064 ;
      RECT 21.18 2.676 21.185 3.055 ;
      RECT 21.175 2.669 21.18 3.03 ;
      RECT 21.17 2.663 21.175 3.015 ;
      RECT 21.165 2.657 21.17 3.003 ;
      RECT 21.155 2.648 21.165 2.985 ;
      RECT 21.15 2.639 21.155 2.963 ;
      RECT 21.125 2.62 21.15 2.913 ;
      RECT 21.12 2.601 21.125 2.863 ;
      RECT 21.105 2.587 21.12 2.823 ;
      RECT 21.1 2.573 21.105 2.79 ;
      RECT 21.095 2.566 21.1 2.783 ;
      RECT 21.08 2.553 21.095 2.775 ;
      RECT 21.035 2.515 21.08 2.748 ;
      RECT 21.005 2.468 21.035 2.713 ;
      RECT 20.985 2.437 21.005 2.69 ;
      RECT 20.905 2.37 20.985 2.643 ;
      RECT 20.875 2.3 20.905 2.59 ;
      RECT 20.87 2.277 20.875 2.573 ;
      RECT 20.84 2.255 20.87 2.558 ;
      RECT 20.81 2.214 20.84 2.53 ;
      RECT 20.805 2.189 20.81 2.515 ;
      RECT 20.8 2.183 20.805 2.508 ;
      RECT 20.79 2.06 20.8 2.5 ;
      RECT 20.78 2.06 20.79 2.493 ;
      RECT 20.775 2.06 20.78 2.485 ;
      RECT 20.755 2.06 20.775 2.473 ;
      RECT 20.705 2.06 20.755 2.443 ;
      RECT 20.65 2.06 20.705 2.393 ;
      RECT 20.62 2.06 20.65 2.353 ;
      RECT 20.595 2.06 20.62 2.33 ;
      RECT 20.465 2.785 20.745 3.065 ;
      RECT 20.43 2.7 20.69 2.96 ;
      RECT 20.43 2.782 20.7 2.96 ;
      RECT 18.63 2.155 18.635 2.64 ;
      RECT 18.52 2.34 18.525 2.64 ;
      RECT 18.43 2.38 18.495 2.64 ;
      RECT 20.105 1.88 20.195 2.51 ;
      RECT 20.07 1.93 20.075 2.51 ;
      RECT 20.015 1.955 20.025 2.51 ;
      RECT 19.97 1.955 19.98 2.51 ;
      RECT 20.34 1.88 20.385 2.16 ;
      RECT 19.19 1.61 19.39 1.75 ;
      RECT 20.306 1.88 20.34 2.172 ;
      RECT 20.22 1.88 20.306 2.212 ;
      RECT 20.205 1.88 20.22 2.253 ;
      RECT 20.2 1.88 20.205 2.273 ;
      RECT 20.195 1.88 20.2 2.293 ;
      RECT 20.075 1.922 20.105 2.51 ;
      RECT 20.025 1.942 20.07 2.51 ;
      RECT 20.01 1.957 20.015 2.51 ;
      RECT 19.98 1.957 20.01 2.51 ;
      RECT 19.935 1.942 19.97 2.51 ;
      RECT 19.93 1.93 19.935 2.29 ;
      RECT 19.925 1.927 19.93 2.27 ;
      RECT 19.91 1.917 19.925 2.223 ;
      RECT 19.905 1.91 19.91 2.186 ;
      RECT 19.9 1.907 19.905 2.169 ;
      RECT 19.885 1.897 19.9 2.125 ;
      RECT 19.88 1.888 19.885 2.085 ;
      RECT 19.875 1.884 19.88 2.07 ;
      RECT 19.865 1.878 19.875 2.053 ;
      RECT 19.825 1.859 19.865 2.028 ;
      RECT 19.82 1.841 19.825 2.008 ;
      RECT 19.81 1.835 19.82 2.003 ;
      RECT 19.78 1.819 19.81 1.99 ;
      RECT 19.765 1.801 19.78 1.973 ;
      RECT 19.75 1.789 19.765 1.96 ;
      RECT 19.745 1.781 19.75 1.953 ;
      RECT 19.715 1.767 19.745 1.94 ;
      RECT 19.71 1.752 19.715 1.928 ;
      RECT 19.7 1.746 19.71 1.92 ;
      RECT 19.68 1.734 19.7 1.908 ;
      RECT 19.67 1.722 19.68 1.895 ;
      RECT 19.64 1.706 19.67 1.88 ;
      RECT 19.62 1.686 19.64 1.863 ;
      RECT 19.615 1.676 19.62 1.853 ;
      RECT 19.59 1.664 19.615 1.84 ;
      RECT 19.585 1.652 19.59 1.828 ;
      RECT 19.58 1.647 19.585 1.824 ;
      RECT 19.565 1.64 19.58 1.816 ;
      RECT 19.555 1.627 19.565 1.806 ;
      RECT 19.55 1.625 19.555 1.8 ;
      RECT 19.525 1.618 19.55 1.789 ;
      RECT 19.52 1.611 19.525 1.778 ;
      RECT 19.495 1.61 19.52 1.765 ;
      RECT 19.476 1.61 19.495 1.755 ;
      RECT 19.39 1.61 19.476 1.752 ;
      RECT 19.16 1.61 19.19 1.755 ;
      RECT 19.12 1.617 19.16 1.768 ;
      RECT 19.095 1.627 19.12 1.781 ;
      RECT 19.08 1.636 19.095 1.791 ;
      RECT 19.05 1.641 19.08 1.81 ;
      RECT 19.045 1.647 19.05 1.828 ;
      RECT 19.025 1.657 19.045 1.843 ;
      RECT 19.015 1.67 19.025 1.863 ;
      RECT 19 1.682 19.015 1.88 ;
      RECT 18.995 1.692 19 1.89 ;
      RECT 18.99 1.697 18.995 1.895 ;
      RECT 18.98 1.705 18.99 1.908 ;
      RECT 18.93 1.737 18.98 1.945 ;
      RECT 18.915 1.772 18.93 1.986 ;
      RECT 18.91 1.782 18.915 2.001 ;
      RECT 18.905 1.787 18.91 2.008 ;
      RECT 18.88 1.803 18.905 2.028 ;
      RECT 18.865 1.824 18.88 2.053 ;
      RECT 18.84 1.845 18.865 2.078 ;
      RECT 18.83 1.864 18.84 2.101 ;
      RECT 18.805 1.882 18.83 2.124 ;
      RECT 18.79 1.902 18.805 2.148 ;
      RECT 18.785 1.912 18.79 2.16 ;
      RECT 18.77 1.924 18.785 2.18 ;
      RECT 18.76 1.939 18.77 2.22 ;
      RECT 18.755 1.947 18.76 2.248 ;
      RECT 18.745 1.957 18.755 2.268 ;
      RECT 18.74 1.97 18.745 2.293 ;
      RECT 18.735 1.983 18.74 2.313 ;
      RECT 18.73 1.989 18.735 2.335 ;
      RECT 18.72 1.998 18.73 2.355 ;
      RECT 18.715 2.018 18.72 2.378 ;
      RECT 18.71 2.024 18.715 2.398 ;
      RECT 18.705 2.031 18.71 2.42 ;
      RECT 18.7 2.042 18.705 2.433 ;
      RECT 18.69 2.052 18.7 2.458 ;
      RECT 18.67 2.077 18.69 2.64 ;
      RECT 18.64 2.117 18.67 2.64 ;
      RECT 18.635 2.147 18.64 2.64 ;
      RECT 18.61 2.175 18.63 2.64 ;
      RECT 18.58 2.22 18.61 2.64 ;
      RECT 18.575 2.247 18.58 2.64 ;
      RECT 18.555 2.265 18.575 2.64 ;
      RECT 18.545 2.29 18.555 2.64 ;
      RECT 18.54 2.302 18.545 2.64 ;
      RECT 18.525 2.325 18.54 2.64 ;
      RECT 18.505 2.352 18.52 2.64 ;
      RECT 18.495 2.375 18.505 2.64 ;
      RECT 20.285 3.26 20.365 3.52 ;
      RECT 19.52 2.48 19.59 2.74 ;
      RECT 20.251 3.227 20.285 3.52 ;
      RECT 20.165 3.13 20.251 3.52 ;
      RECT 20.145 3.042 20.165 3.52 ;
      RECT 20.135 3.012 20.145 3.52 ;
      RECT 20.125 2.992 20.135 3.52 ;
      RECT 20.105 2.979 20.125 3.52 ;
      RECT 20.09 2.969 20.105 3.348 ;
      RECT 20.085 2.962 20.09 3.303 ;
      RECT 20.075 2.956 20.085 3.293 ;
      RECT 20.065 2.948 20.075 3.275 ;
      RECT 20.06 2.942 20.065 3.263 ;
      RECT 20.05 2.937 20.06 3.25 ;
      RECT 20.03 2.927 20.05 3.223 ;
      RECT 19.99 2.906 20.03 3.175 ;
      RECT 19.975 2.887 19.99 3.133 ;
      RECT 19.95 2.873 19.975 3.103 ;
      RECT 19.94 2.861 19.95 3.07 ;
      RECT 19.935 2.856 19.94 3.06 ;
      RECT 19.905 2.842 19.935 3.04 ;
      RECT 19.895 2.826 19.905 3.013 ;
      RECT 19.89 2.821 19.895 3.003 ;
      RECT 19.865 2.812 19.89 2.983 ;
      RECT 19.855 2.8 19.865 2.963 ;
      RECT 19.785 2.768 19.855 2.938 ;
      RECT 19.78 2.737 19.785 2.915 ;
      RECT 19.731 2.48 19.78 2.898 ;
      RECT 19.645 2.48 19.731 2.857 ;
      RECT 19.59 2.48 19.645 2.785 ;
      RECT 19.68 3.265 19.84 3.525 ;
      RECT 19.205 1.88 19.255 2.565 ;
      RECT 18.995 2.305 19.03 2.565 ;
      RECT 19.31 1.88 19.315 2.34 ;
      RECT 19.4 1.88 19.425 2.16 ;
      RECT 19.675 3.262 19.68 3.525 ;
      RECT 19.64 3.25 19.675 3.525 ;
      RECT 19.58 3.223 19.64 3.525 ;
      RECT 19.575 3.206 19.58 3.379 ;
      RECT 19.57 3.203 19.575 3.366 ;
      RECT 19.55 3.196 19.57 3.353 ;
      RECT 19.515 3.179 19.55 3.335 ;
      RECT 19.475 3.158 19.515 3.315 ;
      RECT 19.47 3.146 19.475 3.303 ;
      RECT 19.43 3.132 19.47 3.289 ;
      RECT 19.41 3.115 19.43 3.271 ;
      RECT 19.4 3.107 19.41 3.263 ;
      RECT 19.385 1.88 19.4 2.178 ;
      RECT 19.37 3.097 19.4 3.25 ;
      RECT 19.355 1.88 19.385 2.223 ;
      RECT 19.36 3.087 19.37 3.237 ;
      RECT 19.33 3.072 19.36 3.224 ;
      RECT 19.315 1.88 19.355 2.29 ;
      RECT 19.315 3.04 19.33 3.21 ;
      RECT 19.31 3.012 19.315 3.204 ;
      RECT 19.305 1.88 19.31 2.345 ;
      RECT 19.295 2.982 19.31 3.198 ;
      RECT 19.3 1.88 19.305 2.358 ;
      RECT 19.29 1.88 19.3 2.378 ;
      RECT 19.255 2.895 19.295 3.183 ;
      RECT 19.255 1.88 19.29 2.418 ;
      RECT 19.25 2.827 19.255 3.171 ;
      RECT 19.235 2.782 19.25 3.166 ;
      RECT 19.23 2.72 19.235 3.161 ;
      RECT 19.205 2.627 19.23 3.154 ;
      RECT 19.2 1.88 19.205 3.146 ;
      RECT 19.185 1.88 19.2 3.133 ;
      RECT 19.165 1.88 19.185 3.09 ;
      RECT 19.155 1.88 19.165 3.04 ;
      RECT 19.15 1.88 19.155 3.013 ;
      RECT 19.145 1.88 19.15 2.991 ;
      RECT 19.14 2.106 19.145 2.974 ;
      RECT 19.135 2.128 19.14 2.952 ;
      RECT 19.13 2.17 19.135 2.935 ;
      RECT 19.1 2.22 19.13 2.879 ;
      RECT 19.095 2.247 19.1 2.821 ;
      RECT 19.08 2.265 19.095 2.785 ;
      RECT 19.075 2.283 19.08 2.749 ;
      RECT 19.069 2.29 19.075 2.73 ;
      RECT 19.065 2.297 19.069 2.713 ;
      RECT 19.06 2.302 19.065 2.682 ;
      RECT 19.05 2.305 19.06 2.657 ;
      RECT 19.04 2.305 19.05 2.623 ;
      RECT 19.035 2.305 19.04 2.6 ;
      RECT 19.03 2.305 19.035 2.58 ;
      RECT 17.65 3.47 17.91 3.73 ;
      RECT 17.67 3.397 17.85 3.73 ;
      RECT 17.67 3.14 17.845 3.73 ;
      RECT 17.67 2.932 17.835 3.73 ;
      RECT 17.675 2.85 17.835 3.73 ;
      RECT 17.675 2.615 17.825 3.73 ;
      RECT 17.675 2.462 17.82 3.73 ;
      RECT 17.68 2.447 17.82 3.73 ;
      RECT 17.73 2.162 17.82 3.73 ;
      RECT 17.685 2.397 17.82 3.73 ;
      RECT 17.715 2.215 17.82 3.73 ;
      RECT 17.7 2.327 17.82 3.73 ;
      RECT 17.705 2.285 17.82 3.73 ;
      RECT 17.7 2.327 17.835 2.39 ;
      RECT 17.735 1.915 17.84 2.335 ;
      RECT 17.735 1.915 17.855 2.318 ;
      RECT 17.735 1.915 17.89 2.28 ;
      RECT 17.73 2.162 17.94 2.213 ;
      RECT 17.735 1.915 17.995 2.175 ;
      RECT 16.995 2.62 17.255 2.88 ;
      RECT 16.995 2.62 17.265 2.838 ;
      RECT 16.995 2.62 17.351 2.809 ;
      RECT 16.995 2.62 17.42 2.761 ;
      RECT 16.995 2.62 17.455 2.73 ;
      RECT 17.225 2.44 17.505 2.72 ;
      RECT 17.06 2.605 17.505 2.72 ;
      RECT 17.15 2.482 17.255 2.88 ;
      RECT 17.08 2.545 17.505 2.72 ;
      RECT 12.33 6.655 12.655 6.98 ;
      RECT 11.215 6.745 12.655 6.915 ;
      RECT 11.215 2.395 11.375 6.915 ;
      RECT 11.53 2.365 11.85 2.685 ;
      RECT 11.215 2.395 11.85 2.565 ;
      RECT 10.48 5.86 10.82 6.21 ;
      RECT 10.56 2.705 10.735 6.21 ;
      RECT 10.485 2.705 10.825 3.055 ;
      RECT 9.925 2.705 10.265 3.055 ;
      RECT 9.225 2.77 10.265 2.97 ;
      RECT 9.225 2.765 9.535 2.97 ;
      RECT 9.225 1.04 9.43 2.97 ;
      RECT 10.015 2.7 10.185 3.055 ;
      RECT 3.865 1.04 4.24 1.41 ;
      RECT 3.865 1.04 9.43 1.245 ;
      RECT 8.325 2.44 8.605 2.72 ;
      RECT 8.32 2.44 8.605 2.673 ;
      RECT 8.3 2.44 8.605 2.65 ;
      RECT 8.29 2.44 8.605 2.63 ;
      RECT 8.28 2.44 8.605 2.615 ;
      RECT 8.255 2.44 8.605 2.588 ;
      RECT 8.245 2.44 8.605 2.563 ;
      RECT 8.2 2.295 8.48 2.555 ;
      RECT 8.2 2.39 8.58 2.555 ;
      RECT 8.2 2.335 8.525 2.555 ;
      RECT 8.2 2.327 8.52 2.555 ;
      RECT 8.2 2.317 8.515 2.555 ;
      RECT 8.2 2.305 8.51 2.555 ;
      RECT 7.125 3 7.405 3.28 ;
      RECT 7.125 3 7.44 3.26 ;
      RECT 7.16 2.42 7.21 2.68 ;
      RECT 6.95 2.42 6.955 2.68 ;
      RECT 6.145 1.975 6.175 2.235 ;
      RECT 5.915 1.975 5.99 2.235 ;
      RECT 7.135 2.37 7.16 2.68 ;
      RECT 7.13 2.327 7.135 2.68 ;
      RECT 7.125 2.31 7.13 2.68 ;
      RECT 7.12 2.297 7.125 2.68 ;
      RECT 7.045 2.18 7.12 2.68 ;
      RECT 7 1.997 7.045 2.68 ;
      RECT 6.995 1.925 7 2.68 ;
      RECT 6.98 1.9 6.995 2.68 ;
      RECT 6.955 1.862 6.98 2.68 ;
      RECT 6.945 1.842 6.955 2.402 ;
      RECT 6.93 1.834 6.945 2.357 ;
      RECT 6.925 1.826 6.93 2.328 ;
      RECT 6.92 1.823 6.925 2.308 ;
      RECT 6.915 1.82 6.92 2.288 ;
      RECT 6.91 1.817 6.915 2.268 ;
      RECT 6.88 1.806 6.91 2.205 ;
      RECT 6.86 1.791 6.88 2.12 ;
      RECT 6.855 1.783 6.86 2.083 ;
      RECT 6.845 1.777 6.855 2.05 ;
      RECT 6.83 1.769 6.845 2.01 ;
      RECT 6.825 1.762 6.83 1.97 ;
      RECT 6.82 1.759 6.825 1.948 ;
      RECT 6.815 1.756 6.82 1.935 ;
      RECT 6.81 1.755 6.815 1.925 ;
      RECT 6.795 1.749 6.81 1.915 ;
      RECT 6.77 1.736 6.795 1.9 ;
      RECT 6.72 1.711 6.77 1.871 ;
      RECT 6.705 1.69 6.72 1.846 ;
      RECT 6.695 1.683 6.705 1.835 ;
      RECT 6.64 1.664 6.695 1.808 ;
      RECT 6.615 1.642 6.64 1.781 ;
      RECT 6.61 1.635 6.615 1.776 ;
      RECT 6.595 1.635 6.61 1.774 ;
      RECT 6.57 1.627 6.595 1.77 ;
      RECT 6.555 1.625 6.57 1.766 ;
      RECT 6.525 1.625 6.555 1.763 ;
      RECT 6.515 1.625 6.525 1.758 ;
      RECT 6.47 1.625 6.515 1.756 ;
      RECT 6.441 1.625 6.47 1.757 ;
      RECT 6.355 1.625 6.441 1.759 ;
      RECT 6.341 1.626 6.355 1.761 ;
      RECT 6.255 1.627 6.341 1.763 ;
      RECT 6.24 1.628 6.255 1.773 ;
      RECT 6.235 1.629 6.24 1.782 ;
      RECT 6.215 1.632 6.235 1.792 ;
      RECT 6.2 1.64 6.215 1.807 ;
      RECT 6.18 1.658 6.2 1.822 ;
      RECT 6.17 1.67 6.18 1.845 ;
      RECT 6.16 1.679 6.17 1.875 ;
      RECT 6.145 1.691 6.16 1.92 ;
      RECT 6.09 1.724 6.145 2.235 ;
      RECT 6.085 1.752 6.09 2.235 ;
      RECT 6.065 1.767 6.085 2.235 ;
      RECT 6.03 1.827 6.065 2.235 ;
      RECT 6.028 1.877 6.03 2.235 ;
      RECT 6.025 1.885 6.028 2.235 ;
      RECT 6.015 1.9 6.025 2.235 ;
      RECT 6.01 1.912 6.015 2.235 ;
      RECT 6 1.937 6.01 2.235 ;
      RECT 5.99 1.965 6 2.235 ;
      RECT 3.895 3.47 3.945 3.73 ;
      RECT 6.805 3.02 6.865 3.28 ;
      RECT 6.79 3.02 6.805 3.29 ;
      RECT 6.771 3.02 6.79 3.323 ;
      RECT 6.685 3.02 6.771 3.448 ;
      RECT 6.605 3.02 6.685 3.63 ;
      RECT 6.6 3.257 6.605 3.715 ;
      RECT 6.575 3.327 6.6 3.743 ;
      RECT 6.57 3.397 6.575 3.77 ;
      RECT 6.55 3.469 6.57 3.792 ;
      RECT 6.545 3.536 6.55 3.815 ;
      RECT 6.535 3.565 6.545 3.83 ;
      RECT 6.525 3.587 6.535 3.847 ;
      RECT 6.52 3.597 6.525 3.858 ;
      RECT 6.515 3.605 6.52 3.866 ;
      RECT 6.505 3.613 6.515 3.878 ;
      RECT 6.5 3.625 6.505 3.888 ;
      RECT 6.495 3.633 6.5 3.893 ;
      RECT 6.475 3.651 6.495 3.903 ;
      RECT 6.47 3.668 6.475 3.91 ;
      RECT 6.465 3.676 6.47 3.911 ;
      RECT 6.46 3.687 6.465 3.913 ;
      RECT 6.42 3.725 6.46 3.923 ;
      RECT 6.415 3.76 6.42 3.934 ;
      RECT 6.41 3.765 6.415 3.937 ;
      RECT 6.385 3.775 6.41 3.944 ;
      RECT 6.375 3.789 6.385 3.953 ;
      RECT 6.355 3.801 6.375 3.956 ;
      RECT 6.305 3.82 6.355 3.96 ;
      RECT 6.26 3.835 6.305 3.965 ;
      RECT 6.195 3.838 6.26 3.971 ;
      RECT 6.18 3.836 6.195 3.978 ;
      RECT 6.15 3.835 6.18 3.978 ;
      RECT 6.111 3.834 6.15 3.974 ;
      RECT 6.025 3.831 6.111 3.97 ;
      RECT 6.008 3.829 6.025 3.967 ;
      RECT 5.922 3.827 6.008 3.964 ;
      RECT 5.836 3.824 5.922 3.958 ;
      RECT 5.75 3.82 5.836 3.953 ;
      RECT 5.672 3.817 5.75 3.949 ;
      RECT 5.586 3.814 5.672 3.947 ;
      RECT 5.5 3.811 5.586 3.944 ;
      RECT 5.442 3.809 5.5 3.941 ;
      RECT 5.356 3.806 5.442 3.939 ;
      RECT 5.27 3.802 5.356 3.937 ;
      RECT 5.184 3.799 5.27 3.934 ;
      RECT 5.098 3.795 5.184 3.932 ;
      RECT 5.012 3.791 5.098 3.929 ;
      RECT 4.926 3.788 5.012 3.927 ;
      RECT 4.84 3.784 4.926 3.924 ;
      RECT 4.754 3.781 4.84 3.922 ;
      RECT 4.668 3.777 4.754 3.919 ;
      RECT 4.582 3.774 4.668 3.917 ;
      RECT 4.496 3.77 4.582 3.914 ;
      RECT 4.41 3.767 4.496 3.912 ;
      RECT 4.4 3.765 4.41 3.908 ;
      RECT 4.395 3.765 4.4 3.906 ;
      RECT 4.355 3.76 4.395 3.9 ;
      RECT 4.341 3.751 4.355 3.893 ;
      RECT 4.255 3.721 4.341 3.878 ;
      RECT 4.235 3.687 4.255 3.863 ;
      RECT 4.165 3.656 4.235 3.85 ;
      RECT 4.16 3.631 4.165 3.839 ;
      RECT 4.155 3.625 4.16 3.837 ;
      RECT 4.086 3.47 4.155 3.825 ;
      RECT 4 3.47 4.086 3.799 ;
      RECT 3.975 3.47 4 3.778 ;
      RECT 3.97 3.47 3.975 3.768 ;
      RECT 3.965 3.47 3.97 3.76 ;
      RECT 3.945 3.47 3.965 3.743 ;
      RECT 6.365 2.04 6.625 2.3 ;
      RECT 6.35 2.04 6.625 2.203 ;
      RECT 6.32 2.04 6.625 2.178 ;
      RECT 6.285 1.88 6.565 2.16 ;
      RECT 6.255 3.37 6.315 3.63 ;
      RECT 5.28 2.06 5.335 2.32 ;
      RECT 6.215 3.327 6.255 3.63 ;
      RECT 6.186 3.248 6.215 3.63 ;
      RECT 6.1 3.12 6.186 3.63 ;
      RECT 6.08 3 6.1 3.63 ;
      RECT 6.055 2.951 6.08 3.63 ;
      RECT 6.05 2.916 6.055 3.48 ;
      RECT 6.02 2.876 6.05 3.418 ;
      RECT 5.995 2.813 6.02 3.333 ;
      RECT 5.985 2.775 5.995 3.27 ;
      RECT 5.97 2.75 5.985 3.231 ;
      RECT 5.927 2.708 5.97 3.137 ;
      RECT 5.925 2.681 5.927 3.064 ;
      RECT 5.92 2.676 5.925 3.055 ;
      RECT 5.915 2.669 5.92 3.03 ;
      RECT 5.91 2.663 5.915 3.015 ;
      RECT 5.905 2.657 5.91 3.003 ;
      RECT 5.895 2.648 5.905 2.985 ;
      RECT 5.89 2.639 5.895 2.963 ;
      RECT 5.865 2.62 5.89 2.913 ;
      RECT 5.86 2.601 5.865 2.863 ;
      RECT 5.845 2.587 5.86 2.823 ;
      RECT 5.84 2.573 5.845 2.79 ;
      RECT 5.835 2.566 5.84 2.783 ;
      RECT 5.82 2.553 5.835 2.775 ;
      RECT 5.775 2.515 5.82 2.748 ;
      RECT 5.745 2.468 5.775 2.713 ;
      RECT 5.725 2.437 5.745 2.69 ;
      RECT 5.645 2.37 5.725 2.643 ;
      RECT 5.615 2.3 5.645 2.59 ;
      RECT 5.61 2.277 5.615 2.573 ;
      RECT 5.58 2.255 5.61 2.558 ;
      RECT 5.55 2.214 5.58 2.53 ;
      RECT 5.545 2.189 5.55 2.515 ;
      RECT 5.54 2.183 5.545 2.508 ;
      RECT 5.53 2.06 5.54 2.5 ;
      RECT 5.52 2.06 5.53 2.493 ;
      RECT 5.515 2.06 5.52 2.485 ;
      RECT 5.495 2.06 5.515 2.473 ;
      RECT 5.445 2.06 5.495 2.443 ;
      RECT 5.39 2.06 5.445 2.393 ;
      RECT 5.36 2.06 5.39 2.353 ;
      RECT 5.335 2.06 5.36 2.33 ;
      RECT 5.205 2.785 5.485 3.065 ;
      RECT 5.17 2.7 5.43 2.96 ;
      RECT 5.17 2.782 5.44 2.96 ;
      RECT 3.37 2.155 3.375 2.64 ;
      RECT 3.26 2.34 3.265 2.64 ;
      RECT 3.17 2.38 3.235 2.64 ;
      RECT 4.845 1.88 4.935 2.51 ;
      RECT 4.81 1.93 4.815 2.51 ;
      RECT 4.755 1.955 4.765 2.51 ;
      RECT 4.71 1.955 4.72 2.51 ;
      RECT 5.08 1.88 5.125 2.16 ;
      RECT 3.93 1.61 4.13 1.75 ;
      RECT 5.046 1.88 5.08 2.172 ;
      RECT 4.96 1.88 5.046 2.212 ;
      RECT 4.945 1.88 4.96 2.253 ;
      RECT 4.94 1.88 4.945 2.273 ;
      RECT 4.935 1.88 4.94 2.293 ;
      RECT 4.815 1.922 4.845 2.51 ;
      RECT 4.765 1.942 4.81 2.51 ;
      RECT 4.75 1.957 4.755 2.51 ;
      RECT 4.72 1.957 4.75 2.51 ;
      RECT 4.675 1.942 4.71 2.51 ;
      RECT 4.67 1.93 4.675 2.29 ;
      RECT 4.665 1.927 4.67 2.27 ;
      RECT 4.65 1.917 4.665 2.223 ;
      RECT 4.645 1.91 4.65 2.186 ;
      RECT 4.64 1.907 4.645 2.169 ;
      RECT 4.625 1.897 4.64 2.125 ;
      RECT 4.62 1.888 4.625 2.085 ;
      RECT 4.615 1.884 4.62 2.07 ;
      RECT 4.605 1.878 4.615 2.053 ;
      RECT 4.565 1.859 4.605 2.028 ;
      RECT 4.56 1.841 4.565 2.008 ;
      RECT 4.55 1.835 4.56 2.003 ;
      RECT 4.52 1.819 4.55 1.99 ;
      RECT 4.505 1.801 4.52 1.973 ;
      RECT 4.49 1.789 4.505 1.96 ;
      RECT 4.485 1.781 4.49 1.953 ;
      RECT 4.455 1.767 4.485 1.94 ;
      RECT 4.45 1.752 4.455 1.928 ;
      RECT 4.44 1.746 4.45 1.92 ;
      RECT 4.42 1.734 4.44 1.908 ;
      RECT 4.41 1.722 4.42 1.895 ;
      RECT 4.38 1.706 4.41 1.88 ;
      RECT 4.36 1.686 4.38 1.863 ;
      RECT 4.355 1.676 4.36 1.853 ;
      RECT 4.33 1.664 4.355 1.84 ;
      RECT 4.325 1.652 4.33 1.828 ;
      RECT 4.32 1.647 4.325 1.824 ;
      RECT 4.305 1.64 4.32 1.816 ;
      RECT 4.295 1.627 4.305 1.806 ;
      RECT 4.29 1.625 4.295 1.8 ;
      RECT 4.265 1.618 4.29 1.789 ;
      RECT 4.26 1.611 4.265 1.778 ;
      RECT 4.235 1.61 4.26 1.765 ;
      RECT 4.216 1.61 4.235 1.755 ;
      RECT 4.13 1.61 4.216 1.752 ;
      RECT 3.9 1.61 3.93 1.755 ;
      RECT 3.86 1.617 3.9 1.768 ;
      RECT 3.835 1.627 3.86 1.781 ;
      RECT 3.82 1.636 3.835 1.791 ;
      RECT 3.79 1.641 3.82 1.81 ;
      RECT 3.785 1.647 3.79 1.828 ;
      RECT 3.765 1.657 3.785 1.843 ;
      RECT 3.755 1.67 3.765 1.863 ;
      RECT 3.74 1.682 3.755 1.88 ;
      RECT 3.735 1.692 3.74 1.89 ;
      RECT 3.73 1.697 3.735 1.895 ;
      RECT 3.72 1.705 3.73 1.908 ;
      RECT 3.67 1.737 3.72 1.945 ;
      RECT 3.655 1.772 3.67 1.986 ;
      RECT 3.65 1.782 3.655 2.001 ;
      RECT 3.645 1.787 3.65 2.008 ;
      RECT 3.62 1.803 3.645 2.028 ;
      RECT 3.605 1.824 3.62 2.053 ;
      RECT 3.58 1.845 3.605 2.078 ;
      RECT 3.57 1.864 3.58 2.101 ;
      RECT 3.545 1.882 3.57 2.124 ;
      RECT 3.53 1.902 3.545 2.148 ;
      RECT 3.525 1.912 3.53 2.16 ;
      RECT 3.51 1.924 3.525 2.18 ;
      RECT 3.5 1.939 3.51 2.22 ;
      RECT 3.495 1.947 3.5 2.248 ;
      RECT 3.485 1.957 3.495 2.268 ;
      RECT 3.48 1.97 3.485 2.293 ;
      RECT 3.475 1.983 3.48 2.313 ;
      RECT 3.47 1.989 3.475 2.335 ;
      RECT 3.46 1.998 3.47 2.355 ;
      RECT 3.455 2.018 3.46 2.378 ;
      RECT 3.45 2.024 3.455 2.398 ;
      RECT 3.445 2.031 3.45 2.42 ;
      RECT 3.44 2.042 3.445 2.433 ;
      RECT 3.43 2.052 3.44 2.458 ;
      RECT 3.41 2.077 3.43 2.64 ;
      RECT 3.38 2.117 3.41 2.64 ;
      RECT 3.375 2.147 3.38 2.64 ;
      RECT 3.35 2.175 3.37 2.64 ;
      RECT 3.32 2.22 3.35 2.64 ;
      RECT 3.315 2.247 3.32 2.64 ;
      RECT 3.295 2.265 3.315 2.64 ;
      RECT 3.285 2.29 3.295 2.64 ;
      RECT 3.28 2.302 3.285 2.64 ;
      RECT 3.265 2.325 3.28 2.64 ;
      RECT 3.245 2.352 3.26 2.64 ;
      RECT 3.235 2.375 3.245 2.64 ;
      RECT 5.025 3.26 5.105 3.52 ;
      RECT 4.26 2.48 4.33 2.74 ;
      RECT 4.991 3.227 5.025 3.52 ;
      RECT 4.905 3.13 4.991 3.52 ;
      RECT 4.885 3.042 4.905 3.52 ;
      RECT 4.875 3.012 4.885 3.52 ;
      RECT 4.865 2.992 4.875 3.52 ;
      RECT 4.845 2.979 4.865 3.52 ;
      RECT 4.83 2.969 4.845 3.348 ;
      RECT 4.825 2.962 4.83 3.303 ;
      RECT 4.815 2.956 4.825 3.293 ;
      RECT 4.805 2.948 4.815 3.275 ;
      RECT 4.8 2.942 4.805 3.263 ;
      RECT 4.79 2.937 4.8 3.25 ;
      RECT 4.77 2.927 4.79 3.223 ;
      RECT 4.73 2.906 4.77 3.175 ;
      RECT 4.715 2.887 4.73 3.133 ;
      RECT 4.69 2.873 4.715 3.103 ;
      RECT 4.68 2.861 4.69 3.07 ;
      RECT 4.675 2.856 4.68 3.06 ;
      RECT 4.645 2.842 4.675 3.04 ;
      RECT 4.635 2.826 4.645 3.013 ;
      RECT 4.63 2.821 4.635 3.003 ;
      RECT 4.605 2.812 4.63 2.983 ;
      RECT 4.595 2.8 4.605 2.963 ;
      RECT 4.525 2.768 4.595 2.938 ;
      RECT 4.52 2.737 4.525 2.915 ;
      RECT 4.471 2.48 4.52 2.898 ;
      RECT 4.385 2.48 4.471 2.857 ;
      RECT 4.33 2.48 4.385 2.785 ;
      RECT 4.42 3.265 4.58 3.525 ;
      RECT 3.945 1.88 3.995 2.565 ;
      RECT 3.735 2.305 3.77 2.565 ;
      RECT 4.05 1.88 4.055 2.34 ;
      RECT 4.14 1.88 4.165 2.16 ;
      RECT 4.415 3.262 4.42 3.525 ;
      RECT 4.38 3.25 4.415 3.525 ;
      RECT 4.32 3.223 4.38 3.525 ;
      RECT 4.315 3.206 4.32 3.379 ;
      RECT 4.31 3.203 4.315 3.366 ;
      RECT 4.29 3.196 4.31 3.353 ;
      RECT 4.255 3.179 4.29 3.335 ;
      RECT 4.215 3.158 4.255 3.315 ;
      RECT 4.21 3.146 4.215 3.303 ;
      RECT 4.17 3.132 4.21 3.289 ;
      RECT 4.15 3.115 4.17 3.271 ;
      RECT 4.14 3.107 4.15 3.263 ;
      RECT 4.125 1.88 4.14 2.178 ;
      RECT 4.11 3.097 4.14 3.25 ;
      RECT 4.095 1.88 4.125 2.223 ;
      RECT 4.1 3.087 4.11 3.237 ;
      RECT 4.07 3.072 4.1 3.224 ;
      RECT 4.055 1.88 4.095 2.29 ;
      RECT 4.055 3.04 4.07 3.21 ;
      RECT 4.05 3.012 4.055 3.204 ;
      RECT 4.045 1.88 4.05 2.345 ;
      RECT 4.035 2.982 4.05 3.198 ;
      RECT 4.04 1.88 4.045 2.358 ;
      RECT 4.03 1.88 4.04 2.378 ;
      RECT 3.995 2.895 4.035 3.183 ;
      RECT 3.995 1.88 4.03 2.418 ;
      RECT 3.99 2.827 3.995 3.171 ;
      RECT 3.975 2.782 3.99 3.166 ;
      RECT 3.97 2.72 3.975 3.161 ;
      RECT 3.945 2.627 3.97 3.154 ;
      RECT 3.94 1.88 3.945 3.146 ;
      RECT 3.925 1.88 3.94 3.133 ;
      RECT 3.905 1.88 3.925 3.09 ;
      RECT 3.895 1.88 3.905 3.04 ;
      RECT 3.89 1.88 3.895 3.013 ;
      RECT 3.885 1.88 3.89 2.991 ;
      RECT 3.88 2.106 3.885 2.974 ;
      RECT 3.875 2.128 3.88 2.952 ;
      RECT 3.87 2.17 3.875 2.935 ;
      RECT 3.84 2.22 3.87 2.879 ;
      RECT 3.835 2.247 3.84 2.821 ;
      RECT 3.82 2.265 3.835 2.785 ;
      RECT 3.815 2.283 3.82 2.749 ;
      RECT 3.809 2.29 3.815 2.73 ;
      RECT 3.805 2.297 3.809 2.713 ;
      RECT 3.8 2.302 3.805 2.682 ;
      RECT 3.79 2.305 3.8 2.657 ;
      RECT 3.78 2.305 3.79 2.623 ;
      RECT 3.775 2.305 3.78 2.6 ;
      RECT 3.77 2.305 3.775 2.58 ;
      RECT 2.39 3.47 2.65 3.73 ;
      RECT 2.41 3.397 2.59 3.73 ;
      RECT 2.41 3.14 2.585 3.73 ;
      RECT 2.41 2.932 2.575 3.73 ;
      RECT 2.415 2.85 2.575 3.73 ;
      RECT 2.415 2.615 2.565 3.73 ;
      RECT 2.415 2.462 2.56 3.73 ;
      RECT 2.42 2.447 2.56 3.73 ;
      RECT 2.47 2.162 2.56 3.73 ;
      RECT 2.425 2.397 2.56 3.73 ;
      RECT 2.455 2.215 2.56 3.73 ;
      RECT 2.44 2.327 2.56 3.73 ;
      RECT 2.445 2.285 2.56 3.73 ;
      RECT 2.44 2.327 2.575 2.39 ;
      RECT 2.475 1.915 2.58 2.335 ;
      RECT 2.475 1.915 2.595 2.318 ;
      RECT 2.475 1.915 2.63 2.28 ;
      RECT 2.47 2.162 2.68 2.213 ;
      RECT 2.475 1.915 2.735 2.175 ;
      RECT 1.735 2.62 1.995 2.88 ;
      RECT 1.735 2.62 2.005 2.838 ;
      RECT 1.735 2.62 2.091 2.809 ;
      RECT 1.735 2.62 2.16 2.761 ;
      RECT 1.735 2.62 2.195 2.73 ;
      RECT 1.965 2.44 2.245 2.72 ;
      RECT 1.8 2.605 2.245 2.72 ;
      RECT 1.89 2.482 1.995 2.88 ;
      RECT 1.82 2.545 2.245 2.72 ;
    LAYER via1 ;
      RECT 75.83 1.195 75.98 1.345 ;
      RECT 73.46 6.74 73.61 6.89 ;
      RECT 73.445 2.065 73.595 2.215 ;
      RECT 72.655 2.45 72.805 2.6 ;
      RECT 72.655 6.37 72.805 6.52 ;
      RECT 71.625 2.805 71.775 2.955 ;
      RECT 71.62 5.96 71.77 6.11 ;
      RECT 71.065 2.805 71.215 2.955 ;
      RECT 69.295 2.35 69.445 2.5 ;
      RECT 68.275 3.055 68.425 3.205 ;
      RECT 68.045 2.475 68.195 2.625 ;
      RECT 67.7 3.075 67.85 3.225 ;
      RECT 67.46 2.095 67.61 2.245 ;
      RECT 67.15 3.425 67.3 3.575 ;
      RECT 67.01 2.03 67.16 2.18 ;
      RECT 66.375 2.115 66.525 2.265 ;
      RECT 66.265 2.755 66.415 2.905 ;
      RECT 65.94 3.315 66.09 3.465 ;
      RECT 65.77 2.305 65.92 2.455 ;
      RECT 65.415 3.32 65.565 3.47 ;
      RECT 65.355 2.535 65.505 2.685 ;
      RECT 64.99 3.525 65.14 3.675 ;
      RECT 64.83 2.36 64.98 2.51 ;
      RECT 64.265 2.435 64.415 2.585 ;
      RECT 63.87 2.385 64.02 2.535 ;
      RECT 63.57 1.97 63.72 2.12 ;
      RECT 63.485 3.525 63.635 3.675 ;
      RECT 62.83 2.675 62.98 2.825 ;
      RECT 60.57 1.195 60.72 1.345 ;
      RECT 58.2 6.74 58.35 6.89 ;
      RECT 58.185 2.065 58.335 2.215 ;
      RECT 57.395 2.45 57.545 2.6 ;
      RECT 57.395 6.37 57.545 6.52 ;
      RECT 56.365 2.805 56.515 2.955 ;
      RECT 56.36 5.96 56.51 6.11 ;
      RECT 55.805 2.805 55.955 2.955 ;
      RECT 54.035 2.35 54.185 2.5 ;
      RECT 53.015 3.055 53.165 3.205 ;
      RECT 52.785 2.475 52.935 2.625 ;
      RECT 52.44 3.075 52.59 3.225 ;
      RECT 52.2 2.095 52.35 2.245 ;
      RECT 51.89 3.425 52.04 3.575 ;
      RECT 51.75 2.03 51.9 2.18 ;
      RECT 51.115 2.115 51.265 2.265 ;
      RECT 51.005 2.755 51.155 2.905 ;
      RECT 50.68 3.315 50.83 3.465 ;
      RECT 50.51 2.305 50.66 2.455 ;
      RECT 50.155 3.32 50.305 3.47 ;
      RECT 50.095 2.535 50.245 2.685 ;
      RECT 49.73 3.525 49.88 3.675 ;
      RECT 49.57 2.36 49.72 2.51 ;
      RECT 49.005 2.435 49.155 2.585 ;
      RECT 48.61 2.385 48.76 2.535 ;
      RECT 48.31 1.97 48.46 2.12 ;
      RECT 48.225 3.525 48.375 3.675 ;
      RECT 47.57 2.675 47.72 2.825 ;
      RECT 45.31 1.195 45.46 1.345 ;
      RECT 42.94 6.74 43.09 6.89 ;
      RECT 42.925 2.065 43.075 2.215 ;
      RECT 42.135 2.45 42.285 2.6 ;
      RECT 42.135 6.37 42.285 6.52 ;
      RECT 41.105 2.805 41.255 2.955 ;
      RECT 41.1 5.96 41.25 6.11 ;
      RECT 40.545 2.805 40.695 2.955 ;
      RECT 38.775 2.35 38.925 2.5 ;
      RECT 37.755 3.055 37.905 3.205 ;
      RECT 37.525 2.475 37.675 2.625 ;
      RECT 37.18 3.075 37.33 3.225 ;
      RECT 36.94 2.095 37.09 2.245 ;
      RECT 36.63 3.425 36.78 3.575 ;
      RECT 36.49 2.03 36.64 2.18 ;
      RECT 35.855 2.115 36.005 2.265 ;
      RECT 35.745 2.755 35.895 2.905 ;
      RECT 35.42 3.315 35.57 3.465 ;
      RECT 35.25 2.305 35.4 2.455 ;
      RECT 34.895 3.32 35.045 3.47 ;
      RECT 34.835 2.535 34.985 2.685 ;
      RECT 34.47 3.525 34.62 3.675 ;
      RECT 34.31 2.36 34.46 2.51 ;
      RECT 33.745 2.435 33.895 2.585 ;
      RECT 33.35 2.385 33.5 2.535 ;
      RECT 33.05 1.97 33.2 2.12 ;
      RECT 32.965 3.525 33.115 3.675 ;
      RECT 32.31 2.675 32.46 2.825 ;
      RECT 30.05 1.195 30.2 1.345 ;
      RECT 27.68 6.74 27.83 6.89 ;
      RECT 27.665 2.065 27.815 2.215 ;
      RECT 26.875 2.45 27.025 2.6 ;
      RECT 26.875 6.37 27.025 6.52 ;
      RECT 25.845 2.805 25.995 2.955 ;
      RECT 25.84 5.96 25.99 6.11 ;
      RECT 25.285 2.805 25.435 2.955 ;
      RECT 23.515 2.35 23.665 2.5 ;
      RECT 22.495 3.055 22.645 3.205 ;
      RECT 22.265 2.475 22.415 2.625 ;
      RECT 21.92 3.075 22.07 3.225 ;
      RECT 21.68 2.095 21.83 2.245 ;
      RECT 21.37 3.425 21.52 3.575 ;
      RECT 21.23 2.03 21.38 2.18 ;
      RECT 20.595 2.115 20.745 2.265 ;
      RECT 20.485 2.755 20.635 2.905 ;
      RECT 20.16 3.315 20.31 3.465 ;
      RECT 19.99 2.305 20.14 2.455 ;
      RECT 19.635 3.32 19.785 3.47 ;
      RECT 19.575 2.535 19.725 2.685 ;
      RECT 19.21 3.525 19.36 3.675 ;
      RECT 19.05 2.36 19.2 2.51 ;
      RECT 18.485 2.435 18.635 2.585 ;
      RECT 18.09 2.385 18.24 2.535 ;
      RECT 17.79 1.97 17.94 2.12 ;
      RECT 17.705 3.525 17.855 3.675 ;
      RECT 17.05 2.675 17.2 2.825 ;
      RECT 14.79 1.195 14.94 1.345 ;
      RECT 12.42 6.74 12.57 6.89 ;
      RECT 12.405 2.065 12.555 2.215 ;
      RECT 11.615 2.45 11.765 2.6 ;
      RECT 11.615 6.37 11.765 6.52 ;
      RECT 10.585 2.805 10.735 2.955 ;
      RECT 10.58 5.96 10.73 6.11 ;
      RECT 10.025 2.805 10.175 2.955 ;
      RECT 8.255 2.35 8.405 2.5 ;
      RECT 7.235 3.055 7.385 3.205 ;
      RECT 7.005 2.475 7.155 2.625 ;
      RECT 6.66 3.075 6.81 3.225 ;
      RECT 6.42 2.095 6.57 2.245 ;
      RECT 6.11 3.425 6.26 3.575 ;
      RECT 5.97 2.03 6.12 2.18 ;
      RECT 5.335 2.115 5.485 2.265 ;
      RECT 5.225 2.755 5.375 2.905 ;
      RECT 4.9 3.315 5.05 3.465 ;
      RECT 4.73 2.305 4.88 2.455 ;
      RECT 4.375 3.32 4.525 3.47 ;
      RECT 4.315 2.535 4.465 2.685 ;
      RECT 3.95 3.525 4.1 3.675 ;
      RECT 3.79 2.36 3.94 2.51 ;
      RECT 3.225 2.435 3.375 2.585 ;
      RECT 2.83 2.385 2.98 2.535 ;
      RECT 2.53 1.97 2.68 2.12 ;
      RECT 2.445 3.525 2.595 3.675 ;
      RECT 1.79 2.675 1.94 2.825 ;
    LAYER met1 ;
      RECT 61.79 0 70.53 1.74 ;
      RECT 46.53 0 55.27 1.74 ;
      RECT 31.27 0 40.01 1.74 ;
      RECT 16.01 0 24.75 1.74 ;
      RECT 0.75 0 9.49 1.74 ;
      RECT 0 0 76.3 0.305 ;
      RECT 0 4.14 76.3 4.745 ;
      RECT 61.79 4.135 76.3 4.745 ;
      RECT 46.53 4.135 61.04 4.745 ;
      RECT 31.27 4.135 45.78 4.745 ;
      RECT 16.01 4.135 30.52 4.745 ;
      RECT 0.75 4.135 15.26 4.745 ;
      RECT 61.79 3.98 70.53 4.745 ;
      RECT 46.53 3.98 55.27 4.745 ;
      RECT 31.27 3.98 40.01 4.745 ;
      RECT 16.01 3.98 24.75 4.745 ;
      RECT 0.75 3.98 9.49 4.745 ;
      RECT 75.7 2.365 75.99 2.595 ;
      RECT 75.76 0.885 75.93 2.595 ;
      RECT 75.73 1.095 76.07 1.445 ;
      RECT 75.7 0.885 75.99 1.115 ;
      RECT 75.7 7.765 75.99 7.995 ;
      RECT 75.76 6.285 75.93 7.995 ;
      RECT 75.7 6.285 75.99 6.515 ;
      RECT 75.29 2.735 75.62 2.965 ;
      RECT 75.29 2.765 75.79 2.935 ;
      RECT 75.29 2.395 75.48 2.965 ;
      RECT 74.71 2.365 75 2.595 ;
      RECT 74.71 2.395 75.48 2.565 ;
      RECT 74.77 0.885 74.94 2.595 ;
      RECT 74.71 0.885 75 1.115 ;
      RECT 74.71 7.765 75 7.995 ;
      RECT 74.77 6.285 74.94 7.995 ;
      RECT 74.71 6.285 75 6.515 ;
      RECT 74.71 6.325 75.56 6.485 ;
      RECT 75.39 5.915 75.56 6.485 ;
      RECT 74.71 6.32 75.1 6.485 ;
      RECT 75.33 5.915 75.62 6.145 ;
      RECT 75.33 5.945 75.79 6.115 ;
      RECT 74.34 2.735 74.63 2.965 ;
      RECT 74.34 2.765 74.8 2.935 ;
      RECT 74.4 1.655 74.565 2.965 ;
      RECT 72.915 1.625 73.205 1.855 ;
      RECT 72.915 1.655 74.565 1.825 ;
      RECT 72.975 0.885 73.145 1.855 ;
      RECT 72.915 0.885 73.205 1.115 ;
      RECT 72.915 7.765 73.205 7.995 ;
      RECT 72.975 7.025 73.145 7.995 ;
      RECT 72.975 7.12 74.565 7.29 ;
      RECT 74.395 5.915 74.565 7.29 ;
      RECT 72.915 7.025 73.205 7.255 ;
      RECT 74.34 5.915 74.63 6.145 ;
      RECT 74.34 5.945 74.8 6.115 ;
      RECT 73.345 1.965 73.695 2.315 ;
      RECT 73.175 2.025 73.695 2.195 ;
      RECT 73.37 6.655 73.695 6.98 ;
      RECT 73.345 6.655 73.695 6.885 ;
      RECT 73.175 6.685 73.695 6.855 ;
      RECT 70.965 2.705 71.305 3.055 ;
      RECT 71.055 2.395 71.225 3.055 ;
      RECT 72.57 2.365 72.89 2.685 ;
      RECT 72.54 2.365 72.89 2.595 ;
      RECT 71.055 2.395 72.89 2.565 ;
      RECT 72.57 6.28 72.89 6.605 ;
      RECT 72.54 6.285 72.89 6.515 ;
      RECT 72.37 6.315 72.89 6.485 ;
      RECT 71.525 2.705 71.865 3.055 ;
      RECT 71.525 2.765 72.005 2.935 ;
      RECT 71.52 5.86 71.86 6.21 ;
      RECT 71.52 5.945 72.005 6.115 ;
      RECT 68.26 2.985 68.41 3.26 ;
      RECT 68.8 2.065 68.805 2.285 ;
      RECT 69.95 2.265 69.965 2.463 ;
      RECT 69.915 2.257 69.95 2.47 ;
      RECT 69.885 2.25 69.915 2.47 ;
      RECT 69.83 2.215 69.885 2.47 ;
      RECT 69.765 2.152 69.83 2.47 ;
      RECT 69.76 2.117 69.765 2.468 ;
      RECT 69.755 2.112 69.76 2.46 ;
      RECT 69.75 2.107 69.755 2.446 ;
      RECT 69.745 2.104 69.75 2.439 ;
      RECT 69.7 2.094 69.745 2.39 ;
      RECT 69.68 2.081 69.7 2.325 ;
      RECT 69.675 2.076 69.68 2.298 ;
      RECT 69.67 2.075 69.675 2.291 ;
      RECT 69.665 2.074 69.67 2.284 ;
      RECT 69.58 2.059 69.665 2.23 ;
      RECT 69.55 2.04 69.58 2.18 ;
      RECT 69.47 2.023 69.55 2.165 ;
      RECT 69.435 2.01 69.47 2.15 ;
      RECT 69.427 2.01 69.435 2.145 ;
      RECT 69.341 2.011 69.427 2.145 ;
      RECT 69.255 2.013 69.341 2.145 ;
      RECT 69.23 2.014 69.255 2.149 ;
      RECT 69.155 2.02 69.23 2.164 ;
      RECT 69.072 2.032 69.155 2.188 ;
      RECT 68.986 2.045 69.072 2.214 ;
      RECT 68.9 2.058 68.986 2.24 ;
      RECT 68.865 2.067 68.9 2.259 ;
      RECT 68.815 2.067 68.865 2.272 ;
      RECT 68.805 2.065 68.815 2.283 ;
      RECT 68.79 2.062 68.8 2.285 ;
      RECT 68.775 2.054 68.79 2.293 ;
      RECT 68.76 2.046 68.775 2.313 ;
      RECT 68.755 2.041 68.76 2.37 ;
      RECT 68.74 2.036 68.755 2.443 ;
      RECT 68.735 2.031 68.74 2.485 ;
      RECT 68.73 2.029 68.735 2.513 ;
      RECT 68.725 2.027 68.73 2.535 ;
      RECT 68.715 2.023 68.725 2.578 ;
      RECT 68.71 2.02 68.715 2.603 ;
      RECT 68.705 2.018 68.71 2.623 ;
      RECT 68.7 2.016 68.705 2.647 ;
      RECT 68.695 2.012 68.7 2.67 ;
      RECT 68.69 2.008 68.695 2.693 ;
      RECT 68.655 1.998 68.69 2.8 ;
      RECT 68.65 1.988 68.655 2.898 ;
      RECT 68.645 1.986 68.65 2.925 ;
      RECT 68.64 1.985 68.645 2.945 ;
      RECT 68.635 1.977 68.64 2.965 ;
      RECT 68.63 1.972 68.635 3 ;
      RECT 68.625 1.97 68.63 3.018 ;
      RECT 68.62 1.97 68.625 3.043 ;
      RECT 68.615 1.97 68.62 3.065 ;
      RECT 68.58 1.97 68.615 3.108 ;
      RECT 68.555 1.97 68.58 3.137 ;
      RECT 68.545 1.97 68.555 2.323 ;
      RECT 68.548 2.38 68.555 3.147 ;
      RECT 68.545 2.437 68.548 3.15 ;
      RECT 68.54 1.97 68.545 2.295 ;
      RECT 68.54 2.487 68.545 3.153 ;
      RECT 68.53 1.97 68.54 2.285 ;
      RECT 68.535 2.54 68.54 3.156 ;
      RECT 68.53 2.625 68.535 3.16 ;
      RECT 68.52 1.97 68.53 2.273 ;
      RECT 68.525 2.672 68.53 3.164 ;
      RECT 68.52 2.747 68.525 3.168 ;
      RECT 68.485 1.97 68.52 2.248 ;
      RECT 68.51 2.83 68.52 3.173 ;
      RECT 68.5 2.897 68.51 3.18 ;
      RECT 68.495 2.925 68.5 3.185 ;
      RECT 68.485 2.938 68.495 3.191 ;
      RECT 68.44 1.97 68.485 2.205 ;
      RECT 68.48 2.943 68.485 3.198 ;
      RECT 68.44 2.96 68.48 3.26 ;
      RECT 68.435 1.972 68.44 2.178 ;
      RECT 68.41 2.98 68.44 3.26 ;
      RECT 68.43 1.977 68.435 2.15 ;
      RECT 68.22 2.989 68.26 3.26 ;
      RECT 68.195 2.997 68.22 3.23 ;
      RECT 68.15 3.005 68.195 3.23 ;
      RECT 68.135 3.01 68.15 3.225 ;
      RECT 68.125 3.01 68.135 3.219 ;
      RECT 68.115 3.017 68.125 3.216 ;
      RECT 68.11 3.055 68.115 3.205 ;
      RECT 68.105 3.117 68.11 3.183 ;
      RECT 69.375 2.992 69.56 3.215 ;
      RECT 69.375 3.007 69.565 3.211 ;
      RECT 69.365 2.28 69.45 3.21 ;
      RECT 69.365 3.007 69.57 3.204 ;
      RECT 69.36 3.015 69.57 3.203 ;
      RECT 69.565 2.735 69.885 3.055 ;
      RECT 69.36 2.907 69.53 2.998 ;
      RECT 69.355 2.907 69.53 2.98 ;
      RECT 69.345 2.715 69.48 2.955 ;
      RECT 69.34 2.715 69.48 2.9 ;
      RECT 69.3 2.295 69.47 2.8 ;
      RECT 69.285 2.295 69.47 2.67 ;
      RECT 69.28 2.295 69.47 2.623 ;
      RECT 69.275 2.295 69.47 2.603 ;
      RECT 69.27 2.295 69.47 2.578 ;
      RECT 69.24 2.295 69.5 2.555 ;
      RECT 69.25 2.292 69.46 2.555 ;
      RECT 69.375 2.287 69.46 3.215 ;
      RECT 69.26 2.28 69.45 2.555 ;
      RECT 69.255 2.285 69.45 2.555 ;
      RECT 68.085 2.497 68.27 2.71 ;
      RECT 68.085 2.505 68.28 2.703 ;
      RECT 68.065 2.505 68.28 2.7 ;
      RECT 68.06 2.505 68.28 2.685 ;
      RECT 67.99 2.42 68.25 2.68 ;
      RECT 67.99 2.565 68.285 2.593 ;
      RECT 67.645 3.02 67.905 3.28 ;
      RECT 67.67 2.965 67.865 3.28 ;
      RECT 67.665 2.714 67.845 3.008 ;
      RECT 67.665 2.72 67.855 3.008 ;
      RECT 67.645 2.722 67.855 2.953 ;
      RECT 67.64 2.732 67.855 2.82 ;
      RECT 67.67 2.712 67.845 3.28 ;
      RECT 67.756 2.71 67.845 3.28 ;
      RECT 67.615 1.93 67.65 2.3 ;
      RECT 67.405 2.04 67.41 2.3 ;
      RECT 67.65 1.937 67.665 2.3 ;
      RECT 67.54 1.93 67.615 2.378 ;
      RECT 67.53 1.93 67.54 2.463 ;
      RECT 67.505 1.93 67.53 2.498 ;
      RECT 67.465 1.93 67.505 2.566 ;
      RECT 67.455 1.937 67.465 2.618 ;
      RECT 67.425 2.04 67.455 2.659 ;
      RECT 67.42 2.04 67.425 2.698 ;
      RECT 67.41 2.04 67.42 2.718 ;
      RECT 67.405 2.335 67.41 2.755 ;
      RECT 67.4 2.352 67.405 2.775 ;
      RECT 67.385 2.415 67.4 2.815 ;
      RECT 67.38 2.458 67.385 2.85 ;
      RECT 67.375 2.466 67.38 2.863 ;
      RECT 67.365 2.48 67.375 2.885 ;
      RECT 67.34 2.515 67.365 2.95 ;
      RECT 67.33 2.55 67.34 3.013 ;
      RECT 67.31 2.58 67.33 3.074 ;
      RECT 67.295 2.616 67.31 3.141 ;
      RECT 67.285 2.644 67.295 3.18 ;
      RECT 67.275 2.666 67.285 3.2 ;
      RECT 67.27 2.676 67.275 3.211 ;
      RECT 67.265 2.685 67.27 3.214 ;
      RECT 67.255 2.703 67.265 3.218 ;
      RECT 67.245 2.721 67.255 3.219 ;
      RECT 67.22 2.76 67.245 3.216 ;
      RECT 67.2 2.802 67.22 3.213 ;
      RECT 67.185 2.84 67.2 3.212 ;
      RECT 67.15 2.875 67.185 3.209 ;
      RECT 67.145 2.897 67.15 3.207 ;
      RECT 67.08 2.937 67.145 3.204 ;
      RECT 67.075 2.977 67.08 3.2 ;
      RECT 67.06 2.987 67.075 3.191 ;
      RECT 67.05 3.107 67.06 3.176 ;
      RECT 67.53 3.52 67.54 3.78 ;
      RECT 67.53 3.523 67.55 3.779 ;
      RECT 67.52 3.513 67.53 3.778 ;
      RECT 67.51 3.528 67.59 3.774 ;
      RECT 67.495 3.507 67.51 3.772 ;
      RECT 67.47 3.532 67.595 3.768 ;
      RECT 67.455 3.492 67.47 3.763 ;
      RECT 67.455 3.534 67.605 3.762 ;
      RECT 67.455 3.542 67.62 3.755 ;
      RECT 67.395 3.479 67.455 3.745 ;
      RECT 67.385 3.466 67.395 3.727 ;
      RECT 67.36 3.456 67.385 3.717 ;
      RECT 67.355 3.446 67.36 3.709 ;
      RECT 67.29 3.542 67.62 3.691 ;
      RECT 67.205 3.542 67.62 3.653 ;
      RECT 67.095 3.37 67.355 3.63 ;
      RECT 67.47 3.5 67.495 3.768 ;
      RECT 67.51 3.51 67.52 3.774 ;
      RECT 67.095 3.518 67.535 3.63 ;
      RECT 66.31 3.275 66.34 3.575 ;
      RECT 66.085 3.26 66.09 3.535 ;
      RECT 65.885 3.26 66.04 3.52 ;
      RECT 67.185 1.975 67.215 2.235 ;
      RECT 67.175 1.975 67.185 2.343 ;
      RECT 67.155 1.975 67.175 2.353 ;
      RECT 67.14 1.975 67.155 2.365 ;
      RECT 67.085 1.975 67.14 2.415 ;
      RECT 67.07 1.975 67.085 2.463 ;
      RECT 67.04 1.975 67.07 2.498 ;
      RECT 66.985 1.975 67.04 2.56 ;
      RECT 66.965 1.975 66.985 2.628 ;
      RECT 66.96 1.975 66.965 2.658 ;
      RECT 66.955 1.975 66.96 2.67 ;
      RECT 66.95 2.092 66.955 2.688 ;
      RECT 66.93 2.11 66.95 2.713 ;
      RECT 66.91 2.137 66.93 2.763 ;
      RECT 66.905 2.157 66.91 2.794 ;
      RECT 66.9 2.165 66.905 2.811 ;
      RECT 66.885 2.191 66.9 2.84 ;
      RECT 66.87 2.233 66.885 2.875 ;
      RECT 66.865 2.262 66.87 2.898 ;
      RECT 66.86 2.277 66.865 2.911 ;
      RECT 66.855 2.3 66.86 2.922 ;
      RECT 66.845 2.32 66.855 2.94 ;
      RECT 66.835 2.35 66.845 2.963 ;
      RECT 66.83 2.372 66.835 2.983 ;
      RECT 66.825 2.387 66.83 2.998 ;
      RECT 66.81 2.417 66.825 3.025 ;
      RECT 66.805 2.447 66.81 3.051 ;
      RECT 66.8 2.465 66.805 3.063 ;
      RECT 66.79 2.495 66.8 3.082 ;
      RECT 66.78 2.52 66.79 3.107 ;
      RECT 66.775 2.54 66.78 3.126 ;
      RECT 66.77 2.557 66.775 3.139 ;
      RECT 66.76 2.583 66.77 3.158 ;
      RECT 66.75 2.621 66.76 3.185 ;
      RECT 66.745 2.647 66.75 3.205 ;
      RECT 66.74 2.657 66.745 3.215 ;
      RECT 66.735 2.67 66.74 3.23 ;
      RECT 66.73 2.685 66.735 3.24 ;
      RECT 66.725 2.707 66.73 3.255 ;
      RECT 66.72 2.725 66.725 3.266 ;
      RECT 66.715 2.735 66.72 3.277 ;
      RECT 66.71 2.743 66.715 3.289 ;
      RECT 66.705 2.751 66.71 3.3 ;
      RECT 66.7 2.777 66.705 3.313 ;
      RECT 66.69 2.805 66.7 3.326 ;
      RECT 66.685 2.835 66.69 3.335 ;
      RECT 66.68 2.85 66.685 3.342 ;
      RECT 66.665 2.875 66.68 3.349 ;
      RECT 66.66 2.897 66.665 3.355 ;
      RECT 66.655 2.922 66.66 3.358 ;
      RECT 66.646 2.95 66.655 3.362 ;
      RECT 66.64 2.967 66.646 3.367 ;
      RECT 66.635 2.985 66.64 3.371 ;
      RECT 66.63 2.997 66.635 3.374 ;
      RECT 66.625 3.018 66.63 3.378 ;
      RECT 66.62 3.036 66.625 3.381 ;
      RECT 66.615 3.05 66.62 3.384 ;
      RECT 66.61 3.067 66.615 3.387 ;
      RECT 66.605 3.08 66.61 3.39 ;
      RECT 66.58 3.117 66.605 3.398 ;
      RECT 66.575 3.162 66.58 3.407 ;
      RECT 66.57 3.19 66.575 3.41 ;
      RECT 66.56 3.21 66.57 3.414 ;
      RECT 66.555 3.23 66.56 3.419 ;
      RECT 66.55 3.245 66.555 3.422 ;
      RECT 66.53 3.255 66.55 3.429 ;
      RECT 66.465 3.262 66.53 3.455 ;
      RECT 66.43 3.265 66.465 3.483 ;
      RECT 66.415 3.268 66.43 3.498 ;
      RECT 66.405 3.269 66.415 3.513 ;
      RECT 66.395 3.27 66.405 3.53 ;
      RECT 66.39 3.27 66.395 3.545 ;
      RECT 66.385 3.27 66.39 3.553 ;
      RECT 66.37 3.271 66.385 3.568 ;
      RECT 66.34 3.273 66.37 3.575 ;
      RECT 66.23 3.28 66.31 3.575 ;
      RECT 66.185 3.285 66.23 3.575 ;
      RECT 66.175 3.286 66.185 3.565 ;
      RECT 66.165 3.287 66.175 3.558 ;
      RECT 66.145 3.289 66.165 3.553 ;
      RECT 66.135 3.26 66.145 3.548 ;
      RECT 66.09 3.26 66.135 3.54 ;
      RECT 66.06 3.26 66.085 3.53 ;
      RECT 66.04 3.26 66.06 3.523 ;
      RECT 66.32 2.06 66.58 2.32 ;
      RECT 66.2 2.075 66.21 2.24 ;
      RECT 66.185 2.075 66.19 2.235 ;
      RECT 63.55 1.915 63.735 2.205 ;
      RECT 65.365 2.04 65.38 2.195 ;
      RECT 63.515 1.915 63.54 2.175 ;
      RECT 65.93 1.965 65.935 2.107 ;
      RECT 65.845 1.96 65.87 2.1 ;
      RECT 66.245 2.077 66.32 2.27 ;
      RECT 66.23 2.075 66.245 2.253 ;
      RECT 66.21 2.075 66.23 2.245 ;
      RECT 66.19 2.075 66.2 2.238 ;
      RECT 66.145 2.07 66.185 2.228 ;
      RECT 66.105 2.045 66.145 2.213 ;
      RECT 66.09 2.02 66.105 2.203 ;
      RECT 66.085 2.014 66.09 2.201 ;
      RECT 66.05 2.006 66.085 2.184 ;
      RECT 66.045 1.999 66.05 2.172 ;
      RECT 66.025 1.994 66.045 2.16 ;
      RECT 66.015 1.988 66.025 2.145 ;
      RECT 65.995 1.983 66.015 2.13 ;
      RECT 65.985 1.978 65.995 2.123 ;
      RECT 65.98 1.976 65.985 2.118 ;
      RECT 65.975 1.975 65.98 2.115 ;
      RECT 65.935 1.97 65.975 2.111 ;
      RECT 65.915 1.964 65.93 2.106 ;
      RECT 65.88 1.961 65.915 2.103 ;
      RECT 65.87 1.96 65.88 2.101 ;
      RECT 65.81 1.96 65.845 2.098 ;
      RECT 65.765 1.96 65.81 2.098 ;
      RECT 65.715 1.96 65.765 2.101 ;
      RECT 65.7 1.962 65.715 2.103 ;
      RECT 65.685 1.965 65.7 2.104 ;
      RECT 65.675 1.97 65.685 2.105 ;
      RECT 65.645 1.975 65.675 2.11 ;
      RECT 65.635 1.981 65.645 2.118 ;
      RECT 65.625 1.983 65.635 2.122 ;
      RECT 65.615 1.987 65.625 2.126 ;
      RECT 65.59 1.993 65.615 2.134 ;
      RECT 65.58 1.998 65.59 2.142 ;
      RECT 65.565 2.002 65.58 2.146 ;
      RECT 65.53 2.008 65.565 2.154 ;
      RECT 65.51 2.013 65.53 2.164 ;
      RECT 65.48 2.02 65.51 2.173 ;
      RECT 65.435 2.029 65.48 2.187 ;
      RECT 65.43 2.034 65.435 2.198 ;
      RECT 65.41 2.037 65.43 2.199 ;
      RECT 65.38 2.04 65.41 2.197 ;
      RECT 65.345 2.04 65.365 2.193 ;
      RECT 65.275 2.04 65.345 2.184 ;
      RECT 65.26 2.037 65.275 2.176 ;
      RECT 65.22 2.03 65.26 2.171 ;
      RECT 65.195 2.02 65.22 2.164 ;
      RECT 65.19 2.014 65.195 2.161 ;
      RECT 65.15 2.008 65.19 2.158 ;
      RECT 65.135 2.001 65.15 2.153 ;
      RECT 65.115 1.997 65.135 2.148 ;
      RECT 65.1 1.992 65.115 2.144 ;
      RECT 65.085 1.987 65.1 2.142 ;
      RECT 65.07 1.983 65.085 2.141 ;
      RECT 65.055 1.981 65.07 2.137 ;
      RECT 65.045 1.979 65.055 2.132 ;
      RECT 65.03 1.976 65.045 2.128 ;
      RECT 65.02 1.974 65.03 2.123 ;
      RECT 65 1.971 65.02 2.119 ;
      RECT 64.955 1.97 65 2.117 ;
      RECT 64.895 1.972 64.955 2.118 ;
      RECT 64.875 1.974 64.895 2.12 ;
      RECT 64.845 1.977 64.875 2.121 ;
      RECT 64.795 1.982 64.845 2.123 ;
      RECT 64.79 1.985 64.795 2.125 ;
      RECT 64.78 1.987 64.79 2.128 ;
      RECT 64.775 1.989 64.78 2.131 ;
      RECT 64.725 1.992 64.775 2.138 ;
      RECT 64.705 1.996 64.725 2.15 ;
      RECT 64.695 1.999 64.705 2.156 ;
      RECT 64.685 2 64.695 2.159 ;
      RECT 64.646 2.003 64.685 2.161 ;
      RECT 64.56 2.01 64.646 2.164 ;
      RECT 64.486 2.02 64.56 2.168 ;
      RECT 64.4 2.031 64.486 2.173 ;
      RECT 64.385 2.038 64.4 2.175 ;
      RECT 64.33 2.042 64.385 2.176 ;
      RECT 64.316 2.045 64.33 2.178 ;
      RECT 64.23 2.045 64.316 2.18 ;
      RECT 64.19 2.042 64.23 2.183 ;
      RECT 64.166 2.038 64.19 2.185 ;
      RECT 64.08 2.028 64.166 2.188 ;
      RECT 64.05 2.017 64.08 2.189 ;
      RECT 64.031 2.013 64.05 2.188 ;
      RECT 63.945 2.006 64.031 2.185 ;
      RECT 63.885 1.995 63.945 2.182 ;
      RECT 63.865 1.987 63.885 2.18 ;
      RECT 63.83 1.982 63.865 2.179 ;
      RECT 63.805 1.977 63.83 2.178 ;
      RECT 63.775 1.972 63.805 2.177 ;
      RECT 63.75 1.915 63.775 2.176 ;
      RECT 63.735 1.915 63.75 2.2 ;
      RECT 63.54 1.915 63.55 2.2 ;
      RECT 65.315 2.935 65.32 3.075 ;
      RECT 64.975 2.935 65.01 3.073 ;
      RECT 64.55 2.92 64.565 3.065 ;
      RECT 66.38 2.7 66.47 2.96 ;
      RECT 66.21 2.565 66.31 2.96 ;
      RECT 63.245 2.54 63.325 2.75 ;
      RECT 66.335 2.677 66.38 2.96 ;
      RECT 66.325 2.647 66.335 2.96 ;
      RECT 66.31 2.57 66.325 2.96 ;
      RECT 66.125 2.565 66.21 2.925 ;
      RECT 66.12 2.567 66.125 2.92 ;
      RECT 66.115 2.572 66.12 2.92 ;
      RECT 66.08 2.672 66.115 2.92 ;
      RECT 66.07 2.7 66.08 2.92 ;
      RECT 66.06 2.715 66.07 2.92 ;
      RECT 66.05 2.727 66.06 2.92 ;
      RECT 66.045 2.737 66.05 2.92 ;
      RECT 66.03 2.747 66.045 2.922 ;
      RECT 66.025 2.762 66.03 2.924 ;
      RECT 66.01 2.775 66.025 2.926 ;
      RECT 66.005 2.79 66.01 2.929 ;
      RECT 65.985 2.8 66.005 2.933 ;
      RECT 65.97 2.81 65.985 2.936 ;
      RECT 65.935 2.817 65.97 2.941 ;
      RECT 65.891 2.824 65.935 2.949 ;
      RECT 65.805 2.836 65.891 2.962 ;
      RECT 65.78 2.847 65.805 2.973 ;
      RECT 65.75 2.852 65.78 2.978 ;
      RECT 65.715 2.857 65.75 2.986 ;
      RECT 65.685 2.862 65.715 2.993 ;
      RECT 65.66 2.867 65.685 2.998 ;
      RECT 65.595 2.874 65.66 3.007 ;
      RECT 65.525 2.887 65.595 3.023 ;
      RECT 65.495 2.897 65.525 3.035 ;
      RECT 65.47 2.902 65.495 3.042 ;
      RECT 65.415 2.909 65.47 3.05 ;
      RECT 65.41 2.916 65.415 3.055 ;
      RECT 65.405 2.918 65.41 3.056 ;
      RECT 65.39 2.92 65.405 3.058 ;
      RECT 65.385 2.92 65.39 3.061 ;
      RECT 65.32 2.927 65.385 3.068 ;
      RECT 65.285 2.937 65.315 3.078 ;
      RECT 65.268 2.94 65.285 3.08 ;
      RECT 65.182 2.939 65.268 3.079 ;
      RECT 65.096 2.937 65.182 3.076 ;
      RECT 65.01 2.936 65.096 3.074 ;
      RECT 64.909 2.934 64.975 3.073 ;
      RECT 64.823 2.931 64.909 3.071 ;
      RECT 64.737 2.927 64.823 3.069 ;
      RECT 64.651 2.924 64.737 3.068 ;
      RECT 64.565 2.921 64.651 3.066 ;
      RECT 64.465 2.92 64.55 3.063 ;
      RECT 64.415 2.918 64.465 3.061 ;
      RECT 64.395 2.915 64.415 3.059 ;
      RECT 64.375 2.913 64.395 3.056 ;
      RECT 64.35 2.909 64.375 3.053 ;
      RECT 64.305 2.903 64.35 3.048 ;
      RECT 64.265 2.897 64.305 3.04 ;
      RECT 64.24 2.892 64.265 3.033 ;
      RECT 64.185 2.885 64.24 3.025 ;
      RECT 64.161 2.878 64.185 3.018 ;
      RECT 64.075 2.869 64.161 3.008 ;
      RECT 64.045 2.861 64.075 2.998 ;
      RECT 64.015 2.857 64.045 2.993 ;
      RECT 64.01 2.854 64.015 2.99 ;
      RECT 64.005 2.853 64.01 2.99 ;
      RECT 63.93 2.846 64.005 2.983 ;
      RECT 63.891 2.837 63.93 2.972 ;
      RECT 63.805 2.827 63.891 2.96 ;
      RECT 63.765 2.817 63.805 2.948 ;
      RECT 63.726 2.812 63.765 2.941 ;
      RECT 63.64 2.802 63.726 2.93 ;
      RECT 63.6 2.79 63.64 2.919 ;
      RECT 63.565 2.775 63.6 2.912 ;
      RECT 63.555 2.765 63.565 2.909 ;
      RECT 63.535 2.75 63.555 2.907 ;
      RECT 63.505 2.72 63.535 2.903 ;
      RECT 63.495 2.7 63.505 2.898 ;
      RECT 63.49 2.692 63.495 2.895 ;
      RECT 63.485 2.685 63.49 2.893 ;
      RECT 63.47 2.672 63.485 2.886 ;
      RECT 63.465 2.662 63.47 2.878 ;
      RECT 63.46 2.655 63.465 2.873 ;
      RECT 63.455 2.65 63.46 2.869 ;
      RECT 63.44 2.637 63.455 2.861 ;
      RECT 63.435 2.547 63.44 2.85 ;
      RECT 63.43 2.542 63.435 2.843 ;
      RECT 63.355 2.54 63.43 2.803 ;
      RECT 63.325 2.54 63.355 2.758 ;
      RECT 63.23 2.545 63.245 2.745 ;
      RECT 65.715 2.25 65.975 2.51 ;
      RECT 65.7 2.238 65.88 2.475 ;
      RECT 65.695 2.239 65.88 2.473 ;
      RECT 65.68 2.243 65.89 2.463 ;
      RECT 65.675 2.248 65.895 2.433 ;
      RECT 65.68 2.245 65.895 2.463 ;
      RECT 65.695 2.24 65.89 2.473 ;
      RECT 65.715 2.237 65.88 2.51 ;
      RECT 65.715 2.236 65.87 2.51 ;
      RECT 65.74 2.235 65.87 2.51 ;
      RECT 65.3 2.48 65.56 2.74 ;
      RECT 65.175 2.525 65.56 2.735 ;
      RECT 65.165 2.53 65.56 2.73 ;
      RECT 65.18 3.47 65.195 3.78 ;
      RECT 63.775 3.24 63.785 3.37 ;
      RECT 63.555 3.235 63.66 3.37 ;
      RECT 63.47 3.24 63.52 3.37 ;
      RECT 62.02 1.975 62.025 3.08 ;
      RECT 65.275 3.562 65.28 3.698 ;
      RECT 65.27 3.557 65.275 3.758 ;
      RECT 65.265 3.555 65.27 3.771 ;
      RECT 65.25 3.552 65.265 3.773 ;
      RECT 65.245 3.547 65.25 3.775 ;
      RECT 65.24 3.543 65.245 3.778 ;
      RECT 65.225 3.538 65.24 3.78 ;
      RECT 65.195 3.53 65.225 3.78 ;
      RECT 65.156 3.47 65.18 3.78 ;
      RECT 65.07 3.47 65.156 3.777 ;
      RECT 65.04 3.47 65.07 3.77 ;
      RECT 65.015 3.47 65.04 3.763 ;
      RECT 64.99 3.47 65.015 3.755 ;
      RECT 64.975 3.47 64.99 3.748 ;
      RECT 64.95 3.47 64.975 3.74 ;
      RECT 64.935 3.47 64.95 3.733 ;
      RECT 64.895 3.48 64.935 3.722 ;
      RECT 64.885 3.475 64.895 3.712 ;
      RECT 64.881 3.474 64.885 3.709 ;
      RECT 64.795 3.466 64.881 3.692 ;
      RECT 64.762 3.455 64.795 3.669 ;
      RECT 64.676 3.444 64.762 3.647 ;
      RECT 64.59 3.428 64.676 3.616 ;
      RECT 64.52 3.413 64.59 3.588 ;
      RECT 64.51 3.406 64.52 3.575 ;
      RECT 64.48 3.403 64.51 3.565 ;
      RECT 64.455 3.399 64.48 3.558 ;
      RECT 64.44 3.396 64.455 3.553 ;
      RECT 64.435 3.395 64.44 3.548 ;
      RECT 64.405 3.39 64.435 3.541 ;
      RECT 64.4 3.385 64.405 3.536 ;
      RECT 64.385 3.382 64.4 3.531 ;
      RECT 64.38 3.377 64.385 3.526 ;
      RECT 64.36 3.372 64.38 3.523 ;
      RECT 64.345 3.367 64.36 3.515 ;
      RECT 64.33 3.361 64.345 3.51 ;
      RECT 64.3 3.352 64.33 3.503 ;
      RECT 64.295 3.345 64.3 3.495 ;
      RECT 64.29 3.343 64.295 3.493 ;
      RECT 64.285 3.342 64.29 3.49 ;
      RECT 64.245 3.335 64.285 3.483 ;
      RECT 64.231 3.325 64.245 3.473 ;
      RECT 64.18 3.314 64.231 3.461 ;
      RECT 64.155 3.3 64.18 3.447 ;
      RECT 64.13 3.289 64.155 3.439 ;
      RECT 64.11 3.278 64.13 3.433 ;
      RECT 64.1 3.272 64.11 3.428 ;
      RECT 64.095 3.27 64.1 3.424 ;
      RECT 64.075 3.265 64.095 3.419 ;
      RECT 64.045 3.255 64.075 3.409 ;
      RECT 64.04 3.247 64.045 3.402 ;
      RECT 64.025 3.245 64.04 3.398 ;
      RECT 64.005 3.245 64.025 3.393 ;
      RECT 64 3.244 64.005 3.391 ;
      RECT 63.995 3.244 64 3.388 ;
      RECT 63.955 3.243 63.995 3.383 ;
      RECT 63.93 3.242 63.955 3.378 ;
      RECT 63.87 3.241 63.93 3.375 ;
      RECT 63.785 3.24 63.87 3.373 ;
      RECT 63.746 3.239 63.775 3.37 ;
      RECT 63.66 3.237 63.746 3.37 ;
      RECT 63.52 3.237 63.555 3.37 ;
      RECT 63.43 3.241 63.47 3.373 ;
      RECT 63.415 3.244 63.43 3.38 ;
      RECT 63.405 3.245 63.415 3.387 ;
      RECT 63.38 3.248 63.405 3.392 ;
      RECT 63.375 3.25 63.38 3.395 ;
      RECT 63.325 3.252 63.375 3.396 ;
      RECT 63.286 3.256 63.325 3.398 ;
      RECT 63.2 3.258 63.286 3.401 ;
      RECT 63.182 3.26 63.2 3.403 ;
      RECT 63.096 3.263 63.182 3.405 ;
      RECT 63.01 3.267 63.096 3.408 ;
      RECT 62.973 3.271 63.01 3.411 ;
      RECT 62.887 3.274 62.973 3.414 ;
      RECT 62.801 3.278 62.887 3.417 ;
      RECT 62.715 3.283 62.801 3.421 ;
      RECT 62.695 3.285 62.715 3.424 ;
      RECT 62.675 3.284 62.695 3.425 ;
      RECT 62.626 3.281 62.675 3.426 ;
      RECT 62.54 3.276 62.626 3.429 ;
      RECT 62.49 3.271 62.54 3.431 ;
      RECT 62.466 3.269 62.49 3.432 ;
      RECT 62.38 3.264 62.466 3.434 ;
      RECT 62.355 3.26 62.38 3.433 ;
      RECT 62.345 3.257 62.355 3.431 ;
      RECT 62.335 3.25 62.345 3.428 ;
      RECT 62.33 3.23 62.335 3.423 ;
      RECT 62.32 3.2 62.33 3.418 ;
      RECT 62.305 3.07 62.32 3.409 ;
      RECT 62.3 3.062 62.305 3.402 ;
      RECT 62.28 3.055 62.3 3.394 ;
      RECT 62.275 3.037 62.28 3.386 ;
      RECT 62.265 3.017 62.275 3.381 ;
      RECT 62.26 2.99 62.265 3.377 ;
      RECT 62.255 2.967 62.26 3.374 ;
      RECT 62.235 2.925 62.255 3.366 ;
      RECT 62.2 2.84 62.235 3.35 ;
      RECT 62.195 2.772 62.2 3.338 ;
      RECT 62.18 2.742 62.195 3.332 ;
      RECT 62.175 1.987 62.18 2.233 ;
      RECT 62.165 2.712 62.18 3.323 ;
      RECT 62.17 1.982 62.175 2.265 ;
      RECT 62.165 1.977 62.17 2.308 ;
      RECT 62.16 1.975 62.165 2.343 ;
      RECT 62.145 2.675 62.165 3.313 ;
      RECT 62.155 1.975 62.16 2.38 ;
      RECT 62.14 1.975 62.155 2.478 ;
      RECT 62.14 2.648 62.145 3.306 ;
      RECT 62.135 1.975 62.14 2.553 ;
      RECT 62.135 2.636 62.14 3.303 ;
      RECT 62.13 1.975 62.135 2.585 ;
      RECT 62.13 2.615 62.135 3.3 ;
      RECT 62.125 1.975 62.13 3.297 ;
      RECT 62.09 1.975 62.125 3.283 ;
      RECT 62.075 1.975 62.09 3.265 ;
      RECT 62.055 1.975 62.075 3.255 ;
      RECT 62.03 1.975 62.055 3.238 ;
      RECT 62.025 1.975 62.03 3.188 ;
      RECT 62.015 1.975 62.02 3.018 ;
      RECT 62.01 1.975 62.015 2.925 ;
      RECT 62.005 1.975 62.01 2.838 ;
      RECT 62 1.975 62.005 2.77 ;
      RECT 61.995 1.975 62 2.713 ;
      RECT 61.985 1.975 61.995 2.608 ;
      RECT 61.98 1.975 61.985 2.48 ;
      RECT 61.975 1.975 61.98 2.398 ;
      RECT 61.97 1.977 61.975 2.315 ;
      RECT 61.965 1.982 61.97 2.248 ;
      RECT 61.96 1.987 61.965 2.175 ;
      RECT 64.775 2.305 65.035 2.565 ;
      RECT 64.795 2.272 65.005 2.565 ;
      RECT 64.795 2.27 64.995 2.565 ;
      RECT 64.805 2.257 64.995 2.565 ;
      RECT 64.805 2.255 64.92 2.565 ;
      RECT 64.28 2.38 64.455 2.66 ;
      RECT 64.275 2.38 64.455 2.658 ;
      RECT 64.275 2.38 64.47 2.655 ;
      RECT 64.265 2.38 64.47 2.653 ;
      RECT 64.21 2.38 64.47 2.64 ;
      RECT 64.21 2.455 64.475 2.618 ;
      RECT 63.755 2.392 63.775 2.635 ;
      RECT 63.755 2.392 63.815 2.634 ;
      RECT 63.75 2.394 63.815 2.633 ;
      RECT 63.75 2.394 63.901 2.632 ;
      RECT 63.75 2.394 63.97 2.631 ;
      RECT 63.75 2.394 63.99 2.623 ;
      RECT 63.73 2.397 63.99 2.621 ;
      RECT 63.715 2.407 63.99 2.606 ;
      RECT 63.715 2.407 64.005 2.605 ;
      RECT 63.71 2.416 64.005 2.597 ;
      RECT 63.71 2.416 64.01 2.593 ;
      RECT 63.815 2.33 64.075 2.59 ;
      RECT 63.705 2.418 64.075 2.475 ;
      RECT 63.775 2.385 64.075 2.59 ;
      RECT 63.74 3.578 63.745 3.785 ;
      RECT 63.69 3.572 63.74 3.784 ;
      RECT 63.657 3.586 63.75 3.783 ;
      RECT 63.571 3.586 63.75 3.782 ;
      RECT 63.485 3.586 63.75 3.781 ;
      RECT 63.485 3.685 63.755 3.778 ;
      RECT 63.48 3.685 63.755 3.773 ;
      RECT 63.475 3.685 63.755 3.755 ;
      RECT 63.47 3.685 63.755 3.738 ;
      RECT 63.43 3.47 63.69 3.73 ;
      RECT 62.89 2.62 62.976 3.034 ;
      RECT 62.89 2.62 63.015 3.031 ;
      RECT 62.89 2.62 63.035 3.021 ;
      RECT 62.845 2.62 63.035 3.018 ;
      RECT 62.845 2.772 63.045 3.008 ;
      RECT 62.845 2.793 63.05 3.002 ;
      RECT 62.845 2.811 63.055 2.998 ;
      RECT 62.845 2.831 63.065 2.993 ;
      RECT 62.82 2.831 63.065 2.99 ;
      RECT 62.81 2.831 63.065 2.968 ;
      RECT 62.81 2.847 63.07 2.938 ;
      RECT 62.775 2.62 63.035 2.925 ;
      RECT 62.775 2.859 63.075 2.88 ;
      RECT 60.44 2.365 60.73 2.595 ;
      RECT 60.5 0.885 60.67 2.595 ;
      RECT 60.47 1.095 60.81 1.445 ;
      RECT 60.44 0.885 60.73 1.115 ;
      RECT 60.44 7.765 60.73 7.995 ;
      RECT 60.5 6.285 60.67 7.995 ;
      RECT 60.44 6.285 60.73 6.515 ;
      RECT 60.03 2.735 60.36 2.965 ;
      RECT 60.03 2.765 60.53 2.935 ;
      RECT 60.03 2.395 60.22 2.965 ;
      RECT 59.45 2.365 59.74 2.595 ;
      RECT 59.45 2.395 60.22 2.565 ;
      RECT 59.51 0.885 59.68 2.595 ;
      RECT 59.45 0.885 59.74 1.115 ;
      RECT 59.45 7.765 59.74 7.995 ;
      RECT 59.51 6.285 59.68 7.995 ;
      RECT 59.45 6.285 59.74 6.515 ;
      RECT 59.45 6.325 60.3 6.485 ;
      RECT 60.13 5.915 60.3 6.485 ;
      RECT 59.45 6.32 59.84 6.485 ;
      RECT 60.07 5.915 60.36 6.145 ;
      RECT 60.07 5.945 60.53 6.115 ;
      RECT 59.08 2.735 59.37 2.965 ;
      RECT 59.08 2.765 59.54 2.935 ;
      RECT 59.14 1.655 59.305 2.965 ;
      RECT 57.655 1.625 57.945 1.855 ;
      RECT 57.655 1.655 59.305 1.825 ;
      RECT 57.715 0.885 57.885 1.855 ;
      RECT 57.655 0.885 57.945 1.115 ;
      RECT 57.655 7.765 57.945 7.995 ;
      RECT 57.715 7.025 57.885 7.995 ;
      RECT 57.715 7.12 59.305 7.29 ;
      RECT 59.135 5.915 59.305 7.29 ;
      RECT 57.655 7.025 57.945 7.255 ;
      RECT 59.08 5.915 59.37 6.145 ;
      RECT 59.08 5.945 59.54 6.115 ;
      RECT 58.085 1.965 58.435 2.315 ;
      RECT 57.915 2.025 58.435 2.195 ;
      RECT 58.11 6.655 58.435 6.98 ;
      RECT 58.085 6.655 58.435 6.885 ;
      RECT 57.915 6.685 58.435 6.855 ;
      RECT 55.705 2.705 56.045 3.055 ;
      RECT 55.795 2.395 55.965 3.055 ;
      RECT 57.31 2.365 57.63 2.685 ;
      RECT 57.28 2.365 57.63 2.595 ;
      RECT 55.795 2.395 57.63 2.565 ;
      RECT 57.31 6.28 57.63 6.605 ;
      RECT 57.28 6.285 57.63 6.515 ;
      RECT 57.11 6.315 57.63 6.485 ;
      RECT 56.265 2.705 56.605 3.055 ;
      RECT 56.265 2.765 56.745 2.935 ;
      RECT 56.26 5.86 56.6 6.21 ;
      RECT 56.26 5.945 56.745 6.115 ;
      RECT 53 2.985 53.15 3.26 ;
      RECT 53.54 2.065 53.545 2.285 ;
      RECT 54.69 2.265 54.705 2.463 ;
      RECT 54.655 2.257 54.69 2.47 ;
      RECT 54.625 2.25 54.655 2.47 ;
      RECT 54.57 2.215 54.625 2.47 ;
      RECT 54.505 2.152 54.57 2.47 ;
      RECT 54.5 2.117 54.505 2.468 ;
      RECT 54.495 2.112 54.5 2.46 ;
      RECT 54.49 2.107 54.495 2.446 ;
      RECT 54.485 2.104 54.49 2.439 ;
      RECT 54.44 2.094 54.485 2.39 ;
      RECT 54.42 2.081 54.44 2.325 ;
      RECT 54.415 2.076 54.42 2.298 ;
      RECT 54.41 2.075 54.415 2.291 ;
      RECT 54.405 2.074 54.41 2.284 ;
      RECT 54.32 2.059 54.405 2.23 ;
      RECT 54.29 2.04 54.32 2.18 ;
      RECT 54.21 2.023 54.29 2.165 ;
      RECT 54.175 2.01 54.21 2.15 ;
      RECT 54.167 2.01 54.175 2.145 ;
      RECT 54.081 2.011 54.167 2.145 ;
      RECT 53.995 2.013 54.081 2.145 ;
      RECT 53.97 2.014 53.995 2.149 ;
      RECT 53.895 2.02 53.97 2.164 ;
      RECT 53.812 2.032 53.895 2.188 ;
      RECT 53.726 2.045 53.812 2.214 ;
      RECT 53.64 2.058 53.726 2.24 ;
      RECT 53.605 2.067 53.64 2.259 ;
      RECT 53.555 2.067 53.605 2.272 ;
      RECT 53.545 2.065 53.555 2.283 ;
      RECT 53.53 2.062 53.54 2.285 ;
      RECT 53.515 2.054 53.53 2.293 ;
      RECT 53.5 2.046 53.515 2.313 ;
      RECT 53.495 2.041 53.5 2.37 ;
      RECT 53.48 2.036 53.495 2.443 ;
      RECT 53.475 2.031 53.48 2.485 ;
      RECT 53.47 2.029 53.475 2.513 ;
      RECT 53.465 2.027 53.47 2.535 ;
      RECT 53.455 2.023 53.465 2.578 ;
      RECT 53.45 2.02 53.455 2.603 ;
      RECT 53.445 2.018 53.45 2.623 ;
      RECT 53.44 2.016 53.445 2.647 ;
      RECT 53.435 2.012 53.44 2.67 ;
      RECT 53.43 2.008 53.435 2.693 ;
      RECT 53.395 1.998 53.43 2.8 ;
      RECT 53.39 1.988 53.395 2.898 ;
      RECT 53.385 1.986 53.39 2.925 ;
      RECT 53.38 1.985 53.385 2.945 ;
      RECT 53.375 1.977 53.38 2.965 ;
      RECT 53.37 1.972 53.375 3 ;
      RECT 53.365 1.97 53.37 3.018 ;
      RECT 53.36 1.97 53.365 3.043 ;
      RECT 53.355 1.97 53.36 3.065 ;
      RECT 53.32 1.97 53.355 3.108 ;
      RECT 53.295 1.97 53.32 3.137 ;
      RECT 53.285 1.97 53.295 2.323 ;
      RECT 53.288 2.38 53.295 3.147 ;
      RECT 53.285 2.437 53.288 3.15 ;
      RECT 53.28 1.97 53.285 2.295 ;
      RECT 53.28 2.487 53.285 3.153 ;
      RECT 53.27 1.97 53.28 2.285 ;
      RECT 53.275 2.54 53.28 3.156 ;
      RECT 53.27 2.625 53.275 3.16 ;
      RECT 53.26 1.97 53.27 2.273 ;
      RECT 53.265 2.672 53.27 3.164 ;
      RECT 53.26 2.747 53.265 3.168 ;
      RECT 53.225 1.97 53.26 2.248 ;
      RECT 53.25 2.83 53.26 3.173 ;
      RECT 53.24 2.897 53.25 3.18 ;
      RECT 53.235 2.925 53.24 3.185 ;
      RECT 53.225 2.938 53.235 3.191 ;
      RECT 53.18 1.97 53.225 2.205 ;
      RECT 53.22 2.943 53.225 3.198 ;
      RECT 53.18 2.96 53.22 3.26 ;
      RECT 53.175 1.972 53.18 2.178 ;
      RECT 53.15 2.98 53.18 3.26 ;
      RECT 53.17 1.977 53.175 2.15 ;
      RECT 52.96 2.989 53 3.26 ;
      RECT 52.935 2.997 52.96 3.23 ;
      RECT 52.89 3.005 52.935 3.23 ;
      RECT 52.875 3.01 52.89 3.225 ;
      RECT 52.865 3.01 52.875 3.219 ;
      RECT 52.855 3.017 52.865 3.216 ;
      RECT 52.85 3.055 52.855 3.205 ;
      RECT 52.845 3.117 52.85 3.183 ;
      RECT 54.115 2.992 54.3 3.215 ;
      RECT 54.115 3.007 54.305 3.211 ;
      RECT 54.105 2.28 54.19 3.21 ;
      RECT 54.105 3.007 54.31 3.204 ;
      RECT 54.1 3.015 54.31 3.203 ;
      RECT 54.305 2.735 54.625 3.055 ;
      RECT 54.1 2.907 54.27 2.998 ;
      RECT 54.095 2.907 54.27 2.98 ;
      RECT 54.085 2.715 54.22 2.955 ;
      RECT 54.08 2.715 54.22 2.9 ;
      RECT 54.04 2.295 54.21 2.8 ;
      RECT 54.025 2.295 54.21 2.67 ;
      RECT 54.02 2.295 54.21 2.623 ;
      RECT 54.015 2.295 54.21 2.603 ;
      RECT 54.01 2.295 54.21 2.578 ;
      RECT 53.98 2.295 54.24 2.555 ;
      RECT 53.99 2.292 54.2 2.555 ;
      RECT 54.115 2.287 54.2 3.215 ;
      RECT 54 2.28 54.19 2.555 ;
      RECT 53.995 2.285 54.19 2.555 ;
      RECT 52.825 2.497 53.01 2.71 ;
      RECT 52.825 2.505 53.02 2.703 ;
      RECT 52.805 2.505 53.02 2.7 ;
      RECT 52.8 2.505 53.02 2.685 ;
      RECT 52.73 2.42 52.99 2.68 ;
      RECT 52.73 2.565 53.025 2.593 ;
      RECT 52.385 3.02 52.645 3.28 ;
      RECT 52.41 2.965 52.605 3.28 ;
      RECT 52.405 2.714 52.585 3.008 ;
      RECT 52.405 2.72 52.595 3.008 ;
      RECT 52.385 2.722 52.595 2.953 ;
      RECT 52.38 2.732 52.595 2.82 ;
      RECT 52.41 2.712 52.585 3.28 ;
      RECT 52.496 2.71 52.585 3.28 ;
      RECT 52.355 1.93 52.39 2.3 ;
      RECT 52.145 2.04 52.15 2.3 ;
      RECT 52.39 1.937 52.405 2.3 ;
      RECT 52.28 1.93 52.355 2.378 ;
      RECT 52.27 1.93 52.28 2.463 ;
      RECT 52.245 1.93 52.27 2.498 ;
      RECT 52.205 1.93 52.245 2.566 ;
      RECT 52.195 1.937 52.205 2.618 ;
      RECT 52.165 2.04 52.195 2.659 ;
      RECT 52.16 2.04 52.165 2.698 ;
      RECT 52.15 2.04 52.16 2.718 ;
      RECT 52.145 2.335 52.15 2.755 ;
      RECT 52.14 2.352 52.145 2.775 ;
      RECT 52.125 2.415 52.14 2.815 ;
      RECT 52.12 2.458 52.125 2.85 ;
      RECT 52.115 2.466 52.12 2.863 ;
      RECT 52.105 2.48 52.115 2.885 ;
      RECT 52.08 2.515 52.105 2.95 ;
      RECT 52.07 2.55 52.08 3.013 ;
      RECT 52.05 2.58 52.07 3.074 ;
      RECT 52.035 2.616 52.05 3.141 ;
      RECT 52.025 2.644 52.035 3.18 ;
      RECT 52.015 2.666 52.025 3.2 ;
      RECT 52.01 2.676 52.015 3.211 ;
      RECT 52.005 2.685 52.01 3.214 ;
      RECT 51.995 2.703 52.005 3.218 ;
      RECT 51.985 2.721 51.995 3.219 ;
      RECT 51.96 2.76 51.985 3.216 ;
      RECT 51.94 2.802 51.96 3.213 ;
      RECT 51.925 2.84 51.94 3.212 ;
      RECT 51.89 2.875 51.925 3.209 ;
      RECT 51.885 2.897 51.89 3.207 ;
      RECT 51.82 2.937 51.885 3.204 ;
      RECT 51.815 2.977 51.82 3.2 ;
      RECT 51.8 2.987 51.815 3.191 ;
      RECT 51.79 3.107 51.8 3.176 ;
      RECT 52.27 3.52 52.28 3.78 ;
      RECT 52.27 3.523 52.29 3.779 ;
      RECT 52.26 3.513 52.27 3.778 ;
      RECT 52.25 3.528 52.33 3.774 ;
      RECT 52.235 3.507 52.25 3.772 ;
      RECT 52.21 3.532 52.335 3.768 ;
      RECT 52.195 3.492 52.21 3.763 ;
      RECT 52.195 3.534 52.345 3.762 ;
      RECT 52.195 3.542 52.36 3.755 ;
      RECT 52.135 3.479 52.195 3.745 ;
      RECT 52.125 3.466 52.135 3.727 ;
      RECT 52.1 3.456 52.125 3.717 ;
      RECT 52.095 3.446 52.1 3.709 ;
      RECT 52.03 3.542 52.36 3.691 ;
      RECT 51.945 3.542 52.36 3.653 ;
      RECT 51.835 3.37 52.095 3.63 ;
      RECT 52.21 3.5 52.235 3.768 ;
      RECT 52.25 3.51 52.26 3.774 ;
      RECT 51.835 3.518 52.275 3.63 ;
      RECT 51.05 3.275 51.08 3.575 ;
      RECT 50.825 3.26 50.83 3.535 ;
      RECT 50.625 3.26 50.78 3.52 ;
      RECT 51.925 1.975 51.955 2.235 ;
      RECT 51.915 1.975 51.925 2.343 ;
      RECT 51.895 1.975 51.915 2.353 ;
      RECT 51.88 1.975 51.895 2.365 ;
      RECT 51.825 1.975 51.88 2.415 ;
      RECT 51.81 1.975 51.825 2.463 ;
      RECT 51.78 1.975 51.81 2.498 ;
      RECT 51.725 1.975 51.78 2.56 ;
      RECT 51.705 1.975 51.725 2.628 ;
      RECT 51.7 1.975 51.705 2.658 ;
      RECT 51.695 1.975 51.7 2.67 ;
      RECT 51.69 2.092 51.695 2.688 ;
      RECT 51.67 2.11 51.69 2.713 ;
      RECT 51.65 2.137 51.67 2.763 ;
      RECT 51.645 2.157 51.65 2.794 ;
      RECT 51.64 2.165 51.645 2.811 ;
      RECT 51.625 2.191 51.64 2.84 ;
      RECT 51.61 2.233 51.625 2.875 ;
      RECT 51.605 2.262 51.61 2.898 ;
      RECT 51.6 2.277 51.605 2.911 ;
      RECT 51.595 2.3 51.6 2.922 ;
      RECT 51.585 2.32 51.595 2.94 ;
      RECT 51.575 2.35 51.585 2.963 ;
      RECT 51.57 2.372 51.575 2.983 ;
      RECT 51.565 2.387 51.57 2.998 ;
      RECT 51.55 2.417 51.565 3.025 ;
      RECT 51.545 2.447 51.55 3.051 ;
      RECT 51.54 2.465 51.545 3.063 ;
      RECT 51.53 2.495 51.54 3.082 ;
      RECT 51.52 2.52 51.53 3.107 ;
      RECT 51.515 2.54 51.52 3.126 ;
      RECT 51.51 2.557 51.515 3.139 ;
      RECT 51.5 2.583 51.51 3.158 ;
      RECT 51.49 2.621 51.5 3.185 ;
      RECT 51.485 2.647 51.49 3.205 ;
      RECT 51.48 2.657 51.485 3.215 ;
      RECT 51.475 2.67 51.48 3.23 ;
      RECT 51.47 2.685 51.475 3.24 ;
      RECT 51.465 2.707 51.47 3.255 ;
      RECT 51.46 2.725 51.465 3.266 ;
      RECT 51.455 2.735 51.46 3.277 ;
      RECT 51.45 2.743 51.455 3.289 ;
      RECT 51.445 2.751 51.45 3.3 ;
      RECT 51.44 2.777 51.445 3.313 ;
      RECT 51.43 2.805 51.44 3.326 ;
      RECT 51.425 2.835 51.43 3.335 ;
      RECT 51.42 2.85 51.425 3.342 ;
      RECT 51.405 2.875 51.42 3.349 ;
      RECT 51.4 2.897 51.405 3.355 ;
      RECT 51.395 2.922 51.4 3.358 ;
      RECT 51.386 2.95 51.395 3.362 ;
      RECT 51.38 2.967 51.386 3.367 ;
      RECT 51.375 2.985 51.38 3.371 ;
      RECT 51.37 2.997 51.375 3.374 ;
      RECT 51.365 3.018 51.37 3.378 ;
      RECT 51.36 3.036 51.365 3.381 ;
      RECT 51.355 3.05 51.36 3.384 ;
      RECT 51.35 3.067 51.355 3.387 ;
      RECT 51.345 3.08 51.35 3.39 ;
      RECT 51.32 3.117 51.345 3.398 ;
      RECT 51.315 3.162 51.32 3.407 ;
      RECT 51.31 3.19 51.315 3.41 ;
      RECT 51.3 3.21 51.31 3.414 ;
      RECT 51.295 3.23 51.3 3.419 ;
      RECT 51.29 3.245 51.295 3.422 ;
      RECT 51.27 3.255 51.29 3.429 ;
      RECT 51.205 3.262 51.27 3.455 ;
      RECT 51.17 3.265 51.205 3.483 ;
      RECT 51.155 3.268 51.17 3.498 ;
      RECT 51.145 3.269 51.155 3.513 ;
      RECT 51.135 3.27 51.145 3.53 ;
      RECT 51.13 3.27 51.135 3.545 ;
      RECT 51.125 3.27 51.13 3.553 ;
      RECT 51.11 3.271 51.125 3.568 ;
      RECT 51.08 3.273 51.11 3.575 ;
      RECT 50.97 3.28 51.05 3.575 ;
      RECT 50.925 3.285 50.97 3.575 ;
      RECT 50.915 3.286 50.925 3.565 ;
      RECT 50.905 3.287 50.915 3.558 ;
      RECT 50.885 3.289 50.905 3.553 ;
      RECT 50.875 3.26 50.885 3.548 ;
      RECT 50.83 3.26 50.875 3.54 ;
      RECT 50.8 3.26 50.825 3.53 ;
      RECT 50.78 3.26 50.8 3.523 ;
      RECT 51.06 2.06 51.32 2.32 ;
      RECT 50.94 2.075 50.95 2.24 ;
      RECT 50.925 2.075 50.93 2.235 ;
      RECT 48.29 1.915 48.475 2.205 ;
      RECT 50.105 2.04 50.12 2.195 ;
      RECT 48.255 1.915 48.28 2.175 ;
      RECT 50.67 1.965 50.675 2.107 ;
      RECT 50.585 1.96 50.61 2.1 ;
      RECT 50.985 2.077 51.06 2.27 ;
      RECT 50.97 2.075 50.985 2.253 ;
      RECT 50.95 2.075 50.97 2.245 ;
      RECT 50.93 2.075 50.94 2.238 ;
      RECT 50.885 2.07 50.925 2.228 ;
      RECT 50.845 2.045 50.885 2.213 ;
      RECT 50.83 2.02 50.845 2.203 ;
      RECT 50.825 2.014 50.83 2.201 ;
      RECT 50.79 2.006 50.825 2.184 ;
      RECT 50.785 1.999 50.79 2.172 ;
      RECT 50.765 1.994 50.785 2.16 ;
      RECT 50.755 1.988 50.765 2.145 ;
      RECT 50.735 1.983 50.755 2.13 ;
      RECT 50.725 1.978 50.735 2.123 ;
      RECT 50.72 1.976 50.725 2.118 ;
      RECT 50.715 1.975 50.72 2.115 ;
      RECT 50.675 1.97 50.715 2.111 ;
      RECT 50.655 1.964 50.67 2.106 ;
      RECT 50.62 1.961 50.655 2.103 ;
      RECT 50.61 1.96 50.62 2.101 ;
      RECT 50.55 1.96 50.585 2.098 ;
      RECT 50.505 1.96 50.55 2.098 ;
      RECT 50.455 1.96 50.505 2.101 ;
      RECT 50.44 1.962 50.455 2.103 ;
      RECT 50.425 1.965 50.44 2.104 ;
      RECT 50.415 1.97 50.425 2.105 ;
      RECT 50.385 1.975 50.415 2.11 ;
      RECT 50.375 1.981 50.385 2.118 ;
      RECT 50.365 1.983 50.375 2.122 ;
      RECT 50.355 1.987 50.365 2.126 ;
      RECT 50.33 1.993 50.355 2.134 ;
      RECT 50.32 1.998 50.33 2.142 ;
      RECT 50.305 2.002 50.32 2.146 ;
      RECT 50.27 2.008 50.305 2.154 ;
      RECT 50.25 2.013 50.27 2.164 ;
      RECT 50.22 2.02 50.25 2.173 ;
      RECT 50.175 2.029 50.22 2.187 ;
      RECT 50.17 2.034 50.175 2.198 ;
      RECT 50.15 2.037 50.17 2.199 ;
      RECT 50.12 2.04 50.15 2.197 ;
      RECT 50.085 2.04 50.105 2.193 ;
      RECT 50.015 2.04 50.085 2.184 ;
      RECT 50 2.037 50.015 2.176 ;
      RECT 49.96 2.03 50 2.171 ;
      RECT 49.935 2.02 49.96 2.164 ;
      RECT 49.93 2.014 49.935 2.161 ;
      RECT 49.89 2.008 49.93 2.158 ;
      RECT 49.875 2.001 49.89 2.153 ;
      RECT 49.855 1.997 49.875 2.148 ;
      RECT 49.84 1.992 49.855 2.144 ;
      RECT 49.825 1.987 49.84 2.142 ;
      RECT 49.81 1.983 49.825 2.141 ;
      RECT 49.795 1.981 49.81 2.137 ;
      RECT 49.785 1.979 49.795 2.132 ;
      RECT 49.77 1.976 49.785 2.128 ;
      RECT 49.76 1.974 49.77 2.123 ;
      RECT 49.74 1.971 49.76 2.119 ;
      RECT 49.695 1.97 49.74 2.117 ;
      RECT 49.635 1.972 49.695 2.118 ;
      RECT 49.615 1.974 49.635 2.12 ;
      RECT 49.585 1.977 49.615 2.121 ;
      RECT 49.535 1.982 49.585 2.123 ;
      RECT 49.53 1.985 49.535 2.125 ;
      RECT 49.52 1.987 49.53 2.128 ;
      RECT 49.515 1.989 49.52 2.131 ;
      RECT 49.465 1.992 49.515 2.138 ;
      RECT 49.445 1.996 49.465 2.15 ;
      RECT 49.435 1.999 49.445 2.156 ;
      RECT 49.425 2 49.435 2.159 ;
      RECT 49.386 2.003 49.425 2.161 ;
      RECT 49.3 2.01 49.386 2.164 ;
      RECT 49.226 2.02 49.3 2.168 ;
      RECT 49.14 2.031 49.226 2.173 ;
      RECT 49.125 2.038 49.14 2.175 ;
      RECT 49.07 2.042 49.125 2.176 ;
      RECT 49.056 2.045 49.07 2.178 ;
      RECT 48.97 2.045 49.056 2.18 ;
      RECT 48.93 2.042 48.97 2.183 ;
      RECT 48.906 2.038 48.93 2.185 ;
      RECT 48.82 2.028 48.906 2.188 ;
      RECT 48.79 2.017 48.82 2.189 ;
      RECT 48.771 2.013 48.79 2.188 ;
      RECT 48.685 2.006 48.771 2.185 ;
      RECT 48.625 1.995 48.685 2.182 ;
      RECT 48.605 1.987 48.625 2.18 ;
      RECT 48.57 1.982 48.605 2.179 ;
      RECT 48.545 1.977 48.57 2.178 ;
      RECT 48.515 1.972 48.545 2.177 ;
      RECT 48.49 1.915 48.515 2.176 ;
      RECT 48.475 1.915 48.49 2.2 ;
      RECT 48.28 1.915 48.29 2.2 ;
      RECT 50.055 2.935 50.06 3.075 ;
      RECT 49.715 2.935 49.75 3.073 ;
      RECT 49.29 2.92 49.305 3.065 ;
      RECT 51.12 2.7 51.21 2.96 ;
      RECT 50.95 2.565 51.05 2.96 ;
      RECT 47.985 2.54 48.065 2.75 ;
      RECT 51.075 2.677 51.12 2.96 ;
      RECT 51.065 2.647 51.075 2.96 ;
      RECT 51.05 2.57 51.065 2.96 ;
      RECT 50.865 2.565 50.95 2.925 ;
      RECT 50.86 2.567 50.865 2.92 ;
      RECT 50.855 2.572 50.86 2.92 ;
      RECT 50.82 2.672 50.855 2.92 ;
      RECT 50.81 2.7 50.82 2.92 ;
      RECT 50.8 2.715 50.81 2.92 ;
      RECT 50.79 2.727 50.8 2.92 ;
      RECT 50.785 2.737 50.79 2.92 ;
      RECT 50.77 2.747 50.785 2.922 ;
      RECT 50.765 2.762 50.77 2.924 ;
      RECT 50.75 2.775 50.765 2.926 ;
      RECT 50.745 2.79 50.75 2.929 ;
      RECT 50.725 2.8 50.745 2.933 ;
      RECT 50.71 2.81 50.725 2.936 ;
      RECT 50.675 2.817 50.71 2.941 ;
      RECT 50.631 2.824 50.675 2.949 ;
      RECT 50.545 2.836 50.631 2.962 ;
      RECT 50.52 2.847 50.545 2.973 ;
      RECT 50.49 2.852 50.52 2.978 ;
      RECT 50.455 2.857 50.49 2.986 ;
      RECT 50.425 2.862 50.455 2.993 ;
      RECT 50.4 2.867 50.425 2.998 ;
      RECT 50.335 2.874 50.4 3.007 ;
      RECT 50.265 2.887 50.335 3.023 ;
      RECT 50.235 2.897 50.265 3.035 ;
      RECT 50.21 2.902 50.235 3.042 ;
      RECT 50.155 2.909 50.21 3.05 ;
      RECT 50.15 2.916 50.155 3.055 ;
      RECT 50.145 2.918 50.15 3.056 ;
      RECT 50.13 2.92 50.145 3.058 ;
      RECT 50.125 2.92 50.13 3.061 ;
      RECT 50.06 2.927 50.125 3.068 ;
      RECT 50.025 2.937 50.055 3.078 ;
      RECT 50.008 2.94 50.025 3.08 ;
      RECT 49.922 2.939 50.008 3.079 ;
      RECT 49.836 2.937 49.922 3.076 ;
      RECT 49.75 2.936 49.836 3.074 ;
      RECT 49.649 2.934 49.715 3.073 ;
      RECT 49.563 2.931 49.649 3.071 ;
      RECT 49.477 2.927 49.563 3.069 ;
      RECT 49.391 2.924 49.477 3.068 ;
      RECT 49.305 2.921 49.391 3.066 ;
      RECT 49.205 2.92 49.29 3.063 ;
      RECT 49.155 2.918 49.205 3.061 ;
      RECT 49.135 2.915 49.155 3.059 ;
      RECT 49.115 2.913 49.135 3.056 ;
      RECT 49.09 2.909 49.115 3.053 ;
      RECT 49.045 2.903 49.09 3.048 ;
      RECT 49.005 2.897 49.045 3.04 ;
      RECT 48.98 2.892 49.005 3.033 ;
      RECT 48.925 2.885 48.98 3.025 ;
      RECT 48.901 2.878 48.925 3.018 ;
      RECT 48.815 2.869 48.901 3.008 ;
      RECT 48.785 2.861 48.815 2.998 ;
      RECT 48.755 2.857 48.785 2.993 ;
      RECT 48.75 2.854 48.755 2.99 ;
      RECT 48.745 2.853 48.75 2.99 ;
      RECT 48.67 2.846 48.745 2.983 ;
      RECT 48.631 2.837 48.67 2.972 ;
      RECT 48.545 2.827 48.631 2.96 ;
      RECT 48.505 2.817 48.545 2.948 ;
      RECT 48.466 2.812 48.505 2.941 ;
      RECT 48.38 2.802 48.466 2.93 ;
      RECT 48.34 2.79 48.38 2.919 ;
      RECT 48.305 2.775 48.34 2.912 ;
      RECT 48.295 2.765 48.305 2.909 ;
      RECT 48.275 2.75 48.295 2.907 ;
      RECT 48.245 2.72 48.275 2.903 ;
      RECT 48.235 2.7 48.245 2.898 ;
      RECT 48.23 2.692 48.235 2.895 ;
      RECT 48.225 2.685 48.23 2.893 ;
      RECT 48.21 2.672 48.225 2.886 ;
      RECT 48.205 2.662 48.21 2.878 ;
      RECT 48.2 2.655 48.205 2.873 ;
      RECT 48.195 2.65 48.2 2.869 ;
      RECT 48.18 2.637 48.195 2.861 ;
      RECT 48.175 2.547 48.18 2.85 ;
      RECT 48.17 2.542 48.175 2.843 ;
      RECT 48.095 2.54 48.17 2.803 ;
      RECT 48.065 2.54 48.095 2.758 ;
      RECT 47.97 2.545 47.985 2.745 ;
      RECT 50.455 2.25 50.715 2.51 ;
      RECT 50.44 2.238 50.62 2.475 ;
      RECT 50.435 2.239 50.62 2.473 ;
      RECT 50.42 2.243 50.63 2.463 ;
      RECT 50.415 2.248 50.635 2.433 ;
      RECT 50.42 2.245 50.635 2.463 ;
      RECT 50.435 2.24 50.63 2.473 ;
      RECT 50.455 2.237 50.62 2.51 ;
      RECT 50.455 2.236 50.61 2.51 ;
      RECT 50.48 2.235 50.61 2.51 ;
      RECT 50.04 2.48 50.3 2.74 ;
      RECT 49.915 2.525 50.3 2.735 ;
      RECT 49.905 2.53 50.3 2.73 ;
      RECT 49.92 3.47 49.935 3.78 ;
      RECT 48.515 3.24 48.525 3.37 ;
      RECT 48.295 3.235 48.4 3.37 ;
      RECT 48.21 3.24 48.26 3.37 ;
      RECT 46.76 1.975 46.765 3.08 ;
      RECT 50.015 3.562 50.02 3.698 ;
      RECT 50.01 3.557 50.015 3.758 ;
      RECT 50.005 3.555 50.01 3.771 ;
      RECT 49.99 3.552 50.005 3.773 ;
      RECT 49.985 3.547 49.99 3.775 ;
      RECT 49.98 3.543 49.985 3.778 ;
      RECT 49.965 3.538 49.98 3.78 ;
      RECT 49.935 3.53 49.965 3.78 ;
      RECT 49.896 3.47 49.92 3.78 ;
      RECT 49.81 3.47 49.896 3.777 ;
      RECT 49.78 3.47 49.81 3.77 ;
      RECT 49.755 3.47 49.78 3.763 ;
      RECT 49.73 3.47 49.755 3.755 ;
      RECT 49.715 3.47 49.73 3.748 ;
      RECT 49.69 3.47 49.715 3.74 ;
      RECT 49.675 3.47 49.69 3.733 ;
      RECT 49.635 3.48 49.675 3.722 ;
      RECT 49.625 3.475 49.635 3.712 ;
      RECT 49.621 3.474 49.625 3.709 ;
      RECT 49.535 3.466 49.621 3.692 ;
      RECT 49.502 3.455 49.535 3.669 ;
      RECT 49.416 3.444 49.502 3.647 ;
      RECT 49.33 3.428 49.416 3.616 ;
      RECT 49.26 3.413 49.33 3.588 ;
      RECT 49.25 3.406 49.26 3.575 ;
      RECT 49.22 3.403 49.25 3.565 ;
      RECT 49.195 3.399 49.22 3.558 ;
      RECT 49.18 3.396 49.195 3.553 ;
      RECT 49.175 3.395 49.18 3.548 ;
      RECT 49.145 3.39 49.175 3.541 ;
      RECT 49.14 3.385 49.145 3.536 ;
      RECT 49.125 3.382 49.14 3.531 ;
      RECT 49.12 3.377 49.125 3.526 ;
      RECT 49.1 3.372 49.12 3.523 ;
      RECT 49.085 3.367 49.1 3.515 ;
      RECT 49.07 3.361 49.085 3.51 ;
      RECT 49.04 3.352 49.07 3.503 ;
      RECT 49.035 3.345 49.04 3.495 ;
      RECT 49.03 3.343 49.035 3.493 ;
      RECT 49.025 3.342 49.03 3.49 ;
      RECT 48.985 3.335 49.025 3.483 ;
      RECT 48.971 3.325 48.985 3.473 ;
      RECT 48.92 3.314 48.971 3.461 ;
      RECT 48.895 3.3 48.92 3.447 ;
      RECT 48.87 3.289 48.895 3.439 ;
      RECT 48.85 3.278 48.87 3.433 ;
      RECT 48.84 3.272 48.85 3.428 ;
      RECT 48.835 3.27 48.84 3.424 ;
      RECT 48.815 3.265 48.835 3.419 ;
      RECT 48.785 3.255 48.815 3.409 ;
      RECT 48.78 3.247 48.785 3.402 ;
      RECT 48.765 3.245 48.78 3.398 ;
      RECT 48.745 3.245 48.765 3.393 ;
      RECT 48.74 3.244 48.745 3.391 ;
      RECT 48.735 3.244 48.74 3.388 ;
      RECT 48.695 3.243 48.735 3.383 ;
      RECT 48.67 3.242 48.695 3.378 ;
      RECT 48.61 3.241 48.67 3.375 ;
      RECT 48.525 3.24 48.61 3.373 ;
      RECT 48.486 3.239 48.515 3.37 ;
      RECT 48.4 3.237 48.486 3.37 ;
      RECT 48.26 3.237 48.295 3.37 ;
      RECT 48.17 3.241 48.21 3.373 ;
      RECT 48.155 3.244 48.17 3.38 ;
      RECT 48.145 3.245 48.155 3.387 ;
      RECT 48.12 3.248 48.145 3.392 ;
      RECT 48.115 3.25 48.12 3.395 ;
      RECT 48.065 3.252 48.115 3.396 ;
      RECT 48.026 3.256 48.065 3.398 ;
      RECT 47.94 3.258 48.026 3.401 ;
      RECT 47.922 3.26 47.94 3.403 ;
      RECT 47.836 3.263 47.922 3.405 ;
      RECT 47.75 3.267 47.836 3.408 ;
      RECT 47.713 3.271 47.75 3.411 ;
      RECT 47.627 3.274 47.713 3.414 ;
      RECT 47.541 3.278 47.627 3.417 ;
      RECT 47.455 3.283 47.541 3.421 ;
      RECT 47.435 3.285 47.455 3.424 ;
      RECT 47.415 3.284 47.435 3.425 ;
      RECT 47.366 3.281 47.415 3.426 ;
      RECT 47.28 3.276 47.366 3.429 ;
      RECT 47.23 3.271 47.28 3.431 ;
      RECT 47.206 3.269 47.23 3.432 ;
      RECT 47.12 3.264 47.206 3.434 ;
      RECT 47.095 3.26 47.12 3.433 ;
      RECT 47.085 3.257 47.095 3.431 ;
      RECT 47.075 3.25 47.085 3.428 ;
      RECT 47.07 3.23 47.075 3.423 ;
      RECT 47.06 3.2 47.07 3.418 ;
      RECT 47.045 3.07 47.06 3.409 ;
      RECT 47.04 3.062 47.045 3.402 ;
      RECT 47.02 3.055 47.04 3.394 ;
      RECT 47.015 3.037 47.02 3.386 ;
      RECT 47.005 3.017 47.015 3.381 ;
      RECT 47 2.99 47.005 3.377 ;
      RECT 46.995 2.967 47 3.374 ;
      RECT 46.975 2.925 46.995 3.366 ;
      RECT 46.94 2.84 46.975 3.35 ;
      RECT 46.935 2.772 46.94 3.338 ;
      RECT 46.92 2.742 46.935 3.332 ;
      RECT 46.915 1.987 46.92 2.233 ;
      RECT 46.905 2.712 46.92 3.323 ;
      RECT 46.91 1.982 46.915 2.265 ;
      RECT 46.905 1.977 46.91 2.308 ;
      RECT 46.9 1.975 46.905 2.343 ;
      RECT 46.885 2.675 46.905 3.313 ;
      RECT 46.895 1.975 46.9 2.38 ;
      RECT 46.88 1.975 46.895 2.478 ;
      RECT 46.88 2.648 46.885 3.306 ;
      RECT 46.875 1.975 46.88 2.553 ;
      RECT 46.875 2.636 46.88 3.303 ;
      RECT 46.87 1.975 46.875 2.585 ;
      RECT 46.87 2.615 46.875 3.3 ;
      RECT 46.865 1.975 46.87 3.297 ;
      RECT 46.83 1.975 46.865 3.283 ;
      RECT 46.815 1.975 46.83 3.265 ;
      RECT 46.795 1.975 46.815 3.255 ;
      RECT 46.77 1.975 46.795 3.238 ;
      RECT 46.765 1.975 46.77 3.188 ;
      RECT 46.755 1.975 46.76 3.018 ;
      RECT 46.75 1.975 46.755 2.925 ;
      RECT 46.745 1.975 46.75 2.838 ;
      RECT 46.74 1.975 46.745 2.77 ;
      RECT 46.735 1.975 46.74 2.713 ;
      RECT 46.725 1.975 46.735 2.608 ;
      RECT 46.72 1.975 46.725 2.48 ;
      RECT 46.715 1.975 46.72 2.398 ;
      RECT 46.71 1.977 46.715 2.315 ;
      RECT 46.705 1.982 46.71 2.248 ;
      RECT 46.7 1.987 46.705 2.175 ;
      RECT 49.515 2.305 49.775 2.565 ;
      RECT 49.535 2.272 49.745 2.565 ;
      RECT 49.535 2.27 49.735 2.565 ;
      RECT 49.545 2.257 49.735 2.565 ;
      RECT 49.545 2.255 49.66 2.565 ;
      RECT 49.02 2.38 49.195 2.66 ;
      RECT 49.015 2.38 49.195 2.658 ;
      RECT 49.015 2.38 49.21 2.655 ;
      RECT 49.005 2.38 49.21 2.653 ;
      RECT 48.95 2.38 49.21 2.64 ;
      RECT 48.95 2.455 49.215 2.618 ;
      RECT 48.495 2.392 48.515 2.635 ;
      RECT 48.495 2.392 48.555 2.634 ;
      RECT 48.49 2.394 48.555 2.633 ;
      RECT 48.49 2.394 48.641 2.632 ;
      RECT 48.49 2.394 48.71 2.631 ;
      RECT 48.49 2.394 48.73 2.623 ;
      RECT 48.47 2.397 48.73 2.621 ;
      RECT 48.455 2.407 48.73 2.606 ;
      RECT 48.455 2.407 48.745 2.605 ;
      RECT 48.45 2.416 48.745 2.597 ;
      RECT 48.45 2.416 48.75 2.593 ;
      RECT 48.555 2.33 48.815 2.59 ;
      RECT 48.445 2.418 48.815 2.475 ;
      RECT 48.515 2.385 48.815 2.59 ;
      RECT 48.48 3.578 48.485 3.785 ;
      RECT 48.43 3.572 48.48 3.784 ;
      RECT 48.397 3.586 48.49 3.783 ;
      RECT 48.311 3.586 48.49 3.782 ;
      RECT 48.225 3.586 48.49 3.781 ;
      RECT 48.225 3.685 48.495 3.778 ;
      RECT 48.22 3.685 48.495 3.773 ;
      RECT 48.215 3.685 48.495 3.755 ;
      RECT 48.21 3.685 48.495 3.738 ;
      RECT 48.17 3.47 48.43 3.73 ;
      RECT 47.63 2.62 47.716 3.034 ;
      RECT 47.63 2.62 47.755 3.031 ;
      RECT 47.63 2.62 47.775 3.021 ;
      RECT 47.585 2.62 47.775 3.018 ;
      RECT 47.585 2.772 47.785 3.008 ;
      RECT 47.585 2.793 47.79 3.002 ;
      RECT 47.585 2.811 47.795 2.998 ;
      RECT 47.585 2.831 47.805 2.993 ;
      RECT 47.56 2.831 47.805 2.99 ;
      RECT 47.55 2.831 47.805 2.968 ;
      RECT 47.55 2.847 47.81 2.938 ;
      RECT 47.515 2.62 47.775 2.925 ;
      RECT 47.515 2.859 47.815 2.88 ;
      RECT 45.18 2.365 45.47 2.595 ;
      RECT 45.24 0.885 45.41 2.595 ;
      RECT 45.21 1.095 45.55 1.445 ;
      RECT 45.18 0.885 45.47 1.115 ;
      RECT 45.18 7.765 45.47 7.995 ;
      RECT 45.24 6.285 45.41 7.995 ;
      RECT 45.18 6.285 45.47 6.515 ;
      RECT 44.77 2.735 45.1 2.965 ;
      RECT 44.77 2.765 45.27 2.935 ;
      RECT 44.77 2.395 44.96 2.965 ;
      RECT 44.19 2.365 44.48 2.595 ;
      RECT 44.19 2.395 44.96 2.565 ;
      RECT 44.25 0.885 44.42 2.595 ;
      RECT 44.19 0.885 44.48 1.115 ;
      RECT 44.19 7.765 44.48 7.995 ;
      RECT 44.25 6.285 44.42 7.995 ;
      RECT 44.19 6.285 44.48 6.515 ;
      RECT 44.19 6.325 45.04 6.485 ;
      RECT 44.87 5.915 45.04 6.485 ;
      RECT 44.19 6.32 44.58 6.485 ;
      RECT 44.81 5.915 45.1 6.145 ;
      RECT 44.81 5.945 45.27 6.115 ;
      RECT 43.82 2.735 44.11 2.965 ;
      RECT 43.82 2.765 44.28 2.935 ;
      RECT 43.88 1.655 44.045 2.965 ;
      RECT 42.395 1.625 42.685 1.855 ;
      RECT 42.395 1.655 44.045 1.825 ;
      RECT 42.455 0.885 42.625 1.855 ;
      RECT 42.395 0.885 42.685 1.115 ;
      RECT 42.395 7.765 42.685 7.995 ;
      RECT 42.455 7.025 42.625 7.995 ;
      RECT 42.455 7.12 44.045 7.29 ;
      RECT 43.875 5.915 44.045 7.29 ;
      RECT 42.395 7.025 42.685 7.255 ;
      RECT 43.82 5.915 44.11 6.145 ;
      RECT 43.82 5.945 44.28 6.115 ;
      RECT 42.825 1.965 43.175 2.315 ;
      RECT 42.655 2.025 43.175 2.195 ;
      RECT 42.85 6.655 43.175 6.98 ;
      RECT 42.825 6.655 43.175 6.885 ;
      RECT 42.655 6.685 43.175 6.855 ;
      RECT 40.445 2.705 40.785 3.055 ;
      RECT 40.535 2.395 40.705 3.055 ;
      RECT 42.05 2.365 42.37 2.685 ;
      RECT 42.02 2.365 42.37 2.595 ;
      RECT 40.535 2.395 42.37 2.565 ;
      RECT 42.05 6.28 42.37 6.605 ;
      RECT 42.02 6.285 42.37 6.515 ;
      RECT 41.85 6.315 42.37 6.485 ;
      RECT 41.005 2.705 41.345 3.055 ;
      RECT 41.005 2.765 41.485 2.935 ;
      RECT 41 5.86 41.34 6.21 ;
      RECT 41 5.945 41.485 6.115 ;
      RECT 37.74 2.985 37.89 3.26 ;
      RECT 38.28 2.065 38.285 2.285 ;
      RECT 39.43 2.265 39.445 2.463 ;
      RECT 39.395 2.257 39.43 2.47 ;
      RECT 39.365 2.25 39.395 2.47 ;
      RECT 39.31 2.215 39.365 2.47 ;
      RECT 39.245 2.152 39.31 2.47 ;
      RECT 39.24 2.117 39.245 2.468 ;
      RECT 39.235 2.112 39.24 2.46 ;
      RECT 39.23 2.107 39.235 2.446 ;
      RECT 39.225 2.104 39.23 2.439 ;
      RECT 39.18 2.094 39.225 2.39 ;
      RECT 39.16 2.081 39.18 2.325 ;
      RECT 39.155 2.076 39.16 2.298 ;
      RECT 39.15 2.075 39.155 2.291 ;
      RECT 39.145 2.074 39.15 2.284 ;
      RECT 39.06 2.059 39.145 2.23 ;
      RECT 39.03 2.04 39.06 2.18 ;
      RECT 38.95 2.023 39.03 2.165 ;
      RECT 38.915 2.01 38.95 2.15 ;
      RECT 38.907 2.01 38.915 2.145 ;
      RECT 38.821 2.011 38.907 2.145 ;
      RECT 38.735 2.013 38.821 2.145 ;
      RECT 38.71 2.014 38.735 2.149 ;
      RECT 38.635 2.02 38.71 2.164 ;
      RECT 38.552 2.032 38.635 2.188 ;
      RECT 38.466 2.045 38.552 2.214 ;
      RECT 38.38 2.058 38.466 2.24 ;
      RECT 38.345 2.067 38.38 2.259 ;
      RECT 38.295 2.067 38.345 2.272 ;
      RECT 38.285 2.065 38.295 2.283 ;
      RECT 38.27 2.062 38.28 2.285 ;
      RECT 38.255 2.054 38.27 2.293 ;
      RECT 38.24 2.046 38.255 2.313 ;
      RECT 38.235 2.041 38.24 2.37 ;
      RECT 38.22 2.036 38.235 2.443 ;
      RECT 38.215 2.031 38.22 2.485 ;
      RECT 38.21 2.029 38.215 2.513 ;
      RECT 38.205 2.027 38.21 2.535 ;
      RECT 38.195 2.023 38.205 2.578 ;
      RECT 38.19 2.02 38.195 2.603 ;
      RECT 38.185 2.018 38.19 2.623 ;
      RECT 38.18 2.016 38.185 2.647 ;
      RECT 38.175 2.012 38.18 2.67 ;
      RECT 38.17 2.008 38.175 2.693 ;
      RECT 38.135 1.998 38.17 2.8 ;
      RECT 38.13 1.988 38.135 2.898 ;
      RECT 38.125 1.986 38.13 2.925 ;
      RECT 38.12 1.985 38.125 2.945 ;
      RECT 38.115 1.977 38.12 2.965 ;
      RECT 38.11 1.972 38.115 3 ;
      RECT 38.105 1.97 38.11 3.018 ;
      RECT 38.1 1.97 38.105 3.043 ;
      RECT 38.095 1.97 38.1 3.065 ;
      RECT 38.06 1.97 38.095 3.108 ;
      RECT 38.035 1.97 38.06 3.137 ;
      RECT 38.025 1.97 38.035 2.323 ;
      RECT 38.028 2.38 38.035 3.147 ;
      RECT 38.025 2.437 38.028 3.15 ;
      RECT 38.02 1.97 38.025 2.295 ;
      RECT 38.02 2.487 38.025 3.153 ;
      RECT 38.01 1.97 38.02 2.285 ;
      RECT 38.015 2.54 38.02 3.156 ;
      RECT 38.01 2.625 38.015 3.16 ;
      RECT 38 1.97 38.01 2.273 ;
      RECT 38.005 2.672 38.01 3.164 ;
      RECT 38 2.747 38.005 3.168 ;
      RECT 37.965 1.97 38 2.248 ;
      RECT 37.99 2.83 38 3.173 ;
      RECT 37.98 2.897 37.99 3.18 ;
      RECT 37.975 2.925 37.98 3.185 ;
      RECT 37.965 2.938 37.975 3.191 ;
      RECT 37.92 1.97 37.965 2.205 ;
      RECT 37.96 2.943 37.965 3.198 ;
      RECT 37.92 2.96 37.96 3.26 ;
      RECT 37.915 1.972 37.92 2.178 ;
      RECT 37.89 2.98 37.92 3.26 ;
      RECT 37.91 1.977 37.915 2.15 ;
      RECT 37.7 2.989 37.74 3.26 ;
      RECT 37.675 2.997 37.7 3.23 ;
      RECT 37.63 3.005 37.675 3.23 ;
      RECT 37.615 3.01 37.63 3.225 ;
      RECT 37.605 3.01 37.615 3.219 ;
      RECT 37.595 3.017 37.605 3.216 ;
      RECT 37.59 3.055 37.595 3.205 ;
      RECT 37.585 3.117 37.59 3.183 ;
      RECT 38.855 2.992 39.04 3.215 ;
      RECT 38.855 3.007 39.045 3.211 ;
      RECT 38.845 2.28 38.93 3.21 ;
      RECT 38.845 3.007 39.05 3.204 ;
      RECT 38.84 3.015 39.05 3.203 ;
      RECT 39.045 2.735 39.365 3.055 ;
      RECT 38.84 2.907 39.01 2.998 ;
      RECT 38.835 2.907 39.01 2.98 ;
      RECT 38.825 2.715 38.96 2.955 ;
      RECT 38.82 2.715 38.96 2.9 ;
      RECT 38.78 2.295 38.95 2.8 ;
      RECT 38.765 2.295 38.95 2.67 ;
      RECT 38.76 2.295 38.95 2.623 ;
      RECT 38.755 2.295 38.95 2.603 ;
      RECT 38.75 2.295 38.95 2.578 ;
      RECT 38.72 2.295 38.98 2.555 ;
      RECT 38.73 2.292 38.94 2.555 ;
      RECT 38.855 2.287 38.94 3.215 ;
      RECT 38.74 2.28 38.93 2.555 ;
      RECT 38.735 2.285 38.93 2.555 ;
      RECT 37.565 2.497 37.75 2.71 ;
      RECT 37.565 2.505 37.76 2.703 ;
      RECT 37.545 2.505 37.76 2.7 ;
      RECT 37.54 2.505 37.76 2.685 ;
      RECT 37.47 2.42 37.73 2.68 ;
      RECT 37.47 2.565 37.765 2.593 ;
      RECT 37.125 3.02 37.385 3.28 ;
      RECT 37.15 2.965 37.345 3.28 ;
      RECT 37.145 2.714 37.325 3.008 ;
      RECT 37.145 2.72 37.335 3.008 ;
      RECT 37.125 2.722 37.335 2.953 ;
      RECT 37.12 2.732 37.335 2.82 ;
      RECT 37.15 2.712 37.325 3.28 ;
      RECT 37.236 2.71 37.325 3.28 ;
      RECT 37.095 1.93 37.13 2.3 ;
      RECT 36.885 2.04 36.89 2.3 ;
      RECT 37.13 1.937 37.145 2.3 ;
      RECT 37.02 1.93 37.095 2.378 ;
      RECT 37.01 1.93 37.02 2.463 ;
      RECT 36.985 1.93 37.01 2.498 ;
      RECT 36.945 1.93 36.985 2.566 ;
      RECT 36.935 1.937 36.945 2.618 ;
      RECT 36.905 2.04 36.935 2.659 ;
      RECT 36.9 2.04 36.905 2.698 ;
      RECT 36.89 2.04 36.9 2.718 ;
      RECT 36.885 2.335 36.89 2.755 ;
      RECT 36.88 2.352 36.885 2.775 ;
      RECT 36.865 2.415 36.88 2.815 ;
      RECT 36.86 2.458 36.865 2.85 ;
      RECT 36.855 2.466 36.86 2.863 ;
      RECT 36.845 2.48 36.855 2.885 ;
      RECT 36.82 2.515 36.845 2.95 ;
      RECT 36.81 2.55 36.82 3.013 ;
      RECT 36.79 2.58 36.81 3.074 ;
      RECT 36.775 2.616 36.79 3.141 ;
      RECT 36.765 2.644 36.775 3.18 ;
      RECT 36.755 2.666 36.765 3.2 ;
      RECT 36.75 2.676 36.755 3.211 ;
      RECT 36.745 2.685 36.75 3.214 ;
      RECT 36.735 2.703 36.745 3.218 ;
      RECT 36.725 2.721 36.735 3.219 ;
      RECT 36.7 2.76 36.725 3.216 ;
      RECT 36.68 2.802 36.7 3.213 ;
      RECT 36.665 2.84 36.68 3.212 ;
      RECT 36.63 2.875 36.665 3.209 ;
      RECT 36.625 2.897 36.63 3.207 ;
      RECT 36.56 2.937 36.625 3.204 ;
      RECT 36.555 2.977 36.56 3.2 ;
      RECT 36.54 2.987 36.555 3.191 ;
      RECT 36.53 3.107 36.54 3.176 ;
      RECT 37.01 3.52 37.02 3.78 ;
      RECT 37.01 3.523 37.03 3.779 ;
      RECT 37 3.513 37.01 3.778 ;
      RECT 36.99 3.528 37.07 3.774 ;
      RECT 36.975 3.507 36.99 3.772 ;
      RECT 36.95 3.532 37.075 3.768 ;
      RECT 36.935 3.492 36.95 3.763 ;
      RECT 36.935 3.534 37.085 3.762 ;
      RECT 36.935 3.542 37.1 3.755 ;
      RECT 36.875 3.479 36.935 3.745 ;
      RECT 36.865 3.466 36.875 3.727 ;
      RECT 36.84 3.456 36.865 3.717 ;
      RECT 36.835 3.446 36.84 3.709 ;
      RECT 36.77 3.542 37.1 3.691 ;
      RECT 36.685 3.542 37.1 3.653 ;
      RECT 36.575 3.37 36.835 3.63 ;
      RECT 36.95 3.5 36.975 3.768 ;
      RECT 36.99 3.51 37 3.774 ;
      RECT 36.575 3.518 37.015 3.63 ;
      RECT 35.79 3.275 35.82 3.575 ;
      RECT 35.565 3.26 35.57 3.535 ;
      RECT 35.365 3.26 35.52 3.52 ;
      RECT 36.665 1.975 36.695 2.235 ;
      RECT 36.655 1.975 36.665 2.343 ;
      RECT 36.635 1.975 36.655 2.353 ;
      RECT 36.62 1.975 36.635 2.365 ;
      RECT 36.565 1.975 36.62 2.415 ;
      RECT 36.55 1.975 36.565 2.463 ;
      RECT 36.52 1.975 36.55 2.498 ;
      RECT 36.465 1.975 36.52 2.56 ;
      RECT 36.445 1.975 36.465 2.628 ;
      RECT 36.44 1.975 36.445 2.658 ;
      RECT 36.435 1.975 36.44 2.67 ;
      RECT 36.43 2.092 36.435 2.688 ;
      RECT 36.41 2.11 36.43 2.713 ;
      RECT 36.39 2.137 36.41 2.763 ;
      RECT 36.385 2.157 36.39 2.794 ;
      RECT 36.38 2.165 36.385 2.811 ;
      RECT 36.365 2.191 36.38 2.84 ;
      RECT 36.35 2.233 36.365 2.875 ;
      RECT 36.345 2.262 36.35 2.898 ;
      RECT 36.34 2.277 36.345 2.911 ;
      RECT 36.335 2.3 36.34 2.922 ;
      RECT 36.325 2.32 36.335 2.94 ;
      RECT 36.315 2.35 36.325 2.963 ;
      RECT 36.31 2.372 36.315 2.983 ;
      RECT 36.305 2.387 36.31 2.998 ;
      RECT 36.29 2.417 36.305 3.025 ;
      RECT 36.285 2.447 36.29 3.051 ;
      RECT 36.28 2.465 36.285 3.063 ;
      RECT 36.27 2.495 36.28 3.082 ;
      RECT 36.26 2.52 36.27 3.107 ;
      RECT 36.255 2.54 36.26 3.126 ;
      RECT 36.25 2.557 36.255 3.139 ;
      RECT 36.24 2.583 36.25 3.158 ;
      RECT 36.23 2.621 36.24 3.185 ;
      RECT 36.225 2.647 36.23 3.205 ;
      RECT 36.22 2.657 36.225 3.215 ;
      RECT 36.215 2.67 36.22 3.23 ;
      RECT 36.21 2.685 36.215 3.24 ;
      RECT 36.205 2.707 36.21 3.255 ;
      RECT 36.2 2.725 36.205 3.266 ;
      RECT 36.195 2.735 36.2 3.277 ;
      RECT 36.19 2.743 36.195 3.289 ;
      RECT 36.185 2.751 36.19 3.3 ;
      RECT 36.18 2.777 36.185 3.313 ;
      RECT 36.17 2.805 36.18 3.326 ;
      RECT 36.165 2.835 36.17 3.335 ;
      RECT 36.16 2.85 36.165 3.342 ;
      RECT 36.145 2.875 36.16 3.349 ;
      RECT 36.14 2.897 36.145 3.355 ;
      RECT 36.135 2.922 36.14 3.358 ;
      RECT 36.126 2.95 36.135 3.362 ;
      RECT 36.12 2.967 36.126 3.367 ;
      RECT 36.115 2.985 36.12 3.371 ;
      RECT 36.11 2.997 36.115 3.374 ;
      RECT 36.105 3.018 36.11 3.378 ;
      RECT 36.1 3.036 36.105 3.381 ;
      RECT 36.095 3.05 36.1 3.384 ;
      RECT 36.09 3.067 36.095 3.387 ;
      RECT 36.085 3.08 36.09 3.39 ;
      RECT 36.06 3.117 36.085 3.398 ;
      RECT 36.055 3.162 36.06 3.407 ;
      RECT 36.05 3.19 36.055 3.41 ;
      RECT 36.04 3.21 36.05 3.414 ;
      RECT 36.035 3.23 36.04 3.419 ;
      RECT 36.03 3.245 36.035 3.422 ;
      RECT 36.01 3.255 36.03 3.429 ;
      RECT 35.945 3.262 36.01 3.455 ;
      RECT 35.91 3.265 35.945 3.483 ;
      RECT 35.895 3.268 35.91 3.498 ;
      RECT 35.885 3.269 35.895 3.513 ;
      RECT 35.875 3.27 35.885 3.53 ;
      RECT 35.87 3.27 35.875 3.545 ;
      RECT 35.865 3.27 35.87 3.553 ;
      RECT 35.85 3.271 35.865 3.568 ;
      RECT 35.82 3.273 35.85 3.575 ;
      RECT 35.71 3.28 35.79 3.575 ;
      RECT 35.665 3.285 35.71 3.575 ;
      RECT 35.655 3.286 35.665 3.565 ;
      RECT 35.645 3.287 35.655 3.558 ;
      RECT 35.625 3.289 35.645 3.553 ;
      RECT 35.615 3.26 35.625 3.548 ;
      RECT 35.57 3.26 35.615 3.54 ;
      RECT 35.54 3.26 35.565 3.53 ;
      RECT 35.52 3.26 35.54 3.523 ;
      RECT 35.8 2.06 36.06 2.32 ;
      RECT 35.68 2.075 35.69 2.24 ;
      RECT 35.665 2.075 35.67 2.235 ;
      RECT 33.03 1.915 33.215 2.205 ;
      RECT 34.845 2.04 34.86 2.195 ;
      RECT 32.995 1.915 33.02 2.175 ;
      RECT 35.41 1.965 35.415 2.107 ;
      RECT 35.325 1.96 35.35 2.1 ;
      RECT 35.725 2.077 35.8 2.27 ;
      RECT 35.71 2.075 35.725 2.253 ;
      RECT 35.69 2.075 35.71 2.245 ;
      RECT 35.67 2.075 35.68 2.238 ;
      RECT 35.625 2.07 35.665 2.228 ;
      RECT 35.585 2.045 35.625 2.213 ;
      RECT 35.57 2.02 35.585 2.203 ;
      RECT 35.565 2.014 35.57 2.201 ;
      RECT 35.53 2.006 35.565 2.184 ;
      RECT 35.525 1.999 35.53 2.172 ;
      RECT 35.505 1.994 35.525 2.16 ;
      RECT 35.495 1.988 35.505 2.145 ;
      RECT 35.475 1.983 35.495 2.13 ;
      RECT 35.465 1.978 35.475 2.123 ;
      RECT 35.46 1.976 35.465 2.118 ;
      RECT 35.455 1.975 35.46 2.115 ;
      RECT 35.415 1.97 35.455 2.111 ;
      RECT 35.395 1.964 35.41 2.106 ;
      RECT 35.36 1.961 35.395 2.103 ;
      RECT 35.35 1.96 35.36 2.101 ;
      RECT 35.29 1.96 35.325 2.098 ;
      RECT 35.245 1.96 35.29 2.098 ;
      RECT 35.195 1.96 35.245 2.101 ;
      RECT 35.18 1.962 35.195 2.103 ;
      RECT 35.165 1.965 35.18 2.104 ;
      RECT 35.155 1.97 35.165 2.105 ;
      RECT 35.125 1.975 35.155 2.11 ;
      RECT 35.115 1.981 35.125 2.118 ;
      RECT 35.105 1.983 35.115 2.122 ;
      RECT 35.095 1.987 35.105 2.126 ;
      RECT 35.07 1.993 35.095 2.134 ;
      RECT 35.06 1.998 35.07 2.142 ;
      RECT 35.045 2.002 35.06 2.146 ;
      RECT 35.01 2.008 35.045 2.154 ;
      RECT 34.99 2.013 35.01 2.164 ;
      RECT 34.96 2.02 34.99 2.173 ;
      RECT 34.915 2.029 34.96 2.187 ;
      RECT 34.91 2.034 34.915 2.198 ;
      RECT 34.89 2.037 34.91 2.199 ;
      RECT 34.86 2.04 34.89 2.197 ;
      RECT 34.825 2.04 34.845 2.193 ;
      RECT 34.755 2.04 34.825 2.184 ;
      RECT 34.74 2.037 34.755 2.176 ;
      RECT 34.7 2.03 34.74 2.171 ;
      RECT 34.675 2.02 34.7 2.164 ;
      RECT 34.67 2.014 34.675 2.161 ;
      RECT 34.63 2.008 34.67 2.158 ;
      RECT 34.615 2.001 34.63 2.153 ;
      RECT 34.595 1.997 34.615 2.148 ;
      RECT 34.58 1.992 34.595 2.144 ;
      RECT 34.565 1.987 34.58 2.142 ;
      RECT 34.55 1.983 34.565 2.141 ;
      RECT 34.535 1.981 34.55 2.137 ;
      RECT 34.525 1.979 34.535 2.132 ;
      RECT 34.51 1.976 34.525 2.128 ;
      RECT 34.5 1.974 34.51 2.123 ;
      RECT 34.48 1.971 34.5 2.119 ;
      RECT 34.435 1.97 34.48 2.117 ;
      RECT 34.375 1.972 34.435 2.118 ;
      RECT 34.355 1.974 34.375 2.12 ;
      RECT 34.325 1.977 34.355 2.121 ;
      RECT 34.275 1.982 34.325 2.123 ;
      RECT 34.27 1.985 34.275 2.125 ;
      RECT 34.26 1.987 34.27 2.128 ;
      RECT 34.255 1.989 34.26 2.131 ;
      RECT 34.205 1.992 34.255 2.138 ;
      RECT 34.185 1.996 34.205 2.15 ;
      RECT 34.175 1.999 34.185 2.156 ;
      RECT 34.165 2 34.175 2.159 ;
      RECT 34.126 2.003 34.165 2.161 ;
      RECT 34.04 2.01 34.126 2.164 ;
      RECT 33.966 2.02 34.04 2.168 ;
      RECT 33.88 2.031 33.966 2.173 ;
      RECT 33.865 2.038 33.88 2.175 ;
      RECT 33.81 2.042 33.865 2.176 ;
      RECT 33.796 2.045 33.81 2.178 ;
      RECT 33.71 2.045 33.796 2.18 ;
      RECT 33.67 2.042 33.71 2.183 ;
      RECT 33.646 2.038 33.67 2.185 ;
      RECT 33.56 2.028 33.646 2.188 ;
      RECT 33.53 2.017 33.56 2.189 ;
      RECT 33.511 2.013 33.53 2.188 ;
      RECT 33.425 2.006 33.511 2.185 ;
      RECT 33.365 1.995 33.425 2.182 ;
      RECT 33.345 1.987 33.365 2.18 ;
      RECT 33.31 1.982 33.345 2.179 ;
      RECT 33.285 1.977 33.31 2.178 ;
      RECT 33.255 1.972 33.285 2.177 ;
      RECT 33.23 1.915 33.255 2.176 ;
      RECT 33.215 1.915 33.23 2.2 ;
      RECT 33.02 1.915 33.03 2.2 ;
      RECT 34.795 2.935 34.8 3.075 ;
      RECT 34.455 2.935 34.49 3.073 ;
      RECT 34.03 2.92 34.045 3.065 ;
      RECT 35.86 2.7 35.95 2.96 ;
      RECT 35.69 2.565 35.79 2.96 ;
      RECT 32.725 2.54 32.805 2.75 ;
      RECT 35.815 2.677 35.86 2.96 ;
      RECT 35.805 2.647 35.815 2.96 ;
      RECT 35.79 2.57 35.805 2.96 ;
      RECT 35.605 2.565 35.69 2.925 ;
      RECT 35.6 2.567 35.605 2.92 ;
      RECT 35.595 2.572 35.6 2.92 ;
      RECT 35.56 2.672 35.595 2.92 ;
      RECT 35.55 2.7 35.56 2.92 ;
      RECT 35.54 2.715 35.55 2.92 ;
      RECT 35.53 2.727 35.54 2.92 ;
      RECT 35.525 2.737 35.53 2.92 ;
      RECT 35.51 2.747 35.525 2.922 ;
      RECT 35.505 2.762 35.51 2.924 ;
      RECT 35.49 2.775 35.505 2.926 ;
      RECT 35.485 2.79 35.49 2.929 ;
      RECT 35.465 2.8 35.485 2.933 ;
      RECT 35.45 2.81 35.465 2.936 ;
      RECT 35.415 2.817 35.45 2.941 ;
      RECT 35.371 2.824 35.415 2.949 ;
      RECT 35.285 2.836 35.371 2.962 ;
      RECT 35.26 2.847 35.285 2.973 ;
      RECT 35.23 2.852 35.26 2.978 ;
      RECT 35.195 2.857 35.23 2.986 ;
      RECT 35.165 2.862 35.195 2.993 ;
      RECT 35.14 2.867 35.165 2.998 ;
      RECT 35.075 2.874 35.14 3.007 ;
      RECT 35.005 2.887 35.075 3.023 ;
      RECT 34.975 2.897 35.005 3.035 ;
      RECT 34.95 2.902 34.975 3.042 ;
      RECT 34.895 2.909 34.95 3.05 ;
      RECT 34.89 2.916 34.895 3.055 ;
      RECT 34.885 2.918 34.89 3.056 ;
      RECT 34.87 2.92 34.885 3.058 ;
      RECT 34.865 2.92 34.87 3.061 ;
      RECT 34.8 2.927 34.865 3.068 ;
      RECT 34.765 2.937 34.795 3.078 ;
      RECT 34.748 2.94 34.765 3.08 ;
      RECT 34.662 2.939 34.748 3.079 ;
      RECT 34.576 2.937 34.662 3.076 ;
      RECT 34.49 2.936 34.576 3.074 ;
      RECT 34.389 2.934 34.455 3.073 ;
      RECT 34.303 2.931 34.389 3.071 ;
      RECT 34.217 2.927 34.303 3.069 ;
      RECT 34.131 2.924 34.217 3.068 ;
      RECT 34.045 2.921 34.131 3.066 ;
      RECT 33.945 2.92 34.03 3.063 ;
      RECT 33.895 2.918 33.945 3.061 ;
      RECT 33.875 2.915 33.895 3.059 ;
      RECT 33.855 2.913 33.875 3.056 ;
      RECT 33.83 2.909 33.855 3.053 ;
      RECT 33.785 2.903 33.83 3.048 ;
      RECT 33.745 2.897 33.785 3.04 ;
      RECT 33.72 2.892 33.745 3.033 ;
      RECT 33.665 2.885 33.72 3.025 ;
      RECT 33.641 2.878 33.665 3.018 ;
      RECT 33.555 2.869 33.641 3.008 ;
      RECT 33.525 2.861 33.555 2.998 ;
      RECT 33.495 2.857 33.525 2.993 ;
      RECT 33.49 2.854 33.495 2.99 ;
      RECT 33.485 2.853 33.49 2.99 ;
      RECT 33.41 2.846 33.485 2.983 ;
      RECT 33.371 2.837 33.41 2.972 ;
      RECT 33.285 2.827 33.371 2.96 ;
      RECT 33.245 2.817 33.285 2.948 ;
      RECT 33.206 2.812 33.245 2.941 ;
      RECT 33.12 2.802 33.206 2.93 ;
      RECT 33.08 2.79 33.12 2.919 ;
      RECT 33.045 2.775 33.08 2.912 ;
      RECT 33.035 2.765 33.045 2.909 ;
      RECT 33.015 2.75 33.035 2.907 ;
      RECT 32.985 2.72 33.015 2.903 ;
      RECT 32.975 2.7 32.985 2.898 ;
      RECT 32.97 2.692 32.975 2.895 ;
      RECT 32.965 2.685 32.97 2.893 ;
      RECT 32.95 2.672 32.965 2.886 ;
      RECT 32.945 2.662 32.95 2.878 ;
      RECT 32.94 2.655 32.945 2.873 ;
      RECT 32.935 2.65 32.94 2.869 ;
      RECT 32.92 2.637 32.935 2.861 ;
      RECT 32.915 2.547 32.92 2.85 ;
      RECT 32.91 2.542 32.915 2.843 ;
      RECT 32.835 2.54 32.91 2.803 ;
      RECT 32.805 2.54 32.835 2.758 ;
      RECT 32.71 2.545 32.725 2.745 ;
      RECT 35.195 2.25 35.455 2.51 ;
      RECT 35.18 2.238 35.36 2.475 ;
      RECT 35.175 2.239 35.36 2.473 ;
      RECT 35.16 2.243 35.37 2.463 ;
      RECT 35.155 2.248 35.375 2.433 ;
      RECT 35.16 2.245 35.375 2.463 ;
      RECT 35.175 2.24 35.37 2.473 ;
      RECT 35.195 2.237 35.36 2.51 ;
      RECT 35.195 2.236 35.35 2.51 ;
      RECT 35.22 2.235 35.35 2.51 ;
      RECT 34.78 2.48 35.04 2.74 ;
      RECT 34.655 2.525 35.04 2.735 ;
      RECT 34.645 2.53 35.04 2.73 ;
      RECT 34.66 3.47 34.675 3.78 ;
      RECT 33.255 3.24 33.265 3.37 ;
      RECT 33.035 3.235 33.14 3.37 ;
      RECT 32.95 3.24 33 3.37 ;
      RECT 31.5 1.975 31.505 3.08 ;
      RECT 34.755 3.562 34.76 3.698 ;
      RECT 34.75 3.557 34.755 3.758 ;
      RECT 34.745 3.555 34.75 3.771 ;
      RECT 34.73 3.552 34.745 3.773 ;
      RECT 34.725 3.547 34.73 3.775 ;
      RECT 34.72 3.543 34.725 3.778 ;
      RECT 34.705 3.538 34.72 3.78 ;
      RECT 34.675 3.53 34.705 3.78 ;
      RECT 34.636 3.47 34.66 3.78 ;
      RECT 34.55 3.47 34.636 3.777 ;
      RECT 34.52 3.47 34.55 3.77 ;
      RECT 34.495 3.47 34.52 3.763 ;
      RECT 34.47 3.47 34.495 3.755 ;
      RECT 34.455 3.47 34.47 3.748 ;
      RECT 34.43 3.47 34.455 3.74 ;
      RECT 34.415 3.47 34.43 3.733 ;
      RECT 34.375 3.48 34.415 3.722 ;
      RECT 34.365 3.475 34.375 3.712 ;
      RECT 34.361 3.474 34.365 3.709 ;
      RECT 34.275 3.466 34.361 3.692 ;
      RECT 34.242 3.455 34.275 3.669 ;
      RECT 34.156 3.444 34.242 3.647 ;
      RECT 34.07 3.428 34.156 3.616 ;
      RECT 34 3.413 34.07 3.588 ;
      RECT 33.99 3.406 34 3.575 ;
      RECT 33.96 3.403 33.99 3.565 ;
      RECT 33.935 3.399 33.96 3.558 ;
      RECT 33.92 3.396 33.935 3.553 ;
      RECT 33.915 3.395 33.92 3.548 ;
      RECT 33.885 3.39 33.915 3.541 ;
      RECT 33.88 3.385 33.885 3.536 ;
      RECT 33.865 3.382 33.88 3.531 ;
      RECT 33.86 3.377 33.865 3.526 ;
      RECT 33.84 3.372 33.86 3.523 ;
      RECT 33.825 3.367 33.84 3.515 ;
      RECT 33.81 3.361 33.825 3.51 ;
      RECT 33.78 3.352 33.81 3.503 ;
      RECT 33.775 3.345 33.78 3.495 ;
      RECT 33.77 3.343 33.775 3.493 ;
      RECT 33.765 3.342 33.77 3.49 ;
      RECT 33.725 3.335 33.765 3.483 ;
      RECT 33.711 3.325 33.725 3.473 ;
      RECT 33.66 3.314 33.711 3.461 ;
      RECT 33.635 3.3 33.66 3.447 ;
      RECT 33.61 3.289 33.635 3.439 ;
      RECT 33.59 3.278 33.61 3.433 ;
      RECT 33.58 3.272 33.59 3.428 ;
      RECT 33.575 3.27 33.58 3.424 ;
      RECT 33.555 3.265 33.575 3.419 ;
      RECT 33.525 3.255 33.555 3.409 ;
      RECT 33.52 3.247 33.525 3.402 ;
      RECT 33.505 3.245 33.52 3.398 ;
      RECT 33.485 3.245 33.505 3.393 ;
      RECT 33.48 3.244 33.485 3.391 ;
      RECT 33.475 3.244 33.48 3.388 ;
      RECT 33.435 3.243 33.475 3.383 ;
      RECT 33.41 3.242 33.435 3.378 ;
      RECT 33.35 3.241 33.41 3.375 ;
      RECT 33.265 3.24 33.35 3.373 ;
      RECT 33.226 3.239 33.255 3.37 ;
      RECT 33.14 3.237 33.226 3.37 ;
      RECT 33 3.237 33.035 3.37 ;
      RECT 32.91 3.241 32.95 3.373 ;
      RECT 32.895 3.244 32.91 3.38 ;
      RECT 32.885 3.245 32.895 3.387 ;
      RECT 32.86 3.248 32.885 3.392 ;
      RECT 32.855 3.25 32.86 3.395 ;
      RECT 32.805 3.252 32.855 3.396 ;
      RECT 32.766 3.256 32.805 3.398 ;
      RECT 32.68 3.258 32.766 3.401 ;
      RECT 32.662 3.26 32.68 3.403 ;
      RECT 32.576 3.263 32.662 3.405 ;
      RECT 32.49 3.267 32.576 3.408 ;
      RECT 32.453 3.271 32.49 3.411 ;
      RECT 32.367 3.274 32.453 3.414 ;
      RECT 32.281 3.278 32.367 3.417 ;
      RECT 32.195 3.283 32.281 3.421 ;
      RECT 32.175 3.285 32.195 3.424 ;
      RECT 32.155 3.284 32.175 3.425 ;
      RECT 32.106 3.281 32.155 3.426 ;
      RECT 32.02 3.276 32.106 3.429 ;
      RECT 31.97 3.271 32.02 3.431 ;
      RECT 31.946 3.269 31.97 3.432 ;
      RECT 31.86 3.264 31.946 3.434 ;
      RECT 31.835 3.26 31.86 3.433 ;
      RECT 31.825 3.257 31.835 3.431 ;
      RECT 31.815 3.25 31.825 3.428 ;
      RECT 31.81 3.23 31.815 3.423 ;
      RECT 31.8 3.2 31.81 3.418 ;
      RECT 31.785 3.07 31.8 3.409 ;
      RECT 31.78 3.062 31.785 3.402 ;
      RECT 31.76 3.055 31.78 3.394 ;
      RECT 31.755 3.037 31.76 3.386 ;
      RECT 31.745 3.017 31.755 3.381 ;
      RECT 31.74 2.99 31.745 3.377 ;
      RECT 31.735 2.967 31.74 3.374 ;
      RECT 31.715 2.925 31.735 3.366 ;
      RECT 31.68 2.84 31.715 3.35 ;
      RECT 31.675 2.772 31.68 3.338 ;
      RECT 31.66 2.742 31.675 3.332 ;
      RECT 31.655 1.987 31.66 2.233 ;
      RECT 31.645 2.712 31.66 3.323 ;
      RECT 31.65 1.982 31.655 2.265 ;
      RECT 31.645 1.977 31.65 2.308 ;
      RECT 31.64 1.975 31.645 2.343 ;
      RECT 31.625 2.675 31.645 3.313 ;
      RECT 31.635 1.975 31.64 2.38 ;
      RECT 31.62 1.975 31.635 2.478 ;
      RECT 31.62 2.648 31.625 3.306 ;
      RECT 31.615 1.975 31.62 2.553 ;
      RECT 31.615 2.636 31.62 3.303 ;
      RECT 31.61 1.975 31.615 2.585 ;
      RECT 31.61 2.615 31.615 3.3 ;
      RECT 31.605 1.975 31.61 3.297 ;
      RECT 31.57 1.975 31.605 3.283 ;
      RECT 31.555 1.975 31.57 3.265 ;
      RECT 31.535 1.975 31.555 3.255 ;
      RECT 31.51 1.975 31.535 3.238 ;
      RECT 31.505 1.975 31.51 3.188 ;
      RECT 31.495 1.975 31.5 3.018 ;
      RECT 31.49 1.975 31.495 2.925 ;
      RECT 31.485 1.975 31.49 2.838 ;
      RECT 31.48 1.975 31.485 2.77 ;
      RECT 31.475 1.975 31.48 2.713 ;
      RECT 31.465 1.975 31.475 2.608 ;
      RECT 31.46 1.975 31.465 2.48 ;
      RECT 31.455 1.975 31.46 2.398 ;
      RECT 31.45 1.977 31.455 2.315 ;
      RECT 31.445 1.982 31.45 2.248 ;
      RECT 31.44 1.987 31.445 2.175 ;
      RECT 34.255 2.305 34.515 2.565 ;
      RECT 34.275 2.272 34.485 2.565 ;
      RECT 34.275 2.27 34.475 2.565 ;
      RECT 34.285 2.257 34.475 2.565 ;
      RECT 34.285 2.255 34.4 2.565 ;
      RECT 33.76 2.38 33.935 2.66 ;
      RECT 33.755 2.38 33.935 2.658 ;
      RECT 33.755 2.38 33.95 2.655 ;
      RECT 33.745 2.38 33.95 2.653 ;
      RECT 33.69 2.38 33.95 2.64 ;
      RECT 33.69 2.455 33.955 2.618 ;
      RECT 33.235 2.392 33.255 2.635 ;
      RECT 33.235 2.392 33.295 2.634 ;
      RECT 33.23 2.394 33.295 2.633 ;
      RECT 33.23 2.394 33.381 2.632 ;
      RECT 33.23 2.394 33.45 2.631 ;
      RECT 33.23 2.394 33.47 2.623 ;
      RECT 33.21 2.397 33.47 2.621 ;
      RECT 33.195 2.407 33.47 2.606 ;
      RECT 33.195 2.407 33.485 2.605 ;
      RECT 33.19 2.416 33.485 2.597 ;
      RECT 33.19 2.416 33.49 2.593 ;
      RECT 33.295 2.33 33.555 2.59 ;
      RECT 33.185 2.418 33.555 2.475 ;
      RECT 33.255 2.385 33.555 2.59 ;
      RECT 33.22 3.578 33.225 3.785 ;
      RECT 33.17 3.572 33.22 3.784 ;
      RECT 33.137 3.586 33.23 3.783 ;
      RECT 33.051 3.586 33.23 3.782 ;
      RECT 32.965 3.586 33.23 3.781 ;
      RECT 32.965 3.685 33.235 3.778 ;
      RECT 32.96 3.685 33.235 3.773 ;
      RECT 32.955 3.685 33.235 3.755 ;
      RECT 32.95 3.685 33.235 3.738 ;
      RECT 32.91 3.47 33.17 3.73 ;
      RECT 32.37 2.62 32.456 3.034 ;
      RECT 32.37 2.62 32.495 3.031 ;
      RECT 32.37 2.62 32.515 3.021 ;
      RECT 32.325 2.62 32.515 3.018 ;
      RECT 32.325 2.772 32.525 3.008 ;
      RECT 32.325 2.793 32.53 3.002 ;
      RECT 32.325 2.811 32.535 2.998 ;
      RECT 32.325 2.831 32.545 2.993 ;
      RECT 32.3 2.831 32.545 2.99 ;
      RECT 32.29 2.831 32.545 2.968 ;
      RECT 32.29 2.847 32.55 2.938 ;
      RECT 32.255 2.62 32.515 2.925 ;
      RECT 32.255 2.859 32.555 2.88 ;
      RECT 29.92 2.365 30.21 2.595 ;
      RECT 29.98 0.885 30.15 2.595 ;
      RECT 29.95 1.095 30.29 1.445 ;
      RECT 29.92 0.885 30.21 1.115 ;
      RECT 29.92 7.765 30.21 7.995 ;
      RECT 29.98 6.285 30.15 7.995 ;
      RECT 29.92 6.285 30.21 6.515 ;
      RECT 29.51 2.735 29.84 2.965 ;
      RECT 29.51 2.765 30.01 2.935 ;
      RECT 29.51 2.395 29.7 2.965 ;
      RECT 28.93 2.365 29.22 2.595 ;
      RECT 28.93 2.395 29.7 2.565 ;
      RECT 28.99 0.885 29.16 2.595 ;
      RECT 28.93 0.885 29.22 1.115 ;
      RECT 28.93 7.765 29.22 7.995 ;
      RECT 28.99 6.285 29.16 7.995 ;
      RECT 28.93 6.285 29.22 6.515 ;
      RECT 28.93 6.325 29.78 6.485 ;
      RECT 29.61 5.915 29.78 6.485 ;
      RECT 28.93 6.32 29.32 6.485 ;
      RECT 29.55 5.915 29.84 6.145 ;
      RECT 29.55 5.945 30.01 6.115 ;
      RECT 28.56 2.735 28.85 2.965 ;
      RECT 28.56 2.765 29.02 2.935 ;
      RECT 28.62 1.655 28.785 2.965 ;
      RECT 27.135 1.625 27.425 1.855 ;
      RECT 27.135 1.655 28.785 1.825 ;
      RECT 27.195 0.885 27.365 1.855 ;
      RECT 27.135 0.885 27.425 1.115 ;
      RECT 27.135 7.765 27.425 7.995 ;
      RECT 27.195 7.025 27.365 7.995 ;
      RECT 27.195 7.12 28.785 7.29 ;
      RECT 28.615 5.915 28.785 7.29 ;
      RECT 27.135 7.025 27.425 7.255 ;
      RECT 28.56 5.915 28.85 6.145 ;
      RECT 28.56 5.945 29.02 6.115 ;
      RECT 27.565 1.965 27.915 2.315 ;
      RECT 27.395 2.025 27.915 2.195 ;
      RECT 27.59 6.655 27.915 6.98 ;
      RECT 27.565 6.655 27.915 6.885 ;
      RECT 27.395 6.685 27.915 6.855 ;
      RECT 25.185 2.705 25.525 3.055 ;
      RECT 25.275 2.395 25.445 3.055 ;
      RECT 26.79 2.365 27.11 2.685 ;
      RECT 26.76 2.365 27.11 2.595 ;
      RECT 25.275 2.395 27.11 2.565 ;
      RECT 26.79 6.28 27.11 6.605 ;
      RECT 26.76 6.285 27.11 6.515 ;
      RECT 26.59 6.315 27.11 6.485 ;
      RECT 25.745 2.705 26.085 3.055 ;
      RECT 25.745 2.765 26.225 2.935 ;
      RECT 25.74 5.86 26.08 6.21 ;
      RECT 25.74 5.945 26.225 6.115 ;
      RECT 22.48 2.985 22.63 3.26 ;
      RECT 23.02 2.065 23.025 2.285 ;
      RECT 24.17 2.265 24.185 2.463 ;
      RECT 24.135 2.257 24.17 2.47 ;
      RECT 24.105 2.25 24.135 2.47 ;
      RECT 24.05 2.215 24.105 2.47 ;
      RECT 23.985 2.152 24.05 2.47 ;
      RECT 23.98 2.117 23.985 2.468 ;
      RECT 23.975 2.112 23.98 2.46 ;
      RECT 23.97 2.107 23.975 2.446 ;
      RECT 23.965 2.104 23.97 2.439 ;
      RECT 23.92 2.094 23.965 2.39 ;
      RECT 23.9 2.081 23.92 2.325 ;
      RECT 23.895 2.076 23.9 2.298 ;
      RECT 23.89 2.075 23.895 2.291 ;
      RECT 23.885 2.074 23.89 2.284 ;
      RECT 23.8 2.059 23.885 2.23 ;
      RECT 23.77 2.04 23.8 2.18 ;
      RECT 23.69 2.023 23.77 2.165 ;
      RECT 23.655 2.01 23.69 2.15 ;
      RECT 23.647 2.01 23.655 2.145 ;
      RECT 23.561 2.011 23.647 2.145 ;
      RECT 23.475 2.013 23.561 2.145 ;
      RECT 23.45 2.014 23.475 2.149 ;
      RECT 23.375 2.02 23.45 2.164 ;
      RECT 23.292 2.032 23.375 2.188 ;
      RECT 23.206 2.045 23.292 2.214 ;
      RECT 23.12 2.058 23.206 2.24 ;
      RECT 23.085 2.067 23.12 2.259 ;
      RECT 23.035 2.067 23.085 2.272 ;
      RECT 23.025 2.065 23.035 2.283 ;
      RECT 23.01 2.062 23.02 2.285 ;
      RECT 22.995 2.054 23.01 2.293 ;
      RECT 22.98 2.046 22.995 2.313 ;
      RECT 22.975 2.041 22.98 2.37 ;
      RECT 22.96 2.036 22.975 2.443 ;
      RECT 22.955 2.031 22.96 2.485 ;
      RECT 22.95 2.029 22.955 2.513 ;
      RECT 22.945 2.027 22.95 2.535 ;
      RECT 22.935 2.023 22.945 2.578 ;
      RECT 22.93 2.02 22.935 2.603 ;
      RECT 22.925 2.018 22.93 2.623 ;
      RECT 22.92 2.016 22.925 2.647 ;
      RECT 22.915 2.012 22.92 2.67 ;
      RECT 22.91 2.008 22.915 2.693 ;
      RECT 22.875 1.998 22.91 2.8 ;
      RECT 22.87 1.988 22.875 2.898 ;
      RECT 22.865 1.986 22.87 2.925 ;
      RECT 22.86 1.985 22.865 2.945 ;
      RECT 22.855 1.977 22.86 2.965 ;
      RECT 22.85 1.972 22.855 3 ;
      RECT 22.845 1.97 22.85 3.018 ;
      RECT 22.84 1.97 22.845 3.043 ;
      RECT 22.835 1.97 22.84 3.065 ;
      RECT 22.8 1.97 22.835 3.108 ;
      RECT 22.775 1.97 22.8 3.137 ;
      RECT 22.765 1.97 22.775 2.323 ;
      RECT 22.768 2.38 22.775 3.147 ;
      RECT 22.765 2.437 22.768 3.15 ;
      RECT 22.76 1.97 22.765 2.295 ;
      RECT 22.76 2.487 22.765 3.153 ;
      RECT 22.75 1.97 22.76 2.285 ;
      RECT 22.755 2.54 22.76 3.156 ;
      RECT 22.75 2.625 22.755 3.16 ;
      RECT 22.74 1.97 22.75 2.273 ;
      RECT 22.745 2.672 22.75 3.164 ;
      RECT 22.74 2.747 22.745 3.168 ;
      RECT 22.705 1.97 22.74 2.248 ;
      RECT 22.73 2.83 22.74 3.173 ;
      RECT 22.72 2.897 22.73 3.18 ;
      RECT 22.715 2.925 22.72 3.185 ;
      RECT 22.705 2.938 22.715 3.191 ;
      RECT 22.66 1.97 22.705 2.205 ;
      RECT 22.7 2.943 22.705 3.198 ;
      RECT 22.66 2.96 22.7 3.26 ;
      RECT 22.655 1.972 22.66 2.178 ;
      RECT 22.63 2.98 22.66 3.26 ;
      RECT 22.65 1.977 22.655 2.15 ;
      RECT 22.44 2.989 22.48 3.26 ;
      RECT 22.415 2.997 22.44 3.23 ;
      RECT 22.37 3.005 22.415 3.23 ;
      RECT 22.355 3.01 22.37 3.225 ;
      RECT 22.345 3.01 22.355 3.219 ;
      RECT 22.335 3.017 22.345 3.216 ;
      RECT 22.33 3.055 22.335 3.205 ;
      RECT 22.325 3.117 22.33 3.183 ;
      RECT 23.595 2.992 23.78 3.215 ;
      RECT 23.595 3.007 23.785 3.211 ;
      RECT 23.585 2.28 23.67 3.21 ;
      RECT 23.585 3.007 23.79 3.204 ;
      RECT 23.58 3.015 23.79 3.203 ;
      RECT 23.785 2.735 24.105 3.055 ;
      RECT 23.58 2.907 23.75 2.998 ;
      RECT 23.575 2.907 23.75 2.98 ;
      RECT 23.565 2.715 23.7 2.955 ;
      RECT 23.56 2.715 23.7 2.9 ;
      RECT 23.52 2.295 23.69 2.8 ;
      RECT 23.505 2.295 23.69 2.67 ;
      RECT 23.5 2.295 23.69 2.623 ;
      RECT 23.495 2.295 23.69 2.603 ;
      RECT 23.49 2.295 23.69 2.578 ;
      RECT 23.46 2.295 23.72 2.555 ;
      RECT 23.47 2.292 23.68 2.555 ;
      RECT 23.595 2.287 23.68 3.215 ;
      RECT 23.48 2.28 23.67 2.555 ;
      RECT 23.475 2.285 23.67 2.555 ;
      RECT 22.305 2.497 22.49 2.71 ;
      RECT 22.305 2.505 22.5 2.703 ;
      RECT 22.285 2.505 22.5 2.7 ;
      RECT 22.28 2.505 22.5 2.685 ;
      RECT 22.21 2.42 22.47 2.68 ;
      RECT 22.21 2.565 22.505 2.593 ;
      RECT 21.865 3.02 22.125 3.28 ;
      RECT 21.89 2.965 22.085 3.28 ;
      RECT 21.885 2.714 22.065 3.008 ;
      RECT 21.885 2.72 22.075 3.008 ;
      RECT 21.865 2.722 22.075 2.953 ;
      RECT 21.86 2.732 22.075 2.82 ;
      RECT 21.89 2.712 22.065 3.28 ;
      RECT 21.976 2.71 22.065 3.28 ;
      RECT 21.835 1.93 21.87 2.3 ;
      RECT 21.625 2.04 21.63 2.3 ;
      RECT 21.87 1.937 21.885 2.3 ;
      RECT 21.76 1.93 21.835 2.378 ;
      RECT 21.75 1.93 21.76 2.463 ;
      RECT 21.725 1.93 21.75 2.498 ;
      RECT 21.685 1.93 21.725 2.566 ;
      RECT 21.675 1.937 21.685 2.618 ;
      RECT 21.645 2.04 21.675 2.659 ;
      RECT 21.64 2.04 21.645 2.698 ;
      RECT 21.63 2.04 21.64 2.718 ;
      RECT 21.625 2.335 21.63 2.755 ;
      RECT 21.62 2.352 21.625 2.775 ;
      RECT 21.605 2.415 21.62 2.815 ;
      RECT 21.6 2.458 21.605 2.85 ;
      RECT 21.595 2.466 21.6 2.863 ;
      RECT 21.585 2.48 21.595 2.885 ;
      RECT 21.56 2.515 21.585 2.95 ;
      RECT 21.55 2.55 21.56 3.013 ;
      RECT 21.53 2.58 21.55 3.074 ;
      RECT 21.515 2.616 21.53 3.141 ;
      RECT 21.505 2.644 21.515 3.18 ;
      RECT 21.495 2.666 21.505 3.2 ;
      RECT 21.49 2.676 21.495 3.211 ;
      RECT 21.485 2.685 21.49 3.214 ;
      RECT 21.475 2.703 21.485 3.218 ;
      RECT 21.465 2.721 21.475 3.219 ;
      RECT 21.44 2.76 21.465 3.216 ;
      RECT 21.42 2.802 21.44 3.213 ;
      RECT 21.405 2.84 21.42 3.212 ;
      RECT 21.37 2.875 21.405 3.209 ;
      RECT 21.365 2.897 21.37 3.207 ;
      RECT 21.3 2.937 21.365 3.204 ;
      RECT 21.295 2.977 21.3 3.2 ;
      RECT 21.28 2.987 21.295 3.191 ;
      RECT 21.27 3.107 21.28 3.176 ;
      RECT 21.75 3.52 21.76 3.78 ;
      RECT 21.75 3.523 21.77 3.779 ;
      RECT 21.74 3.513 21.75 3.778 ;
      RECT 21.73 3.528 21.81 3.774 ;
      RECT 21.715 3.507 21.73 3.772 ;
      RECT 21.69 3.532 21.815 3.768 ;
      RECT 21.675 3.492 21.69 3.763 ;
      RECT 21.675 3.534 21.825 3.762 ;
      RECT 21.675 3.542 21.84 3.755 ;
      RECT 21.615 3.479 21.675 3.745 ;
      RECT 21.605 3.466 21.615 3.727 ;
      RECT 21.58 3.456 21.605 3.717 ;
      RECT 21.575 3.446 21.58 3.709 ;
      RECT 21.51 3.542 21.84 3.691 ;
      RECT 21.425 3.542 21.84 3.653 ;
      RECT 21.315 3.37 21.575 3.63 ;
      RECT 21.69 3.5 21.715 3.768 ;
      RECT 21.73 3.51 21.74 3.774 ;
      RECT 21.315 3.518 21.755 3.63 ;
      RECT 20.53 3.275 20.56 3.575 ;
      RECT 20.305 3.26 20.31 3.535 ;
      RECT 20.105 3.26 20.26 3.52 ;
      RECT 21.405 1.975 21.435 2.235 ;
      RECT 21.395 1.975 21.405 2.343 ;
      RECT 21.375 1.975 21.395 2.353 ;
      RECT 21.36 1.975 21.375 2.365 ;
      RECT 21.305 1.975 21.36 2.415 ;
      RECT 21.29 1.975 21.305 2.463 ;
      RECT 21.26 1.975 21.29 2.498 ;
      RECT 21.205 1.975 21.26 2.56 ;
      RECT 21.185 1.975 21.205 2.628 ;
      RECT 21.18 1.975 21.185 2.658 ;
      RECT 21.175 1.975 21.18 2.67 ;
      RECT 21.17 2.092 21.175 2.688 ;
      RECT 21.15 2.11 21.17 2.713 ;
      RECT 21.13 2.137 21.15 2.763 ;
      RECT 21.125 2.157 21.13 2.794 ;
      RECT 21.12 2.165 21.125 2.811 ;
      RECT 21.105 2.191 21.12 2.84 ;
      RECT 21.09 2.233 21.105 2.875 ;
      RECT 21.085 2.262 21.09 2.898 ;
      RECT 21.08 2.277 21.085 2.911 ;
      RECT 21.075 2.3 21.08 2.922 ;
      RECT 21.065 2.32 21.075 2.94 ;
      RECT 21.055 2.35 21.065 2.963 ;
      RECT 21.05 2.372 21.055 2.983 ;
      RECT 21.045 2.387 21.05 2.998 ;
      RECT 21.03 2.417 21.045 3.025 ;
      RECT 21.025 2.447 21.03 3.051 ;
      RECT 21.02 2.465 21.025 3.063 ;
      RECT 21.01 2.495 21.02 3.082 ;
      RECT 21 2.52 21.01 3.107 ;
      RECT 20.995 2.54 21 3.126 ;
      RECT 20.99 2.557 20.995 3.139 ;
      RECT 20.98 2.583 20.99 3.158 ;
      RECT 20.97 2.621 20.98 3.185 ;
      RECT 20.965 2.647 20.97 3.205 ;
      RECT 20.96 2.657 20.965 3.215 ;
      RECT 20.955 2.67 20.96 3.23 ;
      RECT 20.95 2.685 20.955 3.24 ;
      RECT 20.945 2.707 20.95 3.255 ;
      RECT 20.94 2.725 20.945 3.266 ;
      RECT 20.935 2.735 20.94 3.277 ;
      RECT 20.93 2.743 20.935 3.289 ;
      RECT 20.925 2.751 20.93 3.3 ;
      RECT 20.92 2.777 20.925 3.313 ;
      RECT 20.91 2.805 20.92 3.326 ;
      RECT 20.905 2.835 20.91 3.335 ;
      RECT 20.9 2.85 20.905 3.342 ;
      RECT 20.885 2.875 20.9 3.349 ;
      RECT 20.88 2.897 20.885 3.355 ;
      RECT 20.875 2.922 20.88 3.358 ;
      RECT 20.866 2.95 20.875 3.362 ;
      RECT 20.86 2.967 20.866 3.367 ;
      RECT 20.855 2.985 20.86 3.371 ;
      RECT 20.85 2.997 20.855 3.374 ;
      RECT 20.845 3.018 20.85 3.378 ;
      RECT 20.84 3.036 20.845 3.381 ;
      RECT 20.835 3.05 20.84 3.384 ;
      RECT 20.83 3.067 20.835 3.387 ;
      RECT 20.825 3.08 20.83 3.39 ;
      RECT 20.8 3.117 20.825 3.398 ;
      RECT 20.795 3.162 20.8 3.407 ;
      RECT 20.79 3.19 20.795 3.41 ;
      RECT 20.78 3.21 20.79 3.414 ;
      RECT 20.775 3.23 20.78 3.419 ;
      RECT 20.77 3.245 20.775 3.422 ;
      RECT 20.75 3.255 20.77 3.429 ;
      RECT 20.685 3.262 20.75 3.455 ;
      RECT 20.65 3.265 20.685 3.483 ;
      RECT 20.635 3.268 20.65 3.498 ;
      RECT 20.625 3.269 20.635 3.513 ;
      RECT 20.615 3.27 20.625 3.53 ;
      RECT 20.61 3.27 20.615 3.545 ;
      RECT 20.605 3.27 20.61 3.553 ;
      RECT 20.59 3.271 20.605 3.568 ;
      RECT 20.56 3.273 20.59 3.575 ;
      RECT 20.45 3.28 20.53 3.575 ;
      RECT 20.405 3.285 20.45 3.575 ;
      RECT 20.395 3.286 20.405 3.565 ;
      RECT 20.385 3.287 20.395 3.558 ;
      RECT 20.365 3.289 20.385 3.553 ;
      RECT 20.355 3.26 20.365 3.548 ;
      RECT 20.31 3.26 20.355 3.54 ;
      RECT 20.28 3.26 20.305 3.53 ;
      RECT 20.26 3.26 20.28 3.523 ;
      RECT 20.54 2.06 20.8 2.32 ;
      RECT 20.42 2.075 20.43 2.24 ;
      RECT 20.405 2.075 20.41 2.235 ;
      RECT 17.77 1.915 17.955 2.205 ;
      RECT 19.585 2.04 19.6 2.195 ;
      RECT 17.735 1.915 17.76 2.175 ;
      RECT 20.15 1.965 20.155 2.107 ;
      RECT 20.065 1.96 20.09 2.1 ;
      RECT 20.465 2.077 20.54 2.27 ;
      RECT 20.45 2.075 20.465 2.253 ;
      RECT 20.43 2.075 20.45 2.245 ;
      RECT 20.41 2.075 20.42 2.238 ;
      RECT 20.365 2.07 20.405 2.228 ;
      RECT 20.325 2.045 20.365 2.213 ;
      RECT 20.31 2.02 20.325 2.203 ;
      RECT 20.305 2.014 20.31 2.201 ;
      RECT 20.27 2.006 20.305 2.184 ;
      RECT 20.265 1.999 20.27 2.172 ;
      RECT 20.245 1.994 20.265 2.16 ;
      RECT 20.235 1.988 20.245 2.145 ;
      RECT 20.215 1.983 20.235 2.13 ;
      RECT 20.205 1.978 20.215 2.123 ;
      RECT 20.2 1.976 20.205 2.118 ;
      RECT 20.195 1.975 20.2 2.115 ;
      RECT 20.155 1.97 20.195 2.111 ;
      RECT 20.135 1.964 20.15 2.106 ;
      RECT 20.1 1.961 20.135 2.103 ;
      RECT 20.09 1.96 20.1 2.101 ;
      RECT 20.03 1.96 20.065 2.098 ;
      RECT 19.985 1.96 20.03 2.098 ;
      RECT 19.935 1.96 19.985 2.101 ;
      RECT 19.92 1.962 19.935 2.103 ;
      RECT 19.905 1.965 19.92 2.104 ;
      RECT 19.895 1.97 19.905 2.105 ;
      RECT 19.865 1.975 19.895 2.11 ;
      RECT 19.855 1.981 19.865 2.118 ;
      RECT 19.845 1.983 19.855 2.122 ;
      RECT 19.835 1.987 19.845 2.126 ;
      RECT 19.81 1.993 19.835 2.134 ;
      RECT 19.8 1.998 19.81 2.142 ;
      RECT 19.785 2.002 19.8 2.146 ;
      RECT 19.75 2.008 19.785 2.154 ;
      RECT 19.73 2.013 19.75 2.164 ;
      RECT 19.7 2.02 19.73 2.173 ;
      RECT 19.655 2.029 19.7 2.187 ;
      RECT 19.65 2.034 19.655 2.198 ;
      RECT 19.63 2.037 19.65 2.199 ;
      RECT 19.6 2.04 19.63 2.197 ;
      RECT 19.565 2.04 19.585 2.193 ;
      RECT 19.495 2.04 19.565 2.184 ;
      RECT 19.48 2.037 19.495 2.176 ;
      RECT 19.44 2.03 19.48 2.171 ;
      RECT 19.415 2.02 19.44 2.164 ;
      RECT 19.41 2.014 19.415 2.161 ;
      RECT 19.37 2.008 19.41 2.158 ;
      RECT 19.355 2.001 19.37 2.153 ;
      RECT 19.335 1.997 19.355 2.148 ;
      RECT 19.32 1.992 19.335 2.144 ;
      RECT 19.305 1.987 19.32 2.142 ;
      RECT 19.29 1.983 19.305 2.141 ;
      RECT 19.275 1.981 19.29 2.137 ;
      RECT 19.265 1.979 19.275 2.132 ;
      RECT 19.25 1.976 19.265 2.128 ;
      RECT 19.24 1.974 19.25 2.123 ;
      RECT 19.22 1.971 19.24 2.119 ;
      RECT 19.175 1.97 19.22 2.117 ;
      RECT 19.115 1.972 19.175 2.118 ;
      RECT 19.095 1.974 19.115 2.12 ;
      RECT 19.065 1.977 19.095 2.121 ;
      RECT 19.015 1.982 19.065 2.123 ;
      RECT 19.01 1.985 19.015 2.125 ;
      RECT 19 1.987 19.01 2.128 ;
      RECT 18.995 1.989 19 2.131 ;
      RECT 18.945 1.992 18.995 2.138 ;
      RECT 18.925 1.996 18.945 2.15 ;
      RECT 18.915 1.999 18.925 2.156 ;
      RECT 18.905 2 18.915 2.159 ;
      RECT 18.866 2.003 18.905 2.161 ;
      RECT 18.78 2.01 18.866 2.164 ;
      RECT 18.706 2.02 18.78 2.168 ;
      RECT 18.62 2.031 18.706 2.173 ;
      RECT 18.605 2.038 18.62 2.175 ;
      RECT 18.55 2.042 18.605 2.176 ;
      RECT 18.536 2.045 18.55 2.178 ;
      RECT 18.45 2.045 18.536 2.18 ;
      RECT 18.41 2.042 18.45 2.183 ;
      RECT 18.386 2.038 18.41 2.185 ;
      RECT 18.3 2.028 18.386 2.188 ;
      RECT 18.27 2.017 18.3 2.189 ;
      RECT 18.251 2.013 18.27 2.188 ;
      RECT 18.165 2.006 18.251 2.185 ;
      RECT 18.105 1.995 18.165 2.182 ;
      RECT 18.085 1.987 18.105 2.18 ;
      RECT 18.05 1.982 18.085 2.179 ;
      RECT 18.025 1.977 18.05 2.178 ;
      RECT 17.995 1.972 18.025 2.177 ;
      RECT 17.97 1.915 17.995 2.176 ;
      RECT 17.955 1.915 17.97 2.2 ;
      RECT 17.76 1.915 17.77 2.2 ;
      RECT 19.535 2.935 19.54 3.075 ;
      RECT 19.195 2.935 19.23 3.073 ;
      RECT 18.77 2.92 18.785 3.065 ;
      RECT 20.6 2.7 20.69 2.96 ;
      RECT 20.43 2.565 20.53 2.96 ;
      RECT 17.465 2.54 17.545 2.75 ;
      RECT 20.555 2.677 20.6 2.96 ;
      RECT 20.545 2.647 20.555 2.96 ;
      RECT 20.53 2.57 20.545 2.96 ;
      RECT 20.345 2.565 20.43 2.925 ;
      RECT 20.34 2.567 20.345 2.92 ;
      RECT 20.335 2.572 20.34 2.92 ;
      RECT 20.3 2.672 20.335 2.92 ;
      RECT 20.29 2.7 20.3 2.92 ;
      RECT 20.28 2.715 20.29 2.92 ;
      RECT 20.27 2.727 20.28 2.92 ;
      RECT 20.265 2.737 20.27 2.92 ;
      RECT 20.25 2.747 20.265 2.922 ;
      RECT 20.245 2.762 20.25 2.924 ;
      RECT 20.23 2.775 20.245 2.926 ;
      RECT 20.225 2.79 20.23 2.929 ;
      RECT 20.205 2.8 20.225 2.933 ;
      RECT 20.19 2.81 20.205 2.936 ;
      RECT 20.155 2.817 20.19 2.941 ;
      RECT 20.111 2.824 20.155 2.949 ;
      RECT 20.025 2.836 20.111 2.962 ;
      RECT 20 2.847 20.025 2.973 ;
      RECT 19.97 2.852 20 2.978 ;
      RECT 19.935 2.857 19.97 2.986 ;
      RECT 19.905 2.862 19.935 2.993 ;
      RECT 19.88 2.867 19.905 2.998 ;
      RECT 19.815 2.874 19.88 3.007 ;
      RECT 19.745 2.887 19.815 3.023 ;
      RECT 19.715 2.897 19.745 3.035 ;
      RECT 19.69 2.902 19.715 3.042 ;
      RECT 19.635 2.909 19.69 3.05 ;
      RECT 19.63 2.916 19.635 3.055 ;
      RECT 19.625 2.918 19.63 3.056 ;
      RECT 19.61 2.92 19.625 3.058 ;
      RECT 19.605 2.92 19.61 3.061 ;
      RECT 19.54 2.927 19.605 3.068 ;
      RECT 19.505 2.937 19.535 3.078 ;
      RECT 19.488 2.94 19.505 3.08 ;
      RECT 19.402 2.939 19.488 3.079 ;
      RECT 19.316 2.937 19.402 3.076 ;
      RECT 19.23 2.936 19.316 3.074 ;
      RECT 19.129 2.934 19.195 3.073 ;
      RECT 19.043 2.931 19.129 3.071 ;
      RECT 18.957 2.927 19.043 3.069 ;
      RECT 18.871 2.924 18.957 3.068 ;
      RECT 18.785 2.921 18.871 3.066 ;
      RECT 18.685 2.92 18.77 3.063 ;
      RECT 18.635 2.918 18.685 3.061 ;
      RECT 18.615 2.915 18.635 3.059 ;
      RECT 18.595 2.913 18.615 3.056 ;
      RECT 18.57 2.909 18.595 3.053 ;
      RECT 18.525 2.903 18.57 3.048 ;
      RECT 18.485 2.897 18.525 3.04 ;
      RECT 18.46 2.892 18.485 3.033 ;
      RECT 18.405 2.885 18.46 3.025 ;
      RECT 18.381 2.878 18.405 3.018 ;
      RECT 18.295 2.869 18.381 3.008 ;
      RECT 18.265 2.861 18.295 2.998 ;
      RECT 18.235 2.857 18.265 2.993 ;
      RECT 18.23 2.854 18.235 2.99 ;
      RECT 18.225 2.853 18.23 2.99 ;
      RECT 18.15 2.846 18.225 2.983 ;
      RECT 18.111 2.837 18.15 2.972 ;
      RECT 18.025 2.827 18.111 2.96 ;
      RECT 17.985 2.817 18.025 2.948 ;
      RECT 17.946 2.812 17.985 2.941 ;
      RECT 17.86 2.802 17.946 2.93 ;
      RECT 17.82 2.79 17.86 2.919 ;
      RECT 17.785 2.775 17.82 2.912 ;
      RECT 17.775 2.765 17.785 2.909 ;
      RECT 17.755 2.75 17.775 2.907 ;
      RECT 17.725 2.72 17.755 2.903 ;
      RECT 17.715 2.7 17.725 2.898 ;
      RECT 17.71 2.692 17.715 2.895 ;
      RECT 17.705 2.685 17.71 2.893 ;
      RECT 17.69 2.672 17.705 2.886 ;
      RECT 17.685 2.662 17.69 2.878 ;
      RECT 17.68 2.655 17.685 2.873 ;
      RECT 17.675 2.65 17.68 2.869 ;
      RECT 17.66 2.637 17.675 2.861 ;
      RECT 17.655 2.547 17.66 2.85 ;
      RECT 17.65 2.542 17.655 2.843 ;
      RECT 17.575 2.54 17.65 2.803 ;
      RECT 17.545 2.54 17.575 2.758 ;
      RECT 17.45 2.545 17.465 2.745 ;
      RECT 19.935 2.25 20.195 2.51 ;
      RECT 19.92 2.238 20.1 2.475 ;
      RECT 19.915 2.239 20.1 2.473 ;
      RECT 19.9 2.243 20.11 2.463 ;
      RECT 19.895 2.248 20.115 2.433 ;
      RECT 19.9 2.245 20.115 2.463 ;
      RECT 19.915 2.24 20.11 2.473 ;
      RECT 19.935 2.237 20.1 2.51 ;
      RECT 19.935 2.236 20.09 2.51 ;
      RECT 19.96 2.235 20.09 2.51 ;
      RECT 19.52 2.48 19.78 2.74 ;
      RECT 19.395 2.525 19.78 2.735 ;
      RECT 19.385 2.53 19.78 2.73 ;
      RECT 19.4 3.47 19.415 3.78 ;
      RECT 17.995 3.24 18.005 3.37 ;
      RECT 17.775 3.235 17.88 3.37 ;
      RECT 17.69 3.24 17.74 3.37 ;
      RECT 16.24 1.975 16.245 3.08 ;
      RECT 19.495 3.562 19.5 3.698 ;
      RECT 19.49 3.557 19.495 3.758 ;
      RECT 19.485 3.555 19.49 3.771 ;
      RECT 19.47 3.552 19.485 3.773 ;
      RECT 19.465 3.547 19.47 3.775 ;
      RECT 19.46 3.543 19.465 3.778 ;
      RECT 19.445 3.538 19.46 3.78 ;
      RECT 19.415 3.53 19.445 3.78 ;
      RECT 19.376 3.47 19.4 3.78 ;
      RECT 19.29 3.47 19.376 3.777 ;
      RECT 19.26 3.47 19.29 3.77 ;
      RECT 19.235 3.47 19.26 3.763 ;
      RECT 19.21 3.47 19.235 3.755 ;
      RECT 19.195 3.47 19.21 3.748 ;
      RECT 19.17 3.47 19.195 3.74 ;
      RECT 19.155 3.47 19.17 3.733 ;
      RECT 19.115 3.48 19.155 3.722 ;
      RECT 19.105 3.475 19.115 3.712 ;
      RECT 19.101 3.474 19.105 3.709 ;
      RECT 19.015 3.466 19.101 3.692 ;
      RECT 18.982 3.455 19.015 3.669 ;
      RECT 18.896 3.444 18.982 3.647 ;
      RECT 18.81 3.428 18.896 3.616 ;
      RECT 18.74 3.413 18.81 3.588 ;
      RECT 18.73 3.406 18.74 3.575 ;
      RECT 18.7 3.403 18.73 3.565 ;
      RECT 18.675 3.399 18.7 3.558 ;
      RECT 18.66 3.396 18.675 3.553 ;
      RECT 18.655 3.395 18.66 3.548 ;
      RECT 18.625 3.39 18.655 3.541 ;
      RECT 18.62 3.385 18.625 3.536 ;
      RECT 18.605 3.382 18.62 3.531 ;
      RECT 18.6 3.377 18.605 3.526 ;
      RECT 18.58 3.372 18.6 3.523 ;
      RECT 18.565 3.367 18.58 3.515 ;
      RECT 18.55 3.361 18.565 3.51 ;
      RECT 18.52 3.352 18.55 3.503 ;
      RECT 18.515 3.345 18.52 3.495 ;
      RECT 18.51 3.343 18.515 3.493 ;
      RECT 18.505 3.342 18.51 3.49 ;
      RECT 18.465 3.335 18.505 3.483 ;
      RECT 18.451 3.325 18.465 3.473 ;
      RECT 18.4 3.314 18.451 3.461 ;
      RECT 18.375 3.3 18.4 3.447 ;
      RECT 18.35 3.289 18.375 3.439 ;
      RECT 18.33 3.278 18.35 3.433 ;
      RECT 18.32 3.272 18.33 3.428 ;
      RECT 18.315 3.27 18.32 3.424 ;
      RECT 18.295 3.265 18.315 3.419 ;
      RECT 18.265 3.255 18.295 3.409 ;
      RECT 18.26 3.247 18.265 3.402 ;
      RECT 18.245 3.245 18.26 3.398 ;
      RECT 18.225 3.245 18.245 3.393 ;
      RECT 18.22 3.244 18.225 3.391 ;
      RECT 18.215 3.244 18.22 3.388 ;
      RECT 18.175 3.243 18.215 3.383 ;
      RECT 18.15 3.242 18.175 3.378 ;
      RECT 18.09 3.241 18.15 3.375 ;
      RECT 18.005 3.24 18.09 3.373 ;
      RECT 17.966 3.239 17.995 3.37 ;
      RECT 17.88 3.237 17.966 3.37 ;
      RECT 17.74 3.237 17.775 3.37 ;
      RECT 17.65 3.241 17.69 3.373 ;
      RECT 17.635 3.244 17.65 3.38 ;
      RECT 17.625 3.245 17.635 3.387 ;
      RECT 17.6 3.248 17.625 3.392 ;
      RECT 17.595 3.25 17.6 3.395 ;
      RECT 17.545 3.252 17.595 3.396 ;
      RECT 17.506 3.256 17.545 3.398 ;
      RECT 17.42 3.258 17.506 3.401 ;
      RECT 17.402 3.26 17.42 3.403 ;
      RECT 17.316 3.263 17.402 3.405 ;
      RECT 17.23 3.267 17.316 3.408 ;
      RECT 17.193 3.271 17.23 3.411 ;
      RECT 17.107 3.274 17.193 3.414 ;
      RECT 17.021 3.278 17.107 3.417 ;
      RECT 16.935 3.283 17.021 3.421 ;
      RECT 16.915 3.285 16.935 3.424 ;
      RECT 16.895 3.284 16.915 3.425 ;
      RECT 16.846 3.281 16.895 3.426 ;
      RECT 16.76 3.276 16.846 3.429 ;
      RECT 16.71 3.271 16.76 3.431 ;
      RECT 16.686 3.269 16.71 3.432 ;
      RECT 16.6 3.264 16.686 3.434 ;
      RECT 16.575 3.26 16.6 3.433 ;
      RECT 16.565 3.257 16.575 3.431 ;
      RECT 16.555 3.25 16.565 3.428 ;
      RECT 16.55 3.23 16.555 3.423 ;
      RECT 16.54 3.2 16.55 3.418 ;
      RECT 16.525 3.07 16.54 3.409 ;
      RECT 16.52 3.062 16.525 3.402 ;
      RECT 16.5 3.055 16.52 3.394 ;
      RECT 16.495 3.037 16.5 3.386 ;
      RECT 16.485 3.017 16.495 3.381 ;
      RECT 16.48 2.99 16.485 3.377 ;
      RECT 16.475 2.967 16.48 3.374 ;
      RECT 16.455 2.925 16.475 3.366 ;
      RECT 16.42 2.84 16.455 3.35 ;
      RECT 16.415 2.772 16.42 3.338 ;
      RECT 16.4 2.742 16.415 3.332 ;
      RECT 16.395 1.987 16.4 2.233 ;
      RECT 16.385 2.712 16.4 3.323 ;
      RECT 16.39 1.982 16.395 2.265 ;
      RECT 16.385 1.977 16.39 2.308 ;
      RECT 16.38 1.975 16.385 2.343 ;
      RECT 16.365 2.675 16.385 3.313 ;
      RECT 16.375 1.975 16.38 2.38 ;
      RECT 16.36 1.975 16.375 2.478 ;
      RECT 16.36 2.648 16.365 3.306 ;
      RECT 16.355 1.975 16.36 2.553 ;
      RECT 16.355 2.636 16.36 3.303 ;
      RECT 16.35 1.975 16.355 2.585 ;
      RECT 16.35 2.615 16.355 3.3 ;
      RECT 16.345 1.975 16.35 3.297 ;
      RECT 16.31 1.975 16.345 3.283 ;
      RECT 16.295 1.975 16.31 3.265 ;
      RECT 16.275 1.975 16.295 3.255 ;
      RECT 16.25 1.975 16.275 3.238 ;
      RECT 16.245 1.975 16.25 3.188 ;
      RECT 16.235 1.975 16.24 3.018 ;
      RECT 16.23 1.975 16.235 2.925 ;
      RECT 16.225 1.975 16.23 2.838 ;
      RECT 16.22 1.975 16.225 2.77 ;
      RECT 16.215 1.975 16.22 2.713 ;
      RECT 16.205 1.975 16.215 2.608 ;
      RECT 16.2 1.975 16.205 2.48 ;
      RECT 16.195 1.975 16.2 2.398 ;
      RECT 16.19 1.977 16.195 2.315 ;
      RECT 16.185 1.982 16.19 2.248 ;
      RECT 16.18 1.987 16.185 2.175 ;
      RECT 18.995 2.305 19.255 2.565 ;
      RECT 19.015 2.272 19.225 2.565 ;
      RECT 19.015 2.27 19.215 2.565 ;
      RECT 19.025 2.257 19.215 2.565 ;
      RECT 19.025 2.255 19.14 2.565 ;
      RECT 18.5 2.38 18.675 2.66 ;
      RECT 18.495 2.38 18.675 2.658 ;
      RECT 18.495 2.38 18.69 2.655 ;
      RECT 18.485 2.38 18.69 2.653 ;
      RECT 18.43 2.38 18.69 2.64 ;
      RECT 18.43 2.455 18.695 2.618 ;
      RECT 17.975 2.392 17.995 2.635 ;
      RECT 17.975 2.392 18.035 2.634 ;
      RECT 17.97 2.394 18.035 2.633 ;
      RECT 17.97 2.394 18.121 2.632 ;
      RECT 17.97 2.394 18.19 2.631 ;
      RECT 17.97 2.394 18.21 2.623 ;
      RECT 17.95 2.397 18.21 2.621 ;
      RECT 17.935 2.407 18.21 2.606 ;
      RECT 17.935 2.407 18.225 2.605 ;
      RECT 17.93 2.416 18.225 2.597 ;
      RECT 17.93 2.416 18.23 2.593 ;
      RECT 18.035 2.33 18.295 2.59 ;
      RECT 17.925 2.418 18.295 2.475 ;
      RECT 17.995 2.385 18.295 2.59 ;
      RECT 17.96 3.578 17.965 3.785 ;
      RECT 17.91 3.572 17.96 3.784 ;
      RECT 17.877 3.586 17.97 3.783 ;
      RECT 17.791 3.586 17.97 3.782 ;
      RECT 17.705 3.586 17.97 3.781 ;
      RECT 17.705 3.685 17.975 3.778 ;
      RECT 17.7 3.685 17.975 3.773 ;
      RECT 17.695 3.685 17.975 3.755 ;
      RECT 17.69 3.685 17.975 3.738 ;
      RECT 17.65 3.47 17.91 3.73 ;
      RECT 17.11 2.62 17.196 3.034 ;
      RECT 17.11 2.62 17.235 3.031 ;
      RECT 17.11 2.62 17.255 3.021 ;
      RECT 17.065 2.62 17.255 3.018 ;
      RECT 17.065 2.772 17.265 3.008 ;
      RECT 17.065 2.793 17.27 3.002 ;
      RECT 17.065 2.811 17.275 2.998 ;
      RECT 17.065 2.831 17.285 2.993 ;
      RECT 17.04 2.831 17.285 2.99 ;
      RECT 17.03 2.831 17.285 2.968 ;
      RECT 17.03 2.847 17.29 2.938 ;
      RECT 16.995 2.62 17.255 2.925 ;
      RECT 16.995 2.859 17.295 2.88 ;
      RECT 14.66 2.365 14.95 2.595 ;
      RECT 14.72 0.885 14.89 2.595 ;
      RECT 14.69 1.095 15.03 1.445 ;
      RECT 14.66 0.885 14.95 1.115 ;
      RECT 14.66 7.765 14.95 7.995 ;
      RECT 14.72 6.285 14.89 7.995 ;
      RECT 14.66 6.285 14.95 6.515 ;
      RECT 14.25 2.735 14.58 2.965 ;
      RECT 14.25 2.765 14.75 2.935 ;
      RECT 14.25 2.395 14.44 2.965 ;
      RECT 13.67 2.365 13.96 2.595 ;
      RECT 13.67 2.395 14.44 2.565 ;
      RECT 13.73 0.885 13.9 2.595 ;
      RECT 13.67 0.885 13.96 1.115 ;
      RECT 13.67 7.765 13.96 7.995 ;
      RECT 13.73 6.285 13.9 7.995 ;
      RECT 13.67 6.285 13.96 6.515 ;
      RECT 13.67 6.325 14.52 6.485 ;
      RECT 14.35 5.915 14.52 6.485 ;
      RECT 13.67 6.32 14.06 6.485 ;
      RECT 14.29 5.915 14.58 6.145 ;
      RECT 14.29 5.945 14.75 6.115 ;
      RECT 13.3 2.735 13.59 2.965 ;
      RECT 13.3 2.765 13.76 2.935 ;
      RECT 13.36 1.655 13.525 2.965 ;
      RECT 11.875 1.625 12.165 1.855 ;
      RECT 11.875 1.655 13.525 1.825 ;
      RECT 11.935 0.885 12.105 1.855 ;
      RECT 11.875 0.885 12.165 1.115 ;
      RECT 11.875 7.765 12.165 7.995 ;
      RECT 11.935 7.025 12.105 7.995 ;
      RECT 11.935 7.12 13.525 7.29 ;
      RECT 13.355 5.915 13.525 7.29 ;
      RECT 11.875 7.025 12.165 7.255 ;
      RECT 13.3 5.915 13.59 6.145 ;
      RECT 13.3 5.945 13.76 6.115 ;
      RECT 12.305 1.965 12.655 2.315 ;
      RECT 12.135 2.025 12.655 2.195 ;
      RECT 12.33 6.655 12.655 6.98 ;
      RECT 12.305 6.655 12.655 6.885 ;
      RECT 12.135 6.685 12.655 6.855 ;
      RECT 9.925 2.705 10.265 3.055 ;
      RECT 10.015 2.395 10.185 3.055 ;
      RECT 11.53 2.365 11.85 2.685 ;
      RECT 11.5 2.365 11.85 2.595 ;
      RECT 10.015 2.395 11.85 2.565 ;
      RECT 11.53 6.28 11.85 6.605 ;
      RECT 11.5 6.285 11.85 6.515 ;
      RECT 11.33 6.315 11.85 6.485 ;
      RECT 10.485 2.705 10.825 3.055 ;
      RECT 10.485 2.765 10.965 2.935 ;
      RECT 10.48 5.86 10.82 6.21 ;
      RECT 10.48 5.945 10.965 6.115 ;
      RECT 7.22 2.985 7.37 3.26 ;
      RECT 7.76 2.065 7.765 2.285 ;
      RECT 8.91 2.265 8.925 2.463 ;
      RECT 8.875 2.257 8.91 2.47 ;
      RECT 8.845 2.25 8.875 2.47 ;
      RECT 8.79 2.215 8.845 2.47 ;
      RECT 8.725 2.152 8.79 2.47 ;
      RECT 8.72 2.117 8.725 2.468 ;
      RECT 8.715 2.112 8.72 2.46 ;
      RECT 8.71 2.107 8.715 2.446 ;
      RECT 8.705 2.104 8.71 2.439 ;
      RECT 8.66 2.094 8.705 2.39 ;
      RECT 8.64 2.081 8.66 2.325 ;
      RECT 8.635 2.076 8.64 2.298 ;
      RECT 8.63 2.075 8.635 2.291 ;
      RECT 8.625 2.074 8.63 2.284 ;
      RECT 8.54 2.059 8.625 2.23 ;
      RECT 8.51 2.04 8.54 2.18 ;
      RECT 8.43 2.023 8.51 2.165 ;
      RECT 8.395 2.01 8.43 2.15 ;
      RECT 8.387 2.01 8.395 2.145 ;
      RECT 8.301 2.011 8.387 2.145 ;
      RECT 8.215 2.013 8.301 2.145 ;
      RECT 8.19 2.014 8.215 2.149 ;
      RECT 8.115 2.02 8.19 2.164 ;
      RECT 8.032 2.032 8.115 2.188 ;
      RECT 7.946 2.045 8.032 2.214 ;
      RECT 7.86 2.058 7.946 2.24 ;
      RECT 7.825 2.067 7.86 2.259 ;
      RECT 7.775 2.067 7.825 2.272 ;
      RECT 7.765 2.065 7.775 2.283 ;
      RECT 7.75 2.062 7.76 2.285 ;
      RECT 7.735 2.054 7.75 2.293 ;
      RECT 7.72 2.046 7.735 2.313 ;
      RECT 7.715 2.041 7.72 2.37 ;
      RECT 7.7 2.036 7.715 2.443 ;
      RECT 7.695 2.031 7.7 2.485 ;
      RECT 7.69 2.029 7.695 2.513 ;
      RECT 7.685 2.027 7.69 2.535 ;
      RECT 7.675 2.023 7.685 2.578 ;
      RECT 7.67 2.02 7.675 2.603 ;
      RECT 7.665 2.018 7.67 2.623 ;
      RECT 7.66 2.016 7.665 2.647 ;
      RECT 7.655 2.012 7.66 2.67 ;
      RECT 7.65 2.008 7.655 2.693 ;
      RECT 7.615 1.998 7.65 2.8 ;
      RECT 7.61 1.988 7.615 2.898 ;
      RECT 7.605 1.986 7.61 2.925 ;
      RECT 7.6 1.985 7.605 2.945 ;
      RECT 7.595 1.977 7.6 2.965 ;
      RECT 7.59 1.972 7.595 3 ;
      RECT 7.585 1.97 7.59 3.018 ;
      RECT 7.58 1.97 7.585 3.043 ;
      RECT 7.575 1.97 7.58 3.065 ;
      RECT 7.54 1.97 7.575 3.108 ;
      RECT 7.515 1.97 7.54 3.137 ;
      RECT 7.505 1.97 7.515 2.323 ;
      RECT 7.508 2.38 7.515 3.147 ;
      RECT 7.505 2.437 7.508 3.15 ;
      RECT 7.5 1.97 7.505 2.295 ;
      RECT 7.5 2.487 7.505 3.153 ;
      RECT 7.49 1.97 7.5 2.285 ;
      RECT 7.495 2.54 7.5 3.156 ;
      RECT 7.49 2.625 7.495 3.16 ;
      RECT 7.48 1.97 7.49 2.273 ;
      RECT 7.485 2.672 7.49 3.164 ;
      RECT 7.48 2.747 7.485 3.168 ;
      RECT 7.445 1.97 7.48 2.248 ;
      RECT 7.47 2.83 7.48 3.173 ;
      RECT 7.46 2.897 7.47 3.18 ;
      RECT 7.455 2.925 7.46 3.185 ;
      RECT 7.445 2.938 7.455 3.191 ;
      RECT 7.4 1.97 7.445 2.205 ;
      RECT 7.44 2.943 7.445 3.198 ;
      RECT 7.4 2.96 7.44 3.26 ;
      RECT 7.395 1.972 7.4 2.178 ;
      RECT 7.37 2.98 7.4 3.26 ;
      RECT 7.39 1.977 7.395 2.15 ;
      RECT 7.18 2.989 7.22 3.26 ;
      RECT 7.155 2.997 7.18 3.23 ;
      RECT 7.11 3.005 7.155 3.23 ;
      RECT 7.095 3.01 7.11 3.225 ;
      RECT 7.085 3.01 7.095 3.219 ;
      RECT 7.075 3.017 7.085 3.216 ;
      RECT 7.07 3.055 7.075 3.205 ;
      RECT 7.065 3.117 7.07 3.183 ;
      RECT 8.335 2.992 8.52 3.215 ;
      RECT 8.335 3.007 8.525 3.211 ;
      RECT 8.325 2.28 8.41 3.21 ;
      RECT 8.325 3.007 8.53 3.204 ;
      RECT 8.32 3.015 8.53 3.203 ;
      RECT 8.525 2.735 8.845 3.055 ;
      RECT 8.32 2.907 8.49 2.998 ;
      RECT 8.315 2.907 8.49 2.98 ;
      RECT 8.305 2.715 8.44 2.955 ;
      RECT 8.3 2.715 8.44 2.9 ;
      RECT 8.26 2.295 8.43 2.8 ;
      RECT 8.245 2.295 8.43 2.67 ;
      RECT 8.24 2.295 8.43 2.623 ;
      RECT 8.235 2.295 8.43 2.603 ;
      RECT 8.23 2.295 8.43 2.578 ;
      RECT 8.2 2.295 8.46 2.555 ;
      RECT 8.21 2.292 8.42 2.555 ;
      RECT 8.335 2.287 8.42 3.215 ;
      RECT 8.22 2.28 8.41 2.555 ;
      RECT 8.215 2.285 8.41 2.555 ;
      RECT 7.045 2.497 7.23 2.71 ;
      RECT 7.045 2.505 7.24 2.703 ;
      RECT 7.025 2.505 7.24 2.7 ;
      RECT 7.02 2.505 7.24 2.685 ;
      RECT 6.95 2.42 7.21 2.68 ;
      RECT 6.95 2.565 7.245 2.593 ;
      RECT 6.605 3.02 6.865 3.28 ;
      RECT 6.63 2.965 6.825 3.28 ;
      RECT 6.625 2.714 6.805 3.008 ;
      RECT 6.625 2.72 6.815 3.008 ;
      RECT 6.605 2.722 6.815 2.953 ;
      RECT 6.6 2.732 6.815 2.82 ;
      RECT 6.63 2.712 6.805 3.28 ;
      RECT 6.716 2.71 6.805 3.28 ;
      RECT 6.575 1.93 6.61 2.3 ;
      RECT 6.365 2.04 6.37 2.3 ;
      RECT 6.61 1.937 6.625 2.3 ;
      RECT 6.5 1.93 6.575 2.378 ;
      RECT 6.49 1.93 6.5 2.463 ;
      RECT 6.465 1.93 6.49 2.498 ;
      RECT 6.425 1.93 6.465 2.566 ;
      RECT 6.415 1.937 6.425 2.618 ;
      RECT 6.385 2.04 6.415 2.659 ;
      RECT 6.38 2.04 6.385 2.698 ;
      RECT 6.37 2.04 6.38 2.718 ;
      RECT 6.365 2.335 6.37 2.755 ;
      RECT 6.36 2.352 6.365 2.775 ;
      RECT 6.345 2.415 6.36 2.815 ;
      RECT 6.34 2.458 6.345 2.85 ;
      RECT 6.335 2.466 6.34 2.863 ;
      RECT 6.325 2.48 6.335 2.885 ;
      RECT 6.3 2.515 6.325 2.95 ;
      RECT 6.29 2.55 6.3 3.013 ;
      RECT 6.27 2.58 6.29 3.074 ;
      RECT 6.255 2.616 6.27 3.141 ;
      RECT 6.245 2.644 6.255 3.18 ;
      RECT 6.235 2.666 6.245 3.2 ;
      RECT 6.23 2.676 6.235 3.211 ;
      RECT 6.225 2.685 6.23 3.214 ;
      RECT 6.215 2.703 6.225 3.218 ;
      RECT 6.205 2.721 6.215 3.219 ;
      RECT 6.18 2.76 6.205 3.216 ;
      RECT 6.16 2.802 6.18 3.213 ;
      RECT 6.145 2.84 6.16 3.212 ;
      RECT 6.11 2.875 6.145 3.209 ;
      RECT 6.105 2.897 6.11 3.207 ;
      RECT 6.04 2.937 6.105 3.204 ;
      RECT 6.035 2.977 6.04 3.2 ;
      RECT 6.02 2.987 6.035 3.191 ;
      RECT 6.01 3.107 6.02 3.176 ;
      RECT 6.49 3.52 6.5 3.78 ;
      RECT 6.49 3.523 6.51 3.779 ;
      RECT 6.48 3.513 6.49 3.778 ;
      RECT 6.47 3.528 6.55 3.774 ;
      RECT 6.455 3.507 6.47 3.772 ;
      RECT 6.43 3.532 6.555 3.768 ;
      RECT 6.415 3.492 6.43 3.763 ;
      RECT 6.415 3.534 6.565 3.762 ;
      RECT 6.415 3.542 6.58 3.755 ;
      RECT 6.355 3.479 6.415 3.745 ;
      RECT 6.345 3.466 6.355 3.727 ;
      RECT 6.32 3.456 6.345 3.717 ;
      RECT 6.315 3.446 6.32 3.709 ;
      RECT 6.25 3.542 6.58 3.691 ;
      RECT 6.165 3.542 6.58 3.653 ;
      RECT 6.055 3.37 6.315 3.63 ;
      RECT 6.43 3.5 6.455 3.768 ;
      RECT 6.47 3.51 6.48 3.774 ;
      RECT 6.055 3.518 6.495 3.63 ;
      RECT 5.27 3.275 5.3 3.575 ;
      RECT 5.045 3.26 5.05 3.535 ;
      RECT 4.845 3.26 5 3.52 ;
      RECT 6.145 1.975 6.175 2.235 ;
      RECT 6.135 1.975 6.145 2.343 ;
      RECT 6.115 1.975 6.135 2.353 ;
      RECT 6.1 1.975 6.115 2.365 ;
      RECT 6.045 1.975 6.1 2.415 ;
      RECT 6.03 1.975 6.045 2.463 ;
      RECT 6 1.975 6.03 2.498 ;
      RECT 5.945 1.975 6 2.56 ;
      RECT 5.925 1.975 5.945 2.628 ;
      RECT 5.92 1.975 5.925 2.658 ;
      RECT 5.915 1.975 5.92 2.67 ;
      RECT 5.91 2.092 5.915 2.688 ;
      RECT 5.89 2.11 5.91 2.713 ;
      RECT 5.87 2.137 5.89 2.763 ;
      RECT 5.865 2.157 5.87 2.794 ;
      RECT 5.86 2.165 5.865 2.811 ;
      RECT 5.845 2.191 5.86 2.84 ;
      RECT 5.83 2.233 5.845 2.875 ;
      RECT 5.825 2.262 5.83 2.898 ;
      RECT 5.82 2.277 5.825 2.911 ;
      RECT 5.815 2.3 5.82 2.922 ;
      RECT 5.805 2.32 5.815 2.94 ;
      RECT 5.795 2.35 5.805 2.963 ;
      RECT 5.79 2.372 5.795 2.983 ;
      RECT 5.785 2.387 5.79 2.998 ;
      RECT 5.77 2.417 5.785 3.025 ;
      RECT 5.765 2.447 5.77 3.051 ;
      RECT 5.76 2.465 5.765 3.063 ;
      RECT 5.75 2.495 5.76 3.082 ;
      RECT 5.74 2.52 5.75 3.107 ;
      RECT 5.735 2.54 5.74 3.126 ;
      RECT 5.73 2.557 5.735 3.139 ;
      RECT 5.72 2.583 5.73 3.158 ;
      RECT 5.71 2.621 5.72 3.185 ;
      RECT 5.705 2.647 5.71 3.205 ;
      RECT 5.7 2.657 5.705 3.215 ;
      RECT 5.695 2.67 5.7 3.23 ;
      RECT 5.69 2.685 5.695 3.24 ;
      RECT 5.685 2.707 5.69 3.255 ;
      RECT 5.68 2.725 5.685 3.266 ;
      RECT 5.675 2.735 5.68 3.277 ;
      RECT 5.67 2.743 5.675 3.289 ;
      RECT 5.665 2.751 5.67 3.3 ;
      RECT 5.66 2.777 5.665 3.313 ;
      RECT 5.65 2.805 5.66 3.326 ;
      RECT 5.645 2.835 5.65 3.335 ;
      RECT 5.64 2.85 5.645 3.342 ;
      RECT 5.625 2.875 5.64 3.349 ;
      RECT 5.62 2.897 5.625 3.355 ;
      RECT 5.615 2.922 5.62 3.358 ;
      RECT 5.606 2.95 5.615 3.362 ;
      RECT 5.6 2.967 5.606 3.367 ;
      RECT 5.595 2.985 5.6 3.371 ;
      RECT 5.59 2.997 5.595 3.374 ;
      RECT 5.585 3.018 5.59 3.378 ;
      RECT 5.58 3.036 5.585 3.381 ;
      RECT 5.575 3.05 5.58 3.384 ;
      RECT 5.57 3.067 5.575 3.387 ;
      RECT 5.565 3.08 5.57 3.39 ;
      RECT 5.54 3.117 5.565 3.398 ;
      RECT 5.535 3.162 5.54 3.407 ;
      RECT 5.53 3.19 5.535 3.41 ;
      RECT 5.52 3.21 5.53 3.414 ;
      RECT 5.515 3.23 5.52 3.419 ;
      RECT 5.51 3.245 5.515 3.422 ;
      RECT 5.49 3.255 5.51 3.429 ;
      RECT 5.425 3.262 5.49 3.455 ;
      RECT 5.39 3.265 5.425 3.483 ;
      RECT 5.375 3.268 5.39 3.498 ;
      RECT 5.365 3.269 5.375 3.513 ;
      RECT 5.355 3.27 5.365 3.53 ;
      RECT 5.35 3.27 5.355 3.545 ;
      RECT 5.345 3.27 5.35 3.553 ;
      RECT 5.33 3.271 5.345 3.568 ;
      RECT 5.3 3.273 5.33 3.575 ;
      RECT 5.19 3.28 5.27 3.575 ;
      RECT 5.145 3.285 5.19 3.575 ;
      RECT 5.135 3.286 5.145 3.565 ;
      RECT 5.125 3.287 5.135 3.558 ;
      RECT 5.105 3.289 5.125 3.553 ;
      RECT 5.095 3.26 5.105 3.548 ;
      RECT 5.05 3.26 5.095 3.54 ;
      RECT 5.02 3.26 5.045 3.53 ;
      RECT 5 3.26 5.02 3.523 ;
      RECT 5.28 2.06 5.54 2.32 ;
      RECT 5.16 2.075 5.17 2.24 ;
      RECT 5.145 2.075 5.15 2.235 ;
      RECT 2.51 1.915 2.695 2.205 ;
      RECT 4.325 2.04 4.34 2.195 ;
      RECT 2.475 1.915 2.5 2.175 ;
      RECT 4.89 1.965 4.895 2.107 ;
      RECT 4.805 1.96 4.83 2.1 ;
      RECT 5.205 2.077 5.28 2.27 ;
      RECT 5.19 2.075 5.205 2.253 ;
      RECT 5.17 2.075 5.19 2.245 ;
      RECT 5.15 2.075 5.16 2.238 ;
      RECT 5.105 2.07 5.145 2.228 ;
      RECT 5.065 2.045 5.105 2.213 ;
      RECT 5.05 2.02 5.065 2.203 ;
      RECT 5.045 2.014 5.05 2.201 ;
      RECT 5.01 2.006 5.045 2.184 ;
      RECT 5.005 1.999 5.01 2.172 ;
      RECT 4.985 1.994 5.005 2.16 ;
      RECT 4.975 1.988 4.985 2.145 ;
      RECT 4.955 1.983 4.975 2.13 ;
      RECT 4.945 1.978 4.955 2.123 ;
      RECT 4.94 1.976 4.945 2.118 ;
      RECT 4.935 1.975 4.94 2.115 ;
      RECT 4.895 1.97 4.935 2.111 ;
      RECT 4.875 1.964 4.89 2.106 ;
      RECT 4.84 1.961 4.875 2.103 ;
      RECT 4.83 1.96 4.84 2.101 ;
      RECT 4.77 1.96 4.805 2.098 ;
      RECT 4.725 1.96 4.77 2.098 ;
      RECT 4.675 1.96 4.725 2.101 ;
      RECT 4.66 1.962 4.675 2.103 ;
      RECT 4.645 1.965 4.66 2.104 ;
      RECT 4.635 1.97 4.645 2.105 ;
      RECT 4.605 1.975 4.635 2.11 ;
      RECT 4.595 1.981 4.605 2.118 ;
      RECT 4.585 1.983 4.595 2.122 ;
      RECT 4.575 1.987 4.585 2.126 ;
      RECT 4.55 1.993 4.575 2.134 ;
      RECT 4.54 1.998 4.55 2.142 ;
      RECT 4.525 2.002 4.54 2.146 ;
      RECT 4.49 2.008 4.525 2.154 ;
      RECT 4.47 2.013 4.49 2.164 ;
      RECT 4.44 2.02 4.47 2.173 ;
      RECT 4.395 2.029 4.44 2.187 ;
      RECT 4.39 2.034 4.395 2.198 ;
      RECT 4.37 2.037 4.39 2.199 ;
      RECT 4.34 2.04 4.37 2.197 ;
      RECT 4.305 2.04 4.325 2.193 ;
      RECT 4.235 2.04 4.305 2.184 ;
      RECT 4.22 2.037 4.235 2.176 ;
      RECT 4.18 2.03 4.22 2.171 ;
      RECT 4.155 2.02 4.18 2.164 ;
      RECT 4.15 2.014 4.155 2.161 ;
      RECT 4.11 2.008 4.15 2.158 ;
      RECT 4.095 2.001 4.11 2.153 ;
      RECT 4.075 1.997 4.095 2.148 ;
      RECT 4.06 1.992 4.075 2.144 ;
      RECT 4.045 1.987 4.06 2.142 ;
      RECT 4.03 1.983 4.045 2.141 ;
      RECT 4.015 1.981 4.03 2.137 ;
      RECT 4.005 1.979 4.015 2.132 ;
      RECT 3.99 1.976 4.005 2.128 ;
      RECT 3.98 1.974 3.99 2.123 ;
      RECT 3.96 1.971 3.98 2.119 ;
      RECT 3.915 1.97 3.96 2.117 ;
      RECT 3.855 1.972 3.915 2.118 ;
      RECT 3.835 1.974 3.855 2.12 ;
      RECT 3.805 1.977 3.835 2.121 ;
      RECT 3.755 1.982 3.805 2.123 ;
      RECT 3.75 1.985 3.755 2.125 ;
      RECT 3.74 1.987 3.75 2.128 ;
      RECT 3.735 1.989 3.74 2.131 ;
      RECT 3.685 1.992 3.735 2.138 ;
      RECT 3.665 1.996 3.685 2.15 ;
      RECT 3.655 1.999 3.665 2.156 ;
      RECT 3.645 2 3.655 2.159 ;
      RECT 3.606 2.003 3.645 2.161 ;
      RECT 3.52 2.01 3.606 2.164 ;
      RECT 3.446 2.02 3.52 2.168 ;
      RECT 3.36 2.031 3.446 2.173 ;
      RECT 3.345 2.038 3.36 2.175 ;
      RECT 3.29 2.042 3.345 2.176 ;
      RECT 3.276 2.045 3.29 2.178 ;
      RECT 3.19 2.045 3.276 2.18 ;
      RECT 3.15 2.042 3.19 2.183 ;
      RECT 3.126 2.038 3.15 2.185 ;
      RECT 3.04 2.028 3.126 2.188 ;
      RECT 3.01 2.017 3.04 2.189 ;
      RECT 2.991 2.013 3.01 2.188 ;
      RECT 2.905 2.006 2.991 2.185 ;
      RECT 2.845 1.995 2.905 2.182 ;
      RECT 2.825 1.987 2.845 2.18 ;
      RECT 2.79 1.982 2.825 2.179 ;
      RECT 2.765 1.977 2.79 2.178 ;
      RECT 2.735 1.972 2.765 2.177 ;
      RECT 2.71 1.915 2.735 2.176 ;
      RECT 2.695 1.915 2.71 2.2 ;
      RECT 2.5 1.915 2.51 2.2 ;
      RECT 4.275 2.935 4.28 3.075 ;
      RECT 3.935 2.935 3.97 3.073 ;
      RECT 3.51 2.92 3.525 3.065 ;
      RECT 5.34 2.7 5.43 2.96 ;
      RECT 5.17 2.565 5.27 2.96 ;
      RECT 2.205 2.54 2.285 2.75 ;
      RECT 5.295 2.677 5.34 2.96 ;
      RECT 5.285 2.647 5.295 2.96 ;
      RECT 5.27 2.57 5.285 2.96 ;
      RECT 5.085 2.565 5.17 2.925 ;
      RECT 5.08 2.567 5.085 2.92 ;
      RECT 5.075 2.572 5.08 2.92 ;
      RECT 5.04 2.672 5.075 2.92 ;
      RECT 5.03 2.7 5.04 2.92 ;
      RECT 5.02 2.715 5.03 2.92 ;
      RECT 5.01 2.727 5.02 2.92 ;
      RECT 5.005 2.737 5.01 2.92 ;
      RECT 4.99 2.747 5.005 2.922 ;
      RECT 4.985 2.762 4.99 2.924 ;
      RECT 4.97 2.775 4.985 2.926 ;
      RECT 4.965 2.79 4.97 2.929 ;
      RECT 4.945 2.8 4.965 2.933 ;
      RECT 4.93 2.81 4.945 2.936 ;
      RECT 4.895 2.817 4.93 2.941 ;
      RECT 4.851 2.824 4.895 2.949 ;
      RECT 4.765 2.836 4.851 2.962 ;
      RECT 4.74 2.847 4.765 2.973 ;
      RECT 4.71 2.852 4.74 2.978 ;
      RECT 4.675 2.857 4.71 2.986 ;
      RECT 4.645 2.862 4.675 2.993 ;
      RECT 4.62 2.867 4.645 2.998 ;
      RECT 4.555 2.874 4.62 3.007 ;
      RECT 4.485 2.887 4.555 3.023 ;
      RECT 4.455 2.897 4.485 3.035 ;
      RECT 4.43 2.902 4.455 3.042 ;
      RECT 4.375 2.909 4.43 3.05 ;
      RECT 4.37 2.916 4.375 3.055 ;
      RECT 4.365 2.918 4.37 3.056 ;
      RECT 4.35 2.92 4.365 3.058 ;
      RECT 4.345 2.92 4.35 3.061 ;
      RECT 4.28 2.927 4.345 3.068 ;
      RECT 4.245 2.937 4.275 3.078 ;
      RECT 4.228 2.94 4.245 3.08 ;
      RECT 4.142 2.939 4.228 3.079 ;
      RECT 4.056 2.937 4.142 3.076 ;
      RECT 3.97 2.936 4.056 3.074 ;
      RECT 3.869 2.934 3.935 3.073 ;
      RECT 3.783 2.931 3.869 3.071 ;
      RECT 3.697 2.927 3.783 3.069 ;
      RECT 3.611 2.924 3.697 3.068 ;
      RECT 3.525 2.921 3.611 3.066 ;
      RECT 3.425 2.92 3.51 3.063 ;
      RECT 3.375 2.918 3.425 3.061 ;
      RECT 3.355 2.915 3.375 3.059 ;
      RECT 3.335 2.913 3.355 3.056 ;
      RECT 3.31 2.909 3.335 3.053 ;
      RECT 3.265 2.903 3.31 3.048 ;
      RECT 3.225 2.897 3.265 3.04 ;
      RECT 3.2 2.892 3.225 3.033 ;
      RECT 3.145 2.885 3.2 3.025 ;
      RECT 3.121 2.878 3.145 3.018 ;
      RECT 3.035 2.869 3.121 3.008 ;
      RECT 3.005 2.861 3.035 2.998 ;
      RECT 2.975 2.857 3.005 2.993 ;
      RECT 2.97 2.854 2.975 2.99 ;
      RECT 2.965 2.853 2.97 2.99 ;
      RECT 2.89 2.846 2.965 2.983 ;
      RECT 2.851 2.837 2.89 2.972 ;
      RECT 2.765 2.827 2.851 2.96 ;
      RECT 2.725 2.817 2.765 2.948 ;
      RECT 2.686 2.812 2.725 2.941 ;
      RECT 2.6 2.802 2.686 2.93 ;
      RECT 2.56 2.79 2.6 2.919 ;
      RECT 2.525 2.775 2.56 2.912 ;
      RECT 2.515 2.765 2.525 2.909 ;
      RECT 2.495 2.75 2.515 2.907 ;
      RECT 2.465 2.72 2.495 2.903 ;
      RECT 2.455 2.7 2.465 2.898 ;
      RECT 2.45 2.692 2.455 2.895 ;
      RECT 2.445 2.685 2.45 2.893 ;
      RECT 2.43 2.672 2.445 2.886 ;
      RECT 2.425 2.662 2.43 2.878 ;
      RECT 2.42 2.655 2.425 2.873 ;
      RECT 2.415 2.65 2.42 2.869 ;
      RECT 2.4 2.637 2.415 2.861 ;
      RECT 2.395 2.547 2.4 2.85 ;
      RECT 2.39 2.542 2.395 2.843 ;
      RECT 2.315 2.54 2.39 2.803 ;
      RECT 2.285 2.54 2.315 2.758 ;
      RECT 2.19 2.545 2.205 2.745 ;
      RECT 4.675 2.25 4.935 2.51 ;
      RECT 4.66 2.238 4.84 2.475 ;
      RECT 4.655 2.239 4.84 2.473 ;
      RECT 4.64 2.243 4.85 2.463 ;
      RECT 4.635 2.248 4.855 2.433 ;
      RECT 4.64 2.245 4.855 2.463 ;
      RECT 4.655 2.24 4.85 2.473 ;
      RECT 4.675 2.237 4.84 2.51 ;
      RECT 4.675 2.236 4.83 2.51 ;
      RECT 4.7 2.235 4.83 2.51 ;
      RECT 4.26 2.48 4.52 2.74 ;
      RECT 4.135 2.525 4.52 2.735 ;
      RECT 4.125 2.53 4.52 2.73 ;
      RECT 4.14 3.47 4.155 3.78 ;
      RECT 2.735 3.24 2.745 3.37 ;
      RECT 2.515 3.235 2.62 3.37 ;
      RECT 2.43 3.24 2.48 3.37 ;
      RECT 0.98 1.975 0.985 3.08 ;
      RECT 4.235 3.562 4.24 3.698 ;
      RECT 4.23 3.557 4.235 3.758 ;
      RECT 4.225 3.555 4.23 3.771 ;
      RECT 4.21 3.552 4.225 3.773 ;
      RECT 4.205 3.547 4.21 3.775 ;
      RECT 4.2 3.543 4.205 3.778 ;
      RECT 4.185 3.538 4.2 3.78 ;
      RECT 4.155 3.53 4.185 3.78 ;
      RECT 4.116 3.47 4.14 3.78 ;
      RECT 4.03 3.47 4.116 3.777 ;
      RECT 4 3.47 4.03 3.77 ;
      RECT 3.975 3.47 4 3.763 ;
      RECT 3.95 3.47 3.975 3.755 ;
      RECT 3.935 3.47 3.95 3.748 ;
      RECT 3.91 3.47 3.935 3.74 ;
      RECT 3.895 3.47 3.91 3.733 ;
      RECT 3.855 3.48 3.895 3.722 ;
      RECT 3.845 3.475 3.855 3.712 ;
      RECT 3.841 3.474 3.845 3.709 ;
      RECT 3.755 3.466 3.841 3.692 ;
      RECT 3.722 3.455 3.755 3.669 ;
      RECT 3.636 3.444 3.722 3.647 ;
      RECT 3.55 3.428 3.636 3.616 ;
      RECT 3.48 3.413 3.55 3.588 ;
      RECT 3.47 3.406 3.48 3.575 ;
      RECT 3.44 3.403 3.47 3.565 ;
      RECT 3.415 3.399 3.44 3.558 ;
      RECT 3.4 3.396 3.415 3.553 ;
      RECT 3.395 3.395 3.4 3.548 ;
      RECT 3.365 3.39 3.395 3.541 ;
      RECT 3.36 3.385 3.365 3.536 ;
      RECT 3.345 3.382 3.36 3.531 ;
      RECT 3.34 3.377 3.345 3.526 ;
      RECT 3.32 3.372 3.34 3.523 ;
      RECT 3.305 3.367 3.32 3.515 ;
      RECT 3.29 3.361 3.305 3.51 ;
      RECT 3.26 3.352 3.29 3.503 ;
      RECT 3.255 3.345 3.26 3.495 ;
      RECT 3.25 3.343 3.255 3.493 ;
      RECT 3.245 3.342 3.25 3.49 ;
      RECT 3.205 3.335 3.245 3.483 ;
      RECT 3.191 3.325 3.205 3.473 ;
      RECT 3.14 3.314 3.191 3.461 ;
      RECT 3.115 3.3 3.14 3.447 ;
      RECT 3.09 3.289 3.115 3.439 ;
      RECT 3.07 3.278 3.09 3.433 ;
      RECT 3.06 3.272 3.07 3.428 ;
      RECT 3.055 3.27 3.06 3.424 ;
      RECT 3.035 3.265 3.055 3.419 ;
      RECT 3.005 3.255 3.035 3.409 ;
      RECT 3 3.247 3.005 3.402 ;
      RECT 2.985 3.245 3 3.398 ;
      RECT 2.965 3.245 2.985 3.393 ;
      RECT 2.96 3.244 2.965 3.391 ;
      RECT 2.955 3.244 2.96 3.388 ;
      RECT 2.915 3.243 2.955 3.383 ;
      RECT 2.89 3.242 2.915 3.378 ;
      RECT 2.83 3.241 2.89 3.375 ;
      RECT 2.745 3.24 2.83 3.373 ;
      RECT 2.706 3.239 2.735 3.37 ;
      RECT 2.62 3.237 2.706 3.37 ;
      RECT 2.48 3.237 2.515 3.37 ;
      RECT 2.39 3.241 2.43 3.373 ;
      RECT 2.375 3.244 2.39 3.38 ;
      RECT 2.365 3.245 2.375 3.387 ;
      RECT 2.34 3.248 2.365 3.392 ;
      RECT 2.335 3.25 2.34 3.395 ;
      RECT 2.285 3.252 2.335 3.396 ;
      RECT 2.246 3.256 2.285 3.398 ;
      RECT 2.16 3.258 2.246 3.401 ;
      RECT 2.142 3.26 2.16 3.403 ;
      RECT 2.056 3.263 2.142 3.405 ;
      RECT 1.97 3.267 2.056 3.408 ;
      RECT 1.933 3.271 1.97 3.411 ;
      RECT 1.847 3.274 1.933 3.414 ;
      RECT 1.761 3.278 1.847 3.417 ;
      RECT 1.675 3.283 1.761 3.421 ;
      RECT 1.655 3.285 1.675 3.424 ;
      RECT 1.635 3.284 1.655 3.425 ;
      RECT 1.586 3.281 1.635 3.426 ;
      RECT 1.5 3.276 1.586 3.429 ;
      RECT 1.45 3.271 1.5 3.431 ;
      RECT 1.426 3.269 1.45 3.432 ;
      RECT 1.34 3.264 1.426 3.434 ;
      RECT 1.315 3.26 1.34 3.433 ;
      RECT 1.305 3.257 1.315 3.431 ;
      RECT 1.295 3.25 1.305 3.428 ;
      RECT 1.29 3.23 1.295 3.423 ;
      RECT 1.28 3.2 1.29 3.418 ;
      RECT 1.265 3.07 1.28 3.409 ;
      RECT 1.26 3.062 1.265 3.402 ;
      RECT 1.24 3.055 1.26 3.394 ;
      RECT 1.235 3.037 1.24 3.386 ;
      RECT 1.225 3.017 1.235 3.381 ;
      RECT 1.22 2.99 1.225 3.377 ;
      RECT 1.215 2.967 1.22 3.374 ;
      RECT 1.195 2.925 1.215 3.366 ;
      RECT 1.16 2.84 1.195 3.35 ;
      RECT 1.155 2.772 1.16 3.338 ;
      RECT 1.14 2.742 1.155 3.332 ;
      RECT 1.135 1.987 1.14 2.233 ;
      RECT 1.125 2.712 1.14 3.323 ;
      RECT 1.13 1.982 1.135 2.265 ;
      RECT 1.125 1.977 1.13 2.308 ;
      RECT 1.12 1.975 1.125 2.343 ;
      RECT 1.105 2.675 1.125 3.313 ;
      RECT 1.115 1.975 1.12 2.38 ;
      RECT 1.1 1.975 1.115 2.478 ;
      RECT 1.1 2.648 1.105 3.306 ;
      RECT 1.095 1.975 1.1 2.553 ;
      RECT 1.095 2.636 1.1 3.303 ;
      RECT 1.09 1.975 1.095 2.585 ;
      RECT 1.09 2.615 1.095 3.3 ;
      RECT 1.085 1.975 1.09 3.297 ;
      RECT 1.05 1.975 1.085 3.283 ;
      RECT 1.035 1.975 1.05 3.265 ;
      RECT 1.015 1.975 1.035 3.255 ;
      RECT 0.99 1.975 1.015 3.238 ;
      RECT 0.985 1.975 0.99 3.188 ;
      RECT 0.975 1.975 0.98 3.018 ;
      RECT 0.97 1.975 0.975 2.925 ;
      RECT 0.965 1.975 0.97 2.838 ;
      RECT 0.96 1.975 0.965 2.77 ;
      RECT 0.955 1.975 0.96 2.713 ;
      RECT 0.945 1.975 0.955 2.608 ;
      RECT 0.94 1.975 0.945 2.48 ;
      RECT 0.935 1.975 0.94 2.398 ;
      RECT 0.93 1.977 0.935 2.315 ;
      RECT 0.925 1.982 0.93 2.248 ;
      RECT 0.92 1.987 0.925 2.175 ;
      RECT 3.735 2.305 3.995 2.565 ;
      RECT 3.755 2.272 3.965 2.565 ;
      RECT 3.755 2.27 3.955 2.565 ;
      RECT 3.765 2.257 3.955 2.565 ;
      RECT 3.765 2.255 3.88 2.565 ;
      RECT 3.24 2.38 3.415 2.66 ;
      RECT 3.235 2.38 3.415 2.658 ;
      RECT 3.235 2.38 3.43 2.655 ;
      RECT 3.225 2.38 3.43 2.653 ;
      RECT 3.17 2.38 3.43 2.64 ;
      RECT 3.17 2.455 3.435 2.618 ;
      RECT 2.715 2.392 2.735 2.635 ;
      RECT 2.715 2.392 2.775 2.634 ;
      RECT 2.71 2.394 2.775 2.633 ;
      RECT 2.71 2.394 2.861 2.632 ;
      RECT 2.71 2.394 2.93 2.631 ;
      RECT 2.71 2.394 2.95 2.623 ;
      RECT 2.69 2.397 2.95 2.621 ;
      RECT 2.675 2.407 2.95 2.606 ;
      RECT 2.675 2.407 2.965 2.605 ;
      RECT 2.67 2.416 2.965 2.597 ;
      RECT 2.67 2.416 2.97 2.593 ;
      RECT 2.775 2.33 3.035 2.59 ;
      RECT 2.665 2.418 3.035 2.475 ;
      RECT 2.735 2.385 3.035 2.59 ;
      RECT 2.7 3.578 2.705 3.785 ;
      RECT 2.65 3.572 2.7 3.784 ;
      RECT 2.617 3.586 2.71 3.783 ;
      RECT 2.531 3.586 2.71 3.782 ;
      RECT 2.445 3.586 2.71 3.781 ;
      RECT 2.445 3.685 2.715 3.778 ;
      RECT 2.44 3.685 2.715 3.773 ;
      RECT 2.435 3.685 2.715 3.755 ;
      RECT 2.43 3.685 2.715 3.738 ;
      RECT 2.39 3.47 2.65 3.73 ;
      RECT 1.85 2.62 1.936 3.034 ;
      RECT 1.85 2.62 1.975 3.031 ;
      RECT 1.85 2.62 1.995 3.021 ;
      RECT 1.805 2.62 1.995 3.018 ;
      RECT 1.805 2.772 2.005 3.008 ;
      RECT 1.805 2.793 2.01 3.002 ;
      RECT 1.805 2.811 2.015 2.998 ;
      RECT 1.805 2.831 2.025 2.993 ;
      RECT 1.78 2.831 2.025 2.99 ;
      RECT 1.77 2.831 2.025 2.968 ;
      RECT 1.77 2.847 2.03 2.938 ;
      RECT 1.735 2.62 1.995 2.925 ;
      RECT 1.735 2.859 2.035 2.88 ;
      RECT 0 8.575 76.3 8.88 ;
      RECT 65.36 3.265 65.62 3.525 ;
      RECT 50.1 3.265 50.36 3.525 ;
      RECT 34.84 3.265 35.1 3.525 ;
      RECT 19.58 3.265 19.84 3.525 ;
      RECT 4.32 3.265 4.58 3.525 ;
    LAYER mcon ;
      RECT 75.76 0.915 75.93 1.085 ;
      RECT 75.76 2.395 75.93 2.565 ;
      RECT 75.76 6.315 75.93 6.485 ;
      RECT 75.76 7.795 75.93 7.965 ;
      RECT 75.41 0.105 75.58 0.275 ;
      RECT 75.41 4.165 75.58 4.335 ;
      RECT 75.41 4.545 75.58 4.715 ;
      RECT 75.41 8.605 75.58 8.775 ;
      RECT 75.39 2.765 75.56 2.935 ;
      RECT 75.39 5.945 75.56 6.115 ;
      RECT 74.77 0.915 74.94 1.085 ;
      RECT 74.77 2.395 74.94 2.565 ;
      RECT 74.77 6.315 74.94 6.485 ;
      RECT 74.77 7.795 74.94 7.965 ;
      RECT 74.42 0.105 74.59 0.275 ;
      RECT 74.42 4.165 74.59 4.335 ;
      RECT 74.42 4.545 74.59 4.715 ;
      RECT 74.42 8.605 74.59 8.775 ;
      RECT 74.4 2.765 74.57 2.935 ;
      RECT 74.4 5.945 74.57 6.115 ;
      RECT 73.715 0.105 73.885 0.275 ;
      RECT 73.715 4.165 73.885 4.335 ;
      RECT 73.715 4.545 73.885 4.715 ;
      RECT 73.715 8.605 73.885 8.775 ;
      RECT 73.405 2.025 73.575 2.195 ;
      RECT 73.405 6.685 73.575 6.855 ;
      RECT 73.035 0.105 73.205 0.275 ;
      RECT 73.035 8.605 73.205 8.775 ;
      RECT 72.975 0.915 73.145 1.085 ;
      RECT 72.975 1.655 73.145 1.825 ;
      RECT 72.975 7.055 73.145 7.225 ;
      RECT 72.975 7.795 73.145 7.965 ;
      RECT 72.6 2.395 72.77 2.565 ;
      RECT 72.6 6.315 72.77 6.485 ;
      RECT 72.355 0.105 72.525 0.275 ;
      RECT 72.355 8.605 72.525 8.775 ;
      RECT 71.675 0.105 71.845 0.275 ;
      RECT 71.675 8.605 71.845 8.775 ;
      RECT 71.605 2.765 71.775 2.935 ;
      RECT 71.605 5.945 71.775 6.115 ;
      RECT 70.215 1.415 70.385 1.585 ;
      RECT 70.215 4.135 70.385 4.305 ;
      RECT 69.775 2.28 69.945 2.45 ;
      RECT 69.755 1.415 69.925 1.585 ;
      RECT 69.755 4.135 69.925 4.305 ;
      RECT 69.38 3.025 69.55 3.195 ;
      RECT 69.295 1.415 69.465 1.585 ;
      RECT 69.295 4.135 69.465 4.305 ;
      RECT 69.27 2.3 69.44 2.47 ;
      RECT 68.835 1.415 69.005 1.585 ;
      RECT 68.835 4.135 69.005 4.305 ;
      RECT 68.45 1.99 68.62 2.16 ;
      RECT 68.375 1.415 68.545 1.585 ;
      RECT 68.375 4.135 68.545 4.305 ;
      RECT 68.135 3.03 68.305 3.2 ;
      RECT 68.09 2.52 68.26 2.69 ;
      RECT 67.915 1.415 68.085 1.585 ;
      RECT 67.915 4.135 68.085 4.305 ;
      RECT 67.665 2.73 67.835 2.9 ;
      RECT 67.475 1.95 67.645 2.12 ;
      RECT 67.455 1.415 67.625 1.585 ;
      RECT 67.455 4.135 67.625 4.305 ;
      RECT 67.425 3.56 67.595 3.73 ;
      RECT 67.09 3 67.26 3.17 ;
      RECT 66.995 1.415 67.165 1.585 ;
      RECT 66.995 2.16 67.165 2.33 ;
      RECT 66.995 4.135 67.165 4.305 ;
      RECT 66.535 1.415 66.705 1.585 ;
      RECT 66.535 4.135 66.705 4.305 ;
      RECT 66.195 3.385 66.365 3.555 ;
      RECT 66.135 2.585 66.305 2.755 ;
      RECT 66.075 1.415 66.245 1.585 ;
      RECT 66.075 4.135 66.245 4.305 ;
      RECT 65.695 2.255 65.865 2.425 ;
      RECT 65.615 1.415 65.785 1.585 ;
      RECT 65.615 4.135 65.785 4.305 ;
      RECT 65.43 3.305 65.6 3.475 ;
      RECT 65.185 2.545 65.355 2.715 ;
      RECT 65.155 1.415 65.325 1.585 ;
      RECT 65.155 4.135 65.325 4.305 ;
      RECT 65.09 3.575 65.26 3.745 ;
      RECT 64.815 2.27 64.985 2.44 ;
      RECT 64.695 1.415 64.865 1.585 ;
      RECT 64.695 4.135 64.865 4.305 ;
      RECT 64.285 2.47 64.455 2.64 ;
      RECT 64.235 1.415 64.405 1.585 ;
      RECT 64.235 4.135 64.405 4.305 ;
      RECT 63.775 1.415 63.945 1.585 ;
      RECT 63.775 4.135 63.945 4.305 ;
      RECT 63.765 2.415 63.935 2.585 ;
      RECT 63.56 2.015 63.73 2.185 ;
      RECT 63.56 3.595 63.73 3.765 ;
      RECT 63.315 1.415 63.485 1.585 ;
      RECT 63.315 4.135 63.485 4.305 ;
      RECT 63.25 2.56 63.42 2.73 ;
      RECT 62.855 1.415 63.025 1.585 ;
      RECT 62.855 4.135 63.025 4.305 ;
      RECT 62.84 2.785 63.01 2.955 ;
      RECT 62.395 1.415 62.565 1.585 ;
      RECT 62.395 4.135 62.565 4.305 ;
      RECT 62.13 3.085 62.3 3.255 ;
      RECT 61.985 1.995 62.155 2.165 ;
      RECT 61.935 1.415 62.105 1.585 ;
      RECT 61.935 4.135 62.105 4.305 ;
      RECT 60.5 0.915 60.67 1.085 ;
      RECT 60.5 2.395 60.67 2.565 ;
      RECT 60.5 6.315 60.67 6.485 ;
      RECT 60.5 7.795 60.67 7.965 ;
      RECT 60.15 0.105 60.32 0.275 ;
      RECT 60.15 4.165 60.32 4.335 ;
      RECT 60.15 4.545 60.32 4.715 ;
      RECT 60.15 8.605 60.32 8.775 ;
      RECT 60.13 2.765 60.3 2.935 ;
      RECT 60.13 5.945 60.3 6.115 ;
      RECT 59.51 0.915 59.68 1.085 ;
      RECT 59.51 2.395 59.68 2.565 ;
      RECT 59.51 6.315 59.68 6.485 ;
      RECT 59.51 7.795 59.68 7.965 ;
      RECT 59.16 0.105 59.33 0.275 ;
      RECT 59.16 4.165 59.33 4.335 ;
      RECT 59.16 4.545 59.33 4.715 ;
      RECT 59.16 8.605 59.33 8.775 ;
      RECT 59.14 2.765 59.31 2.935 ;
      RECT 59.14 5.945 59.31 6.115 ;
      RECT 58.455 0.105 58.625 0.275 ;
      RECT 58.455 4.165 58.625 4.335 ;
      RECT 58.455 4.545 58.625 4.715 ;
      RECT 58.455 8.605 58.625 8.775 ;
      RECT 58.145 2.025 58.315 2.195 ;
      RECT 58.145 6.685 58.315 6.855 ;
      RECT 57.775 0.105 57.945 0.275 ;
      RECT 57.775 8.605 57.945 8.775 ;
      RECT 57.715 0.915 57.885 1.085 ;
      RECT 57.715 1.655 57.885 1.825 ;
      RECT 57.715 7.055 57.885 7.225 ;
      RECT 57.715 7.795 57.885 7.965 ;
      RECT 57.34 2.395 57.51 2.565 ;
      RECT 57.34 6.315 57.51 6.485 ;
      RECT 57.095 0.105 57.265 0.275 ;
      RECT 57.095 8.605 57.265 8.775 ;
      RECT 56.415 0.105 56.585 0.275 ;
      RECT 56.415 8.605 56.585 8.775 ;
      RECT 56.345 2.765 56.515 2.935 ;
      RECT 56.345 5.945 56.515 6.115 ;
      RECT 54.955 1.415 55.125 1.585 ;
      RECT 54.955 4.135 55.125 4.305 ;
      RECT 54.515 2.28 54.685 2.45 ;
      RECT 54.495 1.415 54.665 1.585 ;
      RECT 54.495 4.135 54.665 4.305 ;
      RECT 54.12 3.025 54.29 3.195 ;
      RECT 54.035 1.415 54.205 1.585 ;
      RECT 54.035 4.135 54.205 4.305 ;
      RECT 54.01 2.3 54.18 2.47 ;
      RECT 53.575 1.415 53.745 1.585 ;
      RECT 53.575 4.135 53.745 4.305 ;
      RECT 53.19 1.99 53.36 2.16 ;
      RECT 53.115 1.415 53.285 1.585 ;
      RECT 53.115 4.135 53.285 4.305 ;
      RECT 52.875 3.03 53.045 3.2 ;
      RECT 52.83 2.52 53 2.69 ;
      RECT 52.655 1.415 52.825 1.585 ;
      RECT 52.655 4.135 52.825 4.305 ;
      RECT 52.405 2.73 52.575 2.9 ;
      RECT 52.215 1.95 52.385 2.12 ;
      RECT 52.195 1.415 52.365 1.585 ;
      RECT 52.195 4.135 52.365 4.305 ;
      RECT 52.165 3.56 52.335 3.73 ;
      RECT 51.83 3 52 3.17 ;
      RECT 51.735 1.415 51.905 1.585 ;
      RECT 51.735 2.16 51.905 2.33 ;
      RECT 51.735 4.135 51.905 4.305 ;
      RECT 51.275 1.415 51.445 1.585 ;
      RECT 51.275 4.135 51.445 4.305 ;
      RECT 50.935 3.385 51.105 3.555 ;
      RECT 50.875 2.585 51.045 2.755 ;
      RECT 50.815 1.415 50.985 1.585 ;
      RECT 50.815 4.135 50.985 4.305 ;
      RECT 50.435 2.255 50.605 2.425 ;
      RECT 50.355 1.415 50.525 1.585 ;
      RECT 50.355 4.135 50.525 4.305 ;
      RECT 50.17 3.305 50.34 3.475 ;
      RECT 49.925 2.545 50.095 2.715 ;
      RECT 49.895 1.415 50.065 1.585 ;
      RECT 49.895 4.135 50.065 4.305 ;
      RECT 49.83 3.575 50 3.745 ;
      RECT 49.555 2.27 49.725 2.44 ;
      RECT 49.435 1.415 49.605 1.585 ;
      RECT 49.435 4.135 49.605 4.305 ;
      RECT 49.025 2.47 49.195 2.64 ;
      RECT 48.975 1.415 49.145 1.585 ;
      RECT 48.975 4.135 49.145 4.305 ;
      RECT 48.515 1.415 48.685 1.585 ;
      RECT 48.515 4.135 48.685 4.305 ;
      RECT 48.505 2.415 48.675 2.585 ;
      RECT 48.3 2.015 48.47 2.185 ;
      RECT 48.3 3.595 48.47 3.765 ;
      RECT 48.055 1.415 48.225 1.585 ;
      RECT 48.055 4.135 48.225 4.305 ;
      RECT 47.99 2.56 48.16 2.73 ;
      RECT 47.595 1.415 47.765 1.585 ;
      RECT 47.595 4.135 47.765 4.305 ;
      RECT 47.58 2.785 47.75 2.955 ;
      RECT 47.135 1.415 47.305 1.585 ;
      RECT 47.135 4.135 47.305 4.305 ;
      RECT 46.87 3.085 47.04 3.255 ;
      RECT 46.725 1.995 46.895 2.165 ;
      RECT 46.675 1.415 46.845 1.585 ;
      RECT 46.675 4.135 46.845 4.305 ;
      RECT 45.24 0.915 45.41 1.085 ;
      RECT 45.24 2.395 45.41 2.565 ;
      RECT 45.24 6.315 45.41 6.485 ;
      RECT 45.24 7.795 45.41 7.965 ;
      RECT 44.89 0.105 45.06 0.275 ;
      RECT 44.89 4.165 45.06 4.335 ;
      RECT 44.89 4.545 45.06 4.715 ;
      RECT 44.89 8.605 45.06 8.775 ;
      RECT 44.87 2.765 45.04 2.935 ;
      RECT 44.87 5.945 45.04 6.115 ;
      RECT 44.25 0.915 44.42 1.085 ;
      RECT 44.25 2.395 44.42 2.565 ;
      RECT 44.25 6.315 44.42 6.485 ;
      RECT 44.25 7.795 44.42 7.965 ;
      RECT 43.9 0.105 44.07 0.275 ;
      RECT 43.9 4.165 44.07 4.335 ;
      RECT 43.9 4.545 44.07 4.715 ;
      RECT 43.9 8.605 44.07 8.775 ;
      RECT 43.88 2.765 44.05 2.935 ;
      RECT 43.88 5.945 44.05 6.115 ;
      RECT 43.195 0.105 43.365 0.275 ;
      RECT 43.195 4.165 43.365 4.335 ;
      RECT 43.195 4.545 43.365 4.715 ;
      RECT 43.195 8.605 43.365 8.775 ;
      RECT 42.885 2.025 43.055 2.195 ;
      RECT 42.885 6.685 43.055 6.855 ;
      RECT 42.515 0.105 42.685 0.275 ;
      RECT 42.515 8.605 42.685 8.775 ;
      RECT 42.455 0.915 42.625 1.085 ;
      RECT 42.455 1.655 42.625 1.825 ;
      RECT 42.455 7.055 42.625 7.225 ;
      RECT 42.455 7.795 42.625 7.965 ;
      RECT 42.08 2.395 42.25 2.565 ;
      RECT 42.08 6.315 42.25 6.485 ;
      RECT 41.835 0.105 42.005 0.275 ;
      RECT 41.835 8.605 42.005 8.775 ;
      RECT 41.155 0.105 41.325 0.275 ;
      RECT 41.155 8.605 41.325 8.775 ;
      RECT 41.085 2.765 41.255 2.935 ;
      RECT 41.085 5.945 41.255 6.115 ;
      RECT 39.695 1.415 39.865 1.585 ;
      RECT 39.695 4.135 39.865 4.305 ;
      RECT 39.255 2.28 39.425 2.45 ;
      RECT 39.235 1.415 39.405 1.585 ;
      RECT 39.235 4.135 39.405 4.305 ;
      RECT 38.86 3.025 39.03 3.195 ;
      RECT 38.775 1.415 38.945 1.585 ;
      RECT 38.775 4.135 38.945 4.305 ;
      RECT 38.75 2.3 38.92 2.47 ;
      RECT 38.315 1.415 38.485 1.585 ;
      RECT 38.315 4.135 38.485 4.305 ;
      RECT 37.93 1.99 38.1 2.16 ;
      RECT 37.855 1.415 38.025 1.585 ;
      RECT 37.855 4.135 38.025 4.305 ;
      RECT 37.615 3.03 37.785 3.2 ;
      RECT 37.57 2.52 37.74 2.69 ;
      RECT 37.395 1.415 37.565 1.585 ;
      RECT 37.395 4.135 37.565 4.305 ;
      RECT 37.145 2.73 37.315 2.9 ;
      RECT 36.955 1.95 37.125 2.12 ;
      RECT 36.935 1.415 37.105 1.585 ;
      RECT 36.935 4.135 37.105 4.305 ;
      RECT 36.905 3.56 37.075 3.73 ;
      RECT 36.57 3 36.74 3.17 ;
      RECT 36.475 1.415 36.645 1.585 ;
      RECT 36.475 2.16 36.645 2.33 ;
      RECT 36.475 4.135 36.645 4.305 ;
      RECT 36.015 1.415 36.185 1.585 ;
      RECT 36.015 4.135 36.185 4.305 ;
      RECT 35.675 3.385 35.845 3.555 ;
      RECT 35.615 2.585 35.785 2.755 ;
      RECT 35.555 1.415 35.725 1.585 ;
      RECT 35.555 4.135 35.725 4.305 ;
      RECT 35.175 2.255 35.345 2.425 ;
      RECT 35.095 1.415 35.265 1.585 ;
      RECT 35.095 4.135 35.265 4.305 ;
      RECT 34.91 3.305 35.08 3.475 ;
      RECT 34.665 2.545 34.835 2.715 ;
      RECT 34.635 1.415 34.805 1.585 ;
      RECT 34.635 4.135 34.805 4.305 ;
      RECT 34.57 3.575 34.74 3.745 ;
      RECT 34.295 2.27 34.465 2.44 ;
      RECT 34.175 1.415 34.345 1.585 ;
      RECT 34.175 4.135 34.345 4.305 ;
      RECT 33.765 2.47 33.935 2.64 ;
      RECT 33.715 1.415 33.885 1.585 ;
      RECT 33.715 4.135 33.885 4.305 ;
      RECT 33.255 1.415 33.425 1.585 ;
      RECT 33.255 4.135 33.425 4.305 ;
      RECT 33.245 2.415 33.415 2.585 ;
      RECT 33.04 2.015 33.21 2.185 ;
      RECT 33.04 3.595 33.21 3.765 ;
      RECT 32.795 1.415 32.965 1.585 ;
      RECT 32.795 4.135 32.965 4.305 ;
      RECT 32.73 2.56 32.9 2.73 ;
      RECT 32.335 1.415 32.505 1.585 ;
      RECT 32.335 4.135 32.505 4.305 ;
      RECT 32.32 2.785 32.49 2.955 ;
      RECT 31.875 1.415 32.045 1.585 ;
      RECT 31.875 4.135 32.045 4.305 ;
      RECT 31.61 3.085 31.78 3.255 ;
      RECT 31.465 1.995 31.635 2.165 ;
      RECT 31.415 1.415 31.585 1.585 ;
      RECT 31.415 4.135 31.585 4.305 ;
      RECT 29.98 0.915 30.15 1.085 ;
      RECT 29.98 2.395 30.15 2.565 ;
      RECT 29.98 6.315 30.15 6.485 ;
      RECT 29.98 7.795 30.15 7.965 ;
      RECT 29.63 0.105 29.8 0.275 ;
      RECT 29.63 4.165 29.8 4.335 ;
      RECT 29.63 4.545 29.8 4.715 ;
      RECT 29.63 8.605 29.8 8.775 ;
      RECT 29.61 2.765 29.78 2.935 ;
      RECT 29.61 5.945 29.78 6.115 ;
      RECT 28.99 0.915 29.16 1.085 ;
      RECT 28.99 2.395 29.16 2.565 ;
      RECT 28.99 6.315 29.16 6.485 ;
      RECT 28.99 7.795 29.16 7.965 ;
      RECT 28.64 0.105 28.81 0.275 ;
      RECT 28.64 4.165 28.81 4.335 ;
      RECT 28.64 4.545 28.81 4.715 ;
      RECT 28.64 8.605 28.81 8.775 ;
      RECT 28.62 2.765 28.79 2.935 ;
      RECT 28.62 5.945 28.79 6.115 ;
      RECT 27.935 0.105 28.105 0.275 ;
      RECT 27.935 4.165 28.105 4.335 ;
      RECT 27.935 4.545 28.105 4.715 ;
      RECT 27.935 8.605 28.105 8.775 ;
      RECT 27.625 2.025 27.795 2.195 ;
      RECT 27.625 6.685 27.795 6.855 ;
      RECT 27.255 0.105 27.425 0.275 ;
      RECT 27.255 8.605 27.425 8.775 ;
      RECT 27.195 0.915 27.365 1.085 ;
      RECT 27.195 1.655 27.365 1.825 ;
      RECT 27.195 7.055 27.365 7.225 ;
      RECT 27.195 7.795 27.365 7.965 ;
      RECT 26.82 2.395 26.99 2.565 ;
      RECT 26.82 6.315 26.99 6.485 ;
      RECT 26.575 0.105 26.745 0.275 ;
      RECT 26.575 8.605 26.745 8.775 ;
      RECT 25.895 0.105 26.065 0.275 ;
      RECT 25.895 8.605 26.065 8.775 ;
      RECT 25.825 2.765 25.995 2.935 ;
      RECT 25.825 5.945 25.995 6.115 ;
      RECT 24.435 1.415 24.605 1.585 ;
      RECT 24.435 4.135 24.605 4.305 ;
      RECT 23.995 2.28 24.165 2.45 ;
      RECT 23.975 1.415 24.145 1.585 ;
      RECT 23.975 4.135 24.145 4.305 ;
      RECT 23.6 3.025 23.77 3.195 ;
      RECT 23.515 1.415 23.685 1.585 ;
      RECT 23.515 4.135 23.685 4.305 ;
      RECT 23.49 2.3 23.66 2.47 ;
      RECT 23.055 1.415 23.225 1.585 ;
      RECT 23.055 4.135 23.225 4.305 ;
      RECT 22.67 1.99 22.84 2.16 ;
      RECT 22.595 1.415 22.765 1.585 ;
      RECT 22.595 4.135 22.765 4.305 ;
      RECT 22.355 3.03 22.525 3.2 ;
      RECT 22.31 2.52 22.48 2.69 ;
      RECT 22.135 1.415 22.305 1.585 ;
      RECT 22.135 4.135 22.305 4.305 ;
      RECT 21.885 2.73 22.055 2.9 ;
      RECT 21.695 1.95 21.865 2.12 ;
      RECT 21.675 1.415 21.845 1.585 ;
      RECT 21.675 4.135 21.845 4.305 ;
      RECT 21.645 3.56 21.815 3.73 ;
      RECT 21.31 3 21.48 3.17 ;
      RECT 21.215 1.415 21.385 1.585 ;
      RECT 21.215 2.16 21.385 2.33 ;
      RECT 21.215 4.135 21.385 4.305 ;
      RECT 20.755 1.415 20.925 1.585 ;
      RECT 20.755 4.135 20.925 4.305 ;
      RECT 20.415 3.385 20.585 3.555 ;
      RECT 20.355 2.585 20.525 2.755 ;
      RECT 20.295 1.415 20.465 1.585 ;
      RECT 20.295 4.135 20.465 4.305 ;
      RECT 19.915 2.255 20.085 2.425 ;
      RECT 19.835 1.415 20.005 1.585 ;
      RECT 19.835 4.135 20.005 4.305 ;
      RECT 19.65 3.305 19.82 3.475 ;
      RECT 19.405 2.545 19.575 2.715 ;
      RECT 19.375 1.415 19.545 1.585 ;
      RECT 19.375 4.135 19.545 4.305 ;
      RECT 19.31 3.575 19.48 3.745 ;
      RECT 19.035 2.27 19.205 2.44 ;
      RECT 18.915 1.415 19.085 1.585 ;
      RECT 18.915 4.135 19.085 4.305 ;
      RECT 18.505 2.47 18.675 2.64 ;
      RECT 18.455 1.415 18.625 1.585 ;
      RECT 18.455 4.135 18.625 4.305 ;
      RECT 17.995 1.415 18.165 1.585 ;
      RECT 17.995 4.135 18.165 4.305 ;
      RECT 17.985 2.415 18.155 2.585 ;
      RECT 17.78 2.015 17.95 2.185 ;
      RECT 17.78 3.595 17.95 3.765 ;
      RECT 17.535 1.415 17.705 1.585 ;
      RECT 17.535 4.135 17.705 4.305 ;
      RECT 17.47 2.56 17.64 2.73 ;
      RECT 17.075 1.415 17.245 1.585 ;
      RECT 17.075 4.135 17.245 4.305 ;
      RECT 17.06 2.785 17.23 2.955 ;
      RECT 16.615 1.415 16.785 1.585 ;
      RECT 16.615 4.135 16.785 4.305 ;
      RECT 16.35 3.085 16.52 3.255 ;
      RECT 16.205 1.995 16.375 2.165 ;
      RECT 16.155 1.415 16.325 1.585 ;
      RECT 16.155 4.135 16.325 4.305 ;
      RECT 14.72 0.915 14.89 1.085 ;
      RECT 14.72 2.395 14.89 2.565 ;
      RECT 14.72 6.315 14.89 6.485 ;
      RECT 14.72 7.795 14.89 7.965 ;
      RECT 14.37 0.105 14.54 0.275 ;
      RECT 14.37 4.165 14.54 4.335 ;
      RECT 14.37 4.545 14.54 4.715 ;
      RECT 14.37 8.605 14.54 8.775 ;
      RECT 14.35 2.765 14.52 2.935 ;
      RECT 14.35 5.945 14.52 6.115 ;
      RECT 13.73 0.915 13.9 1.085 ;
      RECT 13.73 2.395 13.9 2.565 ;
      RECT 13.73 6.315 13.9 6.485 ;
      RECT 13.73 7.795 13.9 7.965 ;
      RECT 13.38 0.105 13.55 0.275 ;
      RECT 13.38 4.165 13.55 4.335 ;
      RECT 13.38 4.545 13.55 4.715 ;
      RECT 13.38 8.605 13.55 8.775 ;
      RECT 13.36 2.765 13.53 2.935 ;
      RECT 13.36 5.945 13.53 6.115 ;
      RECT 12.675 0.105 12.845 0.275 ;
      RECT 12.675 4.165 12.845 4.335 ;
      RECT 12.675 4.545 12.845 4.715 ;
      RECT 12.675 8.605 12.845 8.775 ;
      RECT 12.365 2.025 12.535 2.195 ;
      RECT 12.365 6.685 12.535 6.855 ;
      RECT 11.995 0.105 12.165 0.275 ;
      RECT 11.995 8.605 12.165 8.775 ;
      RECT 11.935 0.915 12.105 1.085 ;
      RECT 11.935 1.655 12.105 1.825 ;
      RECT 11.935 7.055 12.105 7.225 ;
      RECT 11.935 7.795 12.105 7.965 ;
      RECT 11.56 2.395 11.73 2.565 ;
      RECT 11.56 6.315 11.73 6.485 ;
      RECT 11.315 0.105 11.485 0.275 ;
      RECT 11.315 8.605 11.485 8.775 ;
      RECT 10.635 0.105 10.805 0.275 ;
      RECT 10.635 8.605 10.805 8.775 ;
      RECT 10.565 2.765 10.735 2.935 ;
      RECT 10.565 5.945 10.735 6.115 ;
      RECT 9.175 1.415 9.345 1.585 ;
      RECT 9.175 4.135 9.345 4.305 ;
      RECT 8.735 2.28 8.905 2.45 ;
      RECT 8.715 1.415 8.885 1.585 ;
      RECT 8.715 4.135 8.885 4.305 ;
      RECT 8.34 3.025 8.51 3.195 ;
      RECT 8.255 1.415 8.425 1.585 ;
      RECT 8.255 4.135 8.425 4.305 ;
      RECT 8.23 2.3 8.4 2.47 ;
      RECT 7.795 1.415 7.965 1.585 ;
      RECT 7.795 4.135 7.965 4.305 ;
      RECT 7.41 1.99 7.58 2.16 ;
      RECT 7.335 1.415 7.505 1.585 ;
      RECT 7.335 4.135 7.505 4.305 ;
      RECT 7.095 3.03 7.265 3.2 ;
      RECT 7.05 2.52 7.22 2.69 ;
      RECT 6.875 1.415 7.045 1.585 ;
      RECT 6.875 4.135 7.045 4.305 ;
      RECT 6.625 2.73 6.795 2.9 ;
      RECT 6.435 1.95 6.605 2.12 ;
      RECT 6.415 1.415 6.585 1.585 ;
      RECT 6.415 4.135 6.585 4.305 ;
      RECT 6.385 3.56 6.555 3.73 ;
      RECT 6.05 3 6.22 3.17 ;
      RECT 5.955 1.415 6.125 1.585 ;
      RECT 5.955 2.16 6.125 2.33 ;
      RECT 5.955 4.135 6.125 4.305 ;
      RECT 5.495 1.415 5.665 1.585 ;
      RECT 5.495 4.135 5.665 4.305 ;
      RECT 5.155 3.385 5.325 3.555 ;
      RECT 5.095 2.585 5.265 2.755 ;
      RECT 5.035 1.415 5.205 1.585 ;
      RECT 5.035 4.135 5.205 4.305 ;
      RECT 4.655 2.255 4.825 2.425 ;
      RECT 4.575 1.415 4.745 1.585 ;
      RECT 4.575 4.135 4.745 4.305 ;
      RECT 4.39 3.305 4.56 3.475 ;
      RECT 4.145 2.545 4.315 2.715 ;
      RECT 4.115 1.415 4.285 1.585 ;
      RECT 4.115 4.135 4.285 4.305 ;
      RECT 4.05 3.575 4.22 3.745 ;
      RECT 3.775 2.27 3.945 2.44 ;
      RECT 3.655 1.415 3.825 1.585 ;
      RECT 3.655 4.135 3.825 4.305 ;
      RECT 3.245 2.47 3.415 2.64 ;
      RECT 3.195 1.415 3.365 1.585 ;
      RECT 3.195 4.135 3.365 4.305 ;
      RECT 2.735 1.415 2.905 1.585 ;
      RECT 2.735 4.135 2.905 4.305 ;
      RECT 2.725 2.415 2.895 2.585 ;
      RECT 2.52 2.015 2.69 2.185 ;
      RECT 2.52 3.595 2.69 3.765 ;
      RECT 2.275 1.415 2.445 1.585 ;
      RECT 2.275 4.135 2.445 4.305 ;
      RECT 2.21 2.56 2.38 2.73 ;
      RECT 1.815 1.415 1.985 1.585 ;
      RECT 1.815 4.135 1.985 4.305 ;
      RECT 1.8 2.785 1.97 2.955 ;
      RECT 1.355 1.415 1.525 1.585 ;
      RECT 1.355 4.135 1.525 4.305 ;
      RECT 1.09 3.085 1.26 3.255 ;
      RECT 0.945 1.995 1.115 2.165 ;
      RECT 0.895 1.415 1.065 1.585 ;
      RECT 0.895 4.135 1.065 4.305 ;
    LAYER li ;
      RECT 69.76 0 69.93 2.085 ;
      RECT 68.82 0 68.99 2.085 ;
      RECT 67.86 0 68.03 2.085 ;
      RECT 65.94 0 66.11 2.085 ;
      RECT 64.98 0 65.15 2.085 ;
      RECT 63.06 0 63.23 2.085 ;
      RECT 54.5 0 54.67 2.085 ;
      RECT 53.56 0 53.73 2.085 ;
      RECT 52.6 0 52.77 2.085 ;
      RECT 50.68 0 50.85 2.085 ;
      RECT 49.72 0 49.89 2.085 ;
      RECT 47.8 0 47.97 2.085 ;
      RECT 39.24 0 39.41 2.085 ;
      RECT 38.3 0 38.47 2.085 ;
      RECT 37.34 0 37.51 2.085 ;
      RECT 35.42 0 35.59 2.085 ;
      RECT 34.46 0 34.63 2.085 ;
      RECT 32.54 0 32.71 2.085 ;
      RECT 23.98 0 24.15 2.085 ;
      RECT 23.04 0 23.21 2.085 ;
      RECT 22.08 0 22.25 2.085 ;
      RECT 20.16 0 20.33 2.085 ;
      RECT 19.2 0 19.37 2.085 ;
      RECT 17.28 0 17.45 2.085 ;
      RECT 8.72 0 8.89 2.085 ;
      RECT 7.78 0 7.95 2.085 ;
      RECT 6.82 0 6.99 2.085 ;
      RECT 4.9 0 5.07 2.085 ;
      RECT 3.94 0 4.11 2.085 ;
      RECT 2.02 0 2.19 2.085 ;
      RECT 66.815 0 67.01 1.595 ;
      RECT 63.06 0 63.335 1.595 ;
      RECT 51.555 0 51.75 1.595 ;
      RECT 47.8 0 48.075 1.595 ;
      RECT 36.295 0 36.49 1.595 ;
      RECT 32.54 0 32.815 1.595 ;
      RECT 21.035 0 21.23 1.595 ;
      RECT 17.28 0 17.555 1.595 ;
      RECT 5.775 0 5.97 1.595 ;
      RECT 2.02 0 2.295 1.595 ;
      RECT 61.79 0 70.53 1.585 ;
      RECT 46.53 0 55.27 1.585 ;
      RECT 31.27 0 40.01 1.585 ;
      RECT 16.01 0 24.75 1.585 ;
      RECT 0.75 0 9.49 1.585 ;
      RECT 75.33 0 75.5 0.935 ;
      RECT 74.34 0 74.51 0.935 ;
      RECT 71.595 0 71.765 0.935 ;
      RECT 60.07 0 60.24 0.935 ;
      RECT 59.08 0 59.25 0.935 ;
      RECT 56.335 0 56.505 0.935 ;
      RECT 44.81 0 44.98 0.935 ;
      RECT 43.82 0 43.99 0.935 ;
      RECT 41.075 0 41.245 0.935 ;
      RECT 29.55 0 29.72 0.935 ;
      RECT 28.56 0 28.73 0.935 ;
      RECT 25.815 0 25.985 0.935 ;
      RECT 14.29 0 14.46 0.935 ;
      RECT 13.3 0 13.47 0.935 ;
      RECT 10.555 0 10.725 0.935 ;
      RECT 0 0 76.3 0.305 ;
      RECT 75.33 3.405 75.5 5.475 ;
      RECT 74.34 3.405 74.51 5.475 ;
      RECT 71.595 3.405 71.765 5.475 ;
      RECT 60.07 3.405 60.24 5.475 ;
      RECT 59.08 3.405 59.25 5.475 ;
      RECT 56.335 3.405 56.505 5.475 ;
      RECT 44.81 3.405 44.98 5.475 ;
      RECT 43.82 3.405 43.99 5.475 ;
      RECT 41.075 3.405 41.245 5.475 ;
      RECT 29.55 3.405 29.72 5.475 ;
      RECT 28.56 3.405 28.73 5.475 ;
      RECT 25.815 3.405 25.985 5.475 ;
      RECT 14.29 3.405 14.46 5.475 ;
      RECT 13.3 3.405 13.47 5.475 ;
      RECT 10.555 3.405 10.725 5.475 ;
      RECT 0 4.14 76.3 4.745 ;
      RECT 61.79 4.135 76.3 4.745 ;
      RECT 46.53 4.135 61.04 4.745 ;
      RECT 31.27 4.135 45.78 4.745 ;
      RECT 16.01 4.135 30.52 4.745 ;
      RECT 0.75 4.135 15.26 4.745 ;
      RECT 68.82 3.635 68.99 4.745 ;
      RECT 66.9 3.635 67.07 4.745 ;
      RECT 65.96 3.635 66.13 4.745 ;
      RECT 64.5 3.635 64.67 4.745 ;
      RECT 62.58 3.635 62.75 4.745 ;
      RECT 53.56 3.635 53.73 4.745 ;
      RECT 51.64 3.635 51.81 4.745 ;
      RECT 50.7 3.635 50.87 4.745 ;
      RECT 49.24 3.635 49.41 4.745 ;
      RECT 47.32 3.635 47.49 4.745 ;
      RECT 38.3 3.635 38.47 4.745 ;
      RECT 36.38 3.635 36.55 4.745 ;
      RECT 35.44 3.635 35.61 4.745 ;
      RECT 33.98 3.635 34.15 4.745 ;
      RECT 32.06 3.635 32.23 4.745 ;
      RECT 23.04 3.635 23.21 4.745 ;
      RECT 21.12 3.635 21.29 4.745 ;
      RECT 20.18 3.635 20.35 4.745 ;
      RECT 18.72 3.635 18.89 4.745 ;
      RECT 16.8 3.635 16.97 4.745 ;
      RECT 7.78 3.635 7.95 4.745 ;
      RECT 5.86 3.635 6.03 4.745 ;
      RECT 4.92 3.635 5.09 4.745 ;
      RECT 3.46 3.635 3.63 4.745 ;
      RECT 1.54 3.635 1.71 4.745 ;
      RECT 0 8.575 76.3 8.88 ;
      RECT 75.33 7.945 75.5 8.88 ;
      RECT 74.34 7.945 74.51 8.88 ;
      RECT 71.595 7.945 71.765 8.88 ;
      RECT 60.07 7.945 60.24 8.88 ;
      RECT 59.08 7.945 59.25 8.88 ;
      RECT 56.335 7.945 56.505 8.88 ;
      RECT 44.81 7.945 44.98 8.88 ;
      RECT 43.82 7.945 43.99 8.88 ;
      RECT 41.075 7.945 41.245 8.88 ;
      RECT 29.55 7.945 29.72 8.88 ;
      RECT 28.56 7.945 28.73 8.88 ;
      RECT 25.815 7.945 25.985 8.88 ;
      RECT 14.29 7.945 14.46 8.88 ;
      RECT 13.3 7.945 13.47 8.88 ;
      RECT 10.555 7.945 10.725 8.88 ;
      RECT 75.39 1.74 75.56 2.935 ;
      RECT 75.39 1.74 75.855 1.91 ;
      RECT 75.39 6.97 75.855 7.14 ;
      RECT 75.39 5.945 75.56 7.14 ;
      RECT 74.4 1.74 74.57 2.935 ;
      RECT 74.4 1.74 74.865 1.91 ;
      RECT 74.4 6.97 74.865 7.14 ;
      RECT 74.4 5.945 74.57 7.14 ;
      RECT 72.545 2.635 72.715 3.865 ;
      RECT 72.6 0.855 72.77 2.805 ;
      RECT 72.545 0.575 72.715 1.025 ;
      RECT 72.545 7.855 72.715 8.305 ;
      RECT 72.6 6.075 72.77 8.025 ;
      RECT 72.545 5.015 72.715 6.245 ;
      RECT 72.025 0.575 72.195 3.865 ;
      RECT 72.025 2.075 72.43 2.405 ;
      RECT 72.025 1.235 72.43 1.565 ;
      RECT 72.025 5.015 72.195 8.305 ;
      RECT 72.025 7.315 72.43 7.645 ;
      RECT 72.025 6.475 72.43 6.805 ;
      RECT 69.95 3.126 69.955 3.298 ;
      RECT 69.945 3.119 69.95 3.388 ;
      RECT 69.94 3.113 69.945 3.407 ;
      RECT 69.92 3.107 69.94 3.417 ;
      RECT 69.905 3.102 69.92 3.425 ;
      RECT 69.868 3.096 69.905 3.423 ;
      RECT 69.782 3.082 69.868 3.419 ;
      RECT 69.696 3.064 69.782 3.414 ;
      RECT 69.61 3.045 69.696 3.408 ;
      RECT 69.58 3.033 69.61 3.404 ;
      RECT 69.56 3.027 69.58 3.403 ;
      RECT 69.495 3.025 69.56 3.401 ;
      RECT 69.48 3.025 69.495 3.393 ;
      RECT 69.465 3.025 69.48 3.38 ;
      RECT 69.46 3.025 69.465 3.37 ;
      RECT 69.445 3.025 69.46 3.348 ;
      RECT 69.43 3.025 69.445 3.315 ;
      RECT 69.425 3.025 69.43 3.293 ;
      RECT 69.415 3.025 69.425 3.275 ;
      RECT 69.4 3.025 69.415 3.253 ;
      RECT 69.38 3.025 69.4 3.215 ;
      RECT 69.73 2.31 69.765 2.749 ;
      RECT 69.73 2.31 69.77 2.748 ;
      RECT 69.675 2.37 69.77 2.747 ;
      RECT 69.54 2.542 69.77 2.746 ;
      RECT 69.65 2.42 69.77 2.746 ;
      RECT 69.54 2.542 69.795 2.736 ;
      RECT 69.595 2.487 69.875 2.653 ;
      RECT 69.77 2.281 69.775 2.744 ;
      RECT 69.625 2.457 69.915 2.53 ;
      RECT 69.64 2.44 69.77 2.746 ;
      RECT 69.775 2.28 69.945 2.468 ;
      RECT 69.765 2.283 69.945 2.468 ;
      RECT 69.27 2.16 69.44 2.47 ;
      RECT 69.27 2.16 69.445 2.443 ;
      RECT 69.27 2.16 69.45 2.42 ;
      RECT 69.27 2.16 69.46 2.37 ;
      RECT 69.265 2.265 69.46 2.34 ;
      RECT 69.3 1.835 69.47 2.313 ;
      RECT 69.3 1.835 69.485 2.234 ;
      RECT 69.29 2.045 69.485 2.234 ;
      RECT 69.3 1.845 69.495 2.149 ;
      RECT 69.23 2.587 69.235 2.79 ;
      RECT 69.22 2.575 69.23 2.9 ;
      RECT 69.195 2.575 69.22 2.94 ;
      RECT 69.115 2.575 69.195 3.025 ;
      RECT 69.105 2.575 69.115 3.095 ;
      RECT 69.08 2.575 69.105 3.118 ;
      RECT 69.06 2.575 69.08 3.153 ;
      RECT 69.015 2.585 69.06 3.196 ;
      RECT 69.005 2.597 69.015 3.233 ;
      RECT 68.985 2.611 69.005 3.253 ;
      RECT 68.975 2.629 68.985 3.269 ;
      RECT 68.96 2.655 68.975 3.279 ;
      RECT 68.945 2.696 68.96 3.293 ;
      RECT 68.935 2.731 68.945 3.303 ;
      RECT 68.93 2.747 68.935 3.308 ;
      RECT 68.92 2.762 68.93 3.313 ;
      RECT 68.9 2.805 68.92 3.323 ;
      RECT 68.88 2.842 68.9 3.336 ;
      RECT 68.845 2.865 68.88 3.354 ;
      RECT 68.835 2.879 68.845 3.37 ;
      RECT 68.815 2.889 68.835 3.38 ;
      RECT 68.81 2.898 68.815 3.388 ;
      RECT 68.8 2.905 68.81 3.395 ;
      RECT 68.79 2.912 68.8 3.403 ;
      RECT 68.775 2.922 68.79 3.411 ;
      RECT 68.765 2.936 68.775 3.421 ;
      RECT 68.755 2.948 68.765 3.433 ;
      RECT 68.74 2.97 68.755 3.446 ;
      RECT 68.73 2.992 68.74 3.457 ;
      RECT 68.72 3.012 68.73 3.466 ;
      RECT 68.715 3.027 68.72 3.473 ;
      RECT 68.685 3.06 68.715 3.487 ;
      RECT 68.675 3.095 68.685 3.502 ;
      RECT 68.67 3.102 68.675 3.508 ;
      RECT 68.65 3.117 68.67 3.515 ;
      RECT 68.645 3.132 68.65 3.523 ;
      RECT 68.64 3.141 68.645 3.528 ;
      RECT 68.625 3.147 68.64 3.535 ;
      RECT 68.62 3.153 68.625 3.543 ;
      RECT 68.615 3.157 68.62 3.55 ;
      RECT 68.61 3.161 68.615 3.56 ;
      RECT 68.6 3.166 68.61 3.57 ;
      RECT 68.58 3.177 68.6 3.598 ;
      RECT 68.565 3.189 68.58 3.625 ;
      RECT 68.545 3.202 68.565 3.65 ;
      RECT 68.525 3.217 68.545 3.674 ;
      RECT 68.51 3.232 68.525 3.689 ;
      RECT 68.505 3.243 68.51 3.698 ;
      RECT 68.44 3.288 68.505 3.708 ;
      RECT 68.405 3.347 68.44 3.721 ;
      RECT 68.4 3.37 68.405 3.727 ;
      RECT 68.395 3.377 68.4 3.729 ;
      RECT 68.38 3.387 68.395 3.732 ;
      RECT 68.35 3.412 68.38 3.736 ;
      RECT 68.345 3.43 68.35 3.74 ;
      RECT 68.34 3.437 68.345 3.741 ;
      RECT 68.32 3.445 68.34 3.745 ;
      RECT 68.31 3.452 68.32 3.749 ;
      RECT 68.266 3.463 68.31 3.756 ;
      RECT 68.18 3.491 68.266 3.772 ;
      RECT 68.12 3.515 68.18 3.79 ;
      RECT 68.075 3.525 68.12 3.804 ;
      RECT 68.016 3.533 68.075 3.818 ;
      RECT 67.93 3.54 68.016 3.837 ;
      RECT 67.905 3.545 67.93 3.852 ;
      RECT 67.825 3.548 67.905 3.855 ;
      RECT 67.745 3.552 67.825 3.842 ;
      RECT 67.736 3.555 67.745 3.827 ;
      RECT 67.65 3.555 67.736 3.812 ;
      RECT 67.59 3.557 67.65 3.789 ;
      RECT 67.586 3.56 67.59 3.779 ;
      RECT 67.5 3.56 67.586 3.764 ;
      RECT 67.425 3.56 67.5 3.74 ;
      RECT 68.74 2.569 68.75 2.745 ;
      RECT 68.695 2.536 68.74 2.745 ;
      RECT 68.65 2.487 68.695 2.745 ;
      RECT 68.62 2.457 68.65 2.746 ;
      RECT 68.615 2.44 68.62 2.747 ;
      RECT 68.59 2.42 68.615 2.748 ;
      RECT 68.575 2.395 68.59 2.749 ;
      RECT 68.57 2.382 68.575 2.75 ;
      RECT 68.565 2.376 68.57 2.748 ;
      RECT 68.56 2.368 68.565 2.742 ;
      RECT 68.535 2.36 68.56 2.722 ;
      RECT 68.515 2.349 68.535 2.693 ;
      RECT 68.485 2.334 68.515 2.664 ;
      RECT 68.465 2.32 68.485 2.636 ;
      RECT 68.455 2.314 68.465 2.615 ;
      RECT 68.45 2.311 68.455 2.598 ;
      RECT 68.445 2.308 68.45 2.583 ;
      RECT 68.43 2.303 68.445 2.548 ;
      RECT 68.425 2.299 68.43 2.515 ;
      RECT 68.405 2.294 68.425 2.491 ;
      RECT 68.375 2.286 68.405 2.456 ;
      RECT 68.36 2.28 68.375 2.433 ;
      RECT 68.32 2.273 68.36 2.418 ;
      RECT 68.295 2.265 68.32 2.398 ;
      RECT 68.275 2.26 68.295 2.388 ;
      RECT 68.24 2.254 68.275 2.383 ;
      RECT 68.195 2.245 68.24 2.382 ;
      RECT 68.165 2.241 68.195 2.384 ;
      RECT 68.08 2.249 68.165 2.388 ;
      RECT 68.01 2.26 68.08 2.41 ;
      RECT 67.997 2.266 68.01 2.433 ;
      RECT 67.911 2.273 67.997 2.455 ;
      RECT 67.825 2.285 67.911 2.492 ;
      RECT 67.825 2.662 67.835 2.9 ;
      RECT 67.82 2.291 67.825 2.515 ;
      RECT 67.815 2.547 67.825 2.9 ;
      RECT 67.815 2.292 67.82 2.52 ;
      RECT 67.81 2.293 67.815 2.9 ;
      RECT 67.786 2.295 67.81 2.901 ;
      RECT 67.7 2.303 67.786 2.903 ;
      RECT 67.68 2.317 67.7 2.906 ;
      RECT 67.675 2.345 67.68 2.907 ;
      RECT 67.67 2.357 67.675 2.908 ;
      RECT 67.665 2.372 67.67 2.909 ;
      RECT 67.655 2.402 67.665 2.91 ;
      RECT 67.65 2.44 67.655 2.908 ;
      RECT 67.645 2.46 67.65 2.903 ;
      RECT 67.63 2.495 67.645 2.888 ;
      RECT 67.62 2.547 67.63 2.868 ;
      RECT 67.615 2.577 67.62 2.856 ;
      RECT 67.6 2.59 67.615 2.839 ;
      RECT 67.575 2.594 67.6 2.806 ;
      RECT 67.56 2.592 67.575 2.783 ;
      RECT 67.545 2.591 67.56 2.78 ;
      RECT 67.485 2.589 67.545 2.778 ;
      RECT 67.475 2.587 67.485 2.773 ;
      RECT 67.435 2.586 67.475 2.77 ;
      RECT 67.365 2.583 67.435 2.768 ;
      RECT 67.31 2.581 67.365 2.763 ;
      RECT 67.24 2.575 67.31 2.758 ;
      RECT 67.231 2.575 67.24 2.755 ;
      RECT 67.145 2.575 67.231 2.75 ;
      RECT 67.14 2.575 67.145 2.745 ;
      RECT 68.445 1.81 68.62 2.16 ;
      RECT 68.445 1.825 68.63 2.158 ;
      RECT 68.42 1.775 68.565 2.155 ;
      RECT 68.4 1.776 68.565 2.148 ;
      RECT 68.39 1.777 68.575 2.143 ;
      RECT 68.36 1.778 68.575 2.13 ;
      RECT 68.31 1.779 68.575 2.106 ;
      RECT 68.305 1.781 68.575 2.091 ;
      RECT 68.305 1.847 68.635 2.085 ;
      RECT 68.285 1.788 68.59 2.065 ;
      RECT 68.275 1.797 68.6 1.92 ;
      RECT 68.285 1.792 68.6 2.065 ;
      RECT 68.305 1.782 68.59 2.091 ;
      RECT 67.89 3.107 68.06 3.395 ;
      RECT 67.885 3.125 68.07 3.39 ;
      RECT 67.85 3.133 68.135 3.31 ;
      RECT 67.85 3.133 68.221 3.3 ;
      RECT 67.85 3.133 68.275 3.246 ;
      RECT 68.135 3.03 68.305 3.214 ;
      RECT 67.85 3.185 68.31 3.202 ;
      RECT 67.835 3.155 68.305 3.198 ;
      RECT 68.095 3.037 68.135 3.349 ;
      RECT 67.975 3.074 68.305 3.214 ;
      RECT 68.07 3.049 68.095 3.375 ;
      RECT 68.06 3.056 68.305 3.214 ;
      RECT 68.191 2.52 68.26 2.779 ;
      RECT 68.191 2.575 68.265 2.778 ;
      RECT 68.105 2.575 68.265 2.777 ;
      RECT 68.1 2.575 68.27 2.77 ;
      RECT 68.09 2.52 68.26 2.765 ;
      RECT 67.47 1.819 67.645 2.12 ;
      RECT 67.455 1.807 67.47 2.105 ;
      RECT 67.425 1.806 67.455 2.058 ;
      RECT 67.425 1.824 67.65 2.053 ;
      RECT 67.41 1.808 67.47 2.018 ;
      RECT 67.405 1.83 67.66 1.918 ;
      RECT 67.405 1.813 67.556 1.918 ;
      RECT 67.405 1.815 67.56 1.918 ;
      RECT 67.41 1.811 67.556 2.018 ;
      RECT 67.515 3.047 67.52 3.395 ;
      RECT 67.505 3.037 67.515 3.401 ;
      RECT 67.47 3.027 67.505 3.403 ;
      RECT 67.432 3.022 67.47 3.407 ;
      RECT 67.346 3.015 67.432 3.414 ;
      RECT 67.26 3.005 67.346 3.424 ;
      RECT 67.215 3 67.26 3.432 ;
      RECT 67.211 3 67.215 3.436 ;
      RECT 67.125 3 67.211 3.443 ;
      RECT 67.11 3 67.125 3.443 ;
      RECT 67.1 2.998 67.11 3.415 ;
      RECT 67.09 2.994 67.1 3.358 ;
      RECT 67.07 2.988 67.09 3.29 ;
      RECT 67.065 2.984 67.07 3.238 ;
      RECT 67.055 2.983 67.065 3.205 ;
      RECT 67.005 2.981 67.055 3.19 ;
      RECT 66.98 2.979 67.005 3.185 ;
      RECT 66.937 2.977 66.98 3.181 ;
      RECT 66.851 2.973 66.937 3.169 ;
      RECT 66.765 2.968 66.851 3.153 ;
      RECT 66.735 2.965 66.765 3.14 ;
      RECT 66.71 2.964 66.735 3.128 ;
      RECT 66.705 2.964 66.71 3.118 ;
      RECT 66.665 2.963 66.705 3.11 ;
      RECT 66.65 2.962 66.665 3.103 ;
      RECT 66.6 2.961 66.65 3.095 ;
      RECT 66.598 2.96 66.6 3.09 ;
      RECT 66.512 2.958 66.598 3.09 ;
      RECT 66.426 2.953 66.512 3.09 ;
      RECT 66.34 2.949 66.426 3.09 ;
      RECT 66.291 2.945 66.34 3.088 ;
      RECT 66.205 2.942 66.291 3.083 ;
      RECT 66.182 2.939 66.205 3.079 ;
      RECT 66.096 2.936 66.182 3.074 ;
      RECT 66.01 2.932 66.096 3.065 ;
      RECT 65.985 2.925 66.01 3.06 ;
      RECT 65.925 2.89 65.985 3.057 ;
      RECT 65.905 2.815 65.925 3.054 ;
      RECT 65.9 2.757 65.905 3.053 ;
      RECT 65.875 2.697 65.9 3.052 ;
      RECT 65.8 2.575 65.875 3.048 ;
      RECT 65.79 2.575 65.8 3.04 ;
      RECT 65.775 2.575 65.79 3.03 ;
      RECT 65.76 2.575 65.775 3 ;
      RECT 65.745 2.575 65.76 2.945 ;
      RECT 65.73 2.575 65.745 2.883 ;
      RECT 65.705 2.575 65.73 2.808 ;
      RECT 65.7 2.575 65.705 2.758 ;
      RECT 67.045 2.12 67.065 2.429 ;
      RECT 67.031 2.122 67.08 2.426 ;
      RECT 67.031 2.127 67.1 2.417 ;
      RECT 66.945 2.125 67.08 2.411 ;
      RECT 66.945 2.133 67.135 2.394 ;
      RECT 66.91 2.135 67.135 2.393 ;
      RECT 66.88 2.143 67.135 2.384 ;
      RECT 66.87 2.148 67.155 2.37 ;
      RECT 66.91 2.138 67.155 2.37 ;
      RECT 66.91 2.141 67.165 2.358 ;
      RECT 66.88 2.143 67.175 2.345 ;
      RECT 66.88 2.147 67.185 2.288 ;
      RECT 66.87 2.152 67.19 2.203 ;
      RECT 67.031 2.12 67.065 2.426 ;
      RECT 66.47 2.223 66.475 2.435 ;
      RECT 66.345 2.22 66.36 2.435 ;
      RECT 65.81 2.25 65.88 2.435 ;
      RECT 65.695 2.25 65.73 2.43 ;
      RECT 66.816 2.552 66.835 2.746 ;
      RECT 66.73 2.507 66.816 2.747 ;
      RECT 66.72 2.46 66.73 2.749 ;
      RECT 66.715 2.44 66.72 2.75 ;
      RECT 66.695 2.405 66.715 2.751 ;
      RECT 66.68 2.355 66.695 2.752 ;
      RECT 66.66 2.292 66.68 2.753 ;
      RECT 66.65 2.255 66.66 2.754 ;
      RECT 66.635 2.244 66.65 2.755 ;
      RECT 66.63 2.236 66.635 2.753 ;
      RECT 66.62 2.235 66.63 2.745 ;
      RECT 66.59 2.232 66.62 2.724 ;
      RECT 66.515 2.227 66.59 2.669 ;
      RECT 66.5 2.223 66.515 2.615 ;
      RECT 66.49 2.223 66.5 2.51 ;
      RECT 66.475 2.223 66.49 2.443 ;
      RECT 66.46 2.223 66.47 2.433 ;
      RECT 66.405 2.222 66.46 2.43 ;
      RECT 66.36 2.22 66.405 2.433 ;
      RECT 66.332 2.22 66.345 2.436 ;
      RECT 66.246 2.224 66.332 2.438 ;
      RECT 66.16 2.23 66.246 2.443 ;
      RECT 66.14 2.234 66.16 2.445 ;
      RECT 66.138 2.235 66.14 2.444 ;
      RECT 66.052 2.237 66.138 2.443 ;
      RECT 65.966 2.242 66.052 2.44 ;
      RECT 65.88 2.247 65.966 2.437 ;
      RECT 65.73 2.25 65.81 2.433 ;
      RECT 66.506 3.225 66.555 3.559 ;
      RECT 66.506 3.225 66.56 3.558 ;
      RECT 66.42 3.225 66.56 3.557 ;
      RECT 66.195 3.333 66.565 3.555 ;
      RECT 66.42 3.225 66.59 3.548 ;
      RECT 66.39 3.237 66.595 3.539 ;
      RECT 66.375 3.255 66.6 3.536 ;
      RECT 66.19 3.339 66.6 3.463 ;
      RECT 66.185 3.346 66.6 3.423 ;
      RECT 66.2 3.312 66.6 3.536 ;
      RECT 66.361 3.258 66.565 3.555 ;
      RECT 66.275 3.278 66.6 3.536 ;
      RECT 66.375 3.252 66.595 3.539 ;
      RECT 66.145 2.576 66.335 2.77 ;
      RECT 66.14 2.578 66.335 2.769 ;
      RECT 66.135 2.582 66.35 2.766 ;
      RECT 66.15 2.575 66.35 2.766 ;
      RECT 66.135 2.685 66.355 2.761 ;
      RECT 65.43 3.185 65.521 3.483 ;
      RECT 65.425 3.187 65.6 3.478 ;
      RECT 65.43 3.185 65.6 3.478 ;
      RECT 65.425 3.191 65.62 3.476 ;
      RECT 65.425 3.246 65.66 3.475 ;
      RECT 65.425 3.281 65.675 3.469 ;
      RECT 65.425 3.315 65.685 3.459 ;
      RECT 65.415 3.195 65.62 3.31 ;
      RECT 65.415 3.215 65.635 3.31 ;
      RECT 65.415 3.198 65.625 3.31 ;
      RECT 65.64 1.966 65.645 2.028 ;
      RECT 65.635 1.888 65.64 2.051 ;
      RECT 65.63 1.845 65.635 2.062 ;
      RECT 65.625 1.835 65.63 2.074 ;
      RECT 65.62 1.835 65.625 2.083 ;
      RECT 65.595 1.835 65.62 2.115 ;
      RECT 65.59 1.835 65.595 2.148 ;
      RECT 65.575 1.835 65.59 2.173 ;
      RECT 65.565 1.835 65.575 2.2 ;
      RECT 65.56 1.835 65.565 2.213 ;
      RECT 65.555 1.835 65.56 2.228 ;
      RECT 65.545 1.835 65.555 2.243 ;
      RECT 65.54 1.835 65.545 2.263 ;
      RECT 65.515 1.835 65.54 2.298 ;
      RECT 65.47 1.835 65.515 2.343 ;
      RECT 65.46 1.835 65.47 2.356 ;
      RECT 65.375 1.92 65.46 2.363 ;
      RECT 65.34 2.042 65.375 2.372 ;
      RECT 65.335 2.082 65.34 2.376 ;
      RECT 65.315 2.105 65.335 2.378 ;
      RECT 65.31 2.135 65.315 2.381 ;
      RECT 65.3 2.147 65.31 2.382 ;
      RECT 65.255 2.17 65.3 2.387 ;
      RECT 65.215 2.2 65.255 2.395 ;
      RECT 65.18 2.212 65.215 2.401 ;
      RECT 65.175 2.217 65.18 2.405 ;
      RECT 65.105 2.227 65.175 2.412 ;
      RECT 65.065 2.237 65.105 2.422 ;
      RECT 65.045 2.242 65.065 2.428 ;
      RECT 65.035 2.246 65.045 2.433 ;
      RECT 65.03 2.249 65.035 2.436 ;
      RECT 65.02 2.25 65.03 2.437 ;
      RECT 64.995 2.252 65.02 2.441 ;
      RECT 64.985 2.257 64.995 2.444 ;
      RECT 64.94 2.265 64.985 2.445 ;
      RECT 64.815 2.27 64.94 2.445 ;
      RECT 65.37 2.567 65.39 2.749 ;
      RECT 65.321 2.552 65.37 2.748 ;
      RECT 65.235 2.567 65.39 2.746 ;
      RECT 65.22 2.567 65.39 2.745 ;
      RECT 65.185 2.545 65.355 2.73 ;
      RECT 65.255 3.565 65.27 3.774 ;
      RECT 65.255 3.573 65.275 3.773 ;
      RECT 65.2 3.573 65.275 3.772 ;
      RECT 65.18 3.577 65.28 3.77 ;
      RECT 65.16 3.527 65.2 3.769 ;
      RECT 65.105 3.585 65.285 3.767 ;
      RECT 65.07 3.542 65.2 3.765 ;
      RECT 65.066 3.545 65.255 3.764 ;
      RECT 64.98 3.553 65.255 3.762 ;
      RECT 64.98 3.597 65.29 3.755 ;
      RECT 64.97 3.69 65.29 3.753 ;
      RECT 64.98 3.609 65.295 3.738 ;
      RECT 64.98 3.63 65.31 3.708 ;
      RECT 64.98 3.657 65.315 3.678 ;
      RECT 65.105 3.535 65.2 3.767 ;
      RECT 64.735 2.58 64.74 3.118 ;
      RECT 64.54 2.91 64.545 3.105 ;
      RECT 62.84 2.575 62.855 2.955 ;
      RECT 64.905 2.575 64.91 2.745 ;
      RECT 64.9 2.575 64.905 2.755 ;
      RECT 64.895 2.575 64.9 2.768 ;
      RECT 64.87 2.575 64.895 2.81 ;
      RECT 64.845 2.575 64.87 2.883 ;
      RECT 64.83 2.575 64.845 2.935 ;
      RECT 64.825 2.575 64.83 2.965 ;
      RECT 64.8 2.575 64.825 3.005 ;
      RECT 64.785 2.575 64.8 3.06 ;
      RECT 64.78 2.575 64.785 3.093 ;
      RECT 64.755 2.575 64.78 3.113 ;
      RECT 64.74 2.575 64.755 3.119 ;
      RECT 64.67 2.61 64.735 3.115 ;
      RECT 64.62 2.665 64.67 3.11 ;
      RECT 64.61 2.697 64.62 3.108 ;
      RECT 64.605 2.722 64.61 3.108 ;
      RECT 64.585 2.795 64.605 3.108 ;
      RECT 64.575 2.875 64.585 3.107 ;
      RECT 64.56 2.905 64.575 3.107 ;
      RECT 64.545 2.91 64.56 3.106 ;
      RECT 64.485 2.912 64.54 3.103 ;
      RECT 64.455 2.917 64.485 3.099 ;
      RECT 64.453 2.92 64.455 3.098 ;
      RECT 64.367 2.922 64.453 3.095 ;
      RECT 64.281 2.928 64.367 3.089 ;
      RECT 64.195 2.933 64.281 3.083 ;
      RECT 64.122 2.938 64.195 3.084 ;
      RECT 64.036 2.944 64.122 3.092 ;
      RECT 63.95 2.95 64.036 3.101 ;
      RECT 63.93 2.954 63.95 3.106 ;
      RECT 63.883 2.956 63.93 3.109 ;
      RECT 63.797 2.961 63.883 3.115 ;
      RECT 63.711 2.966 63.797 3.124 ;
      RECT 63.625 2.972 63.711 3.132 ;
      RECT 63.54 2.97 63.625 3.141 ;
      RECT 63.536 2.965 63.54 3.145 ;
      RECT 63.45 2.96 63.536 3.137 ;
      RECT 63.386 2.951 63.45 3.125 ;
      RECT 63.3 2.942 63.386 3.112 ;
      RECT 63.276 2.935 63.3 3.103 ;
      RECT 63.19 2.929 63.276 3.09 ;
      RECT 63.15 2.922 63.19 3.076 ;
      RECT 63.145 2.912 63.15 3.072 ;
      RECT 63.135 2.9 63.145 3.071 ;
      RECT 63.115 2.87 63.135 3.068 ;
      RECT 63.06 2.79 63.115 3.062 ;
      RECT 63.04 2.709 63.06 3.057 ;
      RECT 63.02 2.667 63.04 3.053 ;
      RECT 62.995 2.62 63.02 3.047 ;
      RECT 62.99 2.595 62.995 3.044 ;
      RECT 62.955 2.575 62.99 3.039 ;
      RECT 62.946 2.575 62.955 3.032 ;
      RECT 62.86 2.575 62.946 3.002 ;
      RECT 62.855 2.575 62.86 2.965 ;
      RECT 62.82 2.575 62.84 2.887 ;
      RECT 62.815 2.617 62.82 2.852 ;
      RECT 62.81 2.692 62.815 2.808 ;
      RECT 64.26 2.497 64.435 2.745 ;
      RECT 64.26 2.497 64.44 2.743 ;
      RECT 64.255 2.529 64.44 2.703 ;
      RECT 64.285 2.47 64.455 2.69 ;
      RECT 64.25 2.547 64.455 2.623 ;
      RECT 63.56 2.01 63.73 2.185 ;
      RECT 63.56 2.01 63.902 2.177 ;
      RECT 63.56 2.01 63.985 2.171 ;
      RECT 63.56 2.01 64.02 2.167 ;
      RECT 63.56 2.01 64.04 2.166 ;
      RECT 63.56 2.01 64.126 2.162 ;
      RECT 64.02 1.835 64.19 2.157 ;
      RECT 63.595 1.942 64.22 2.155 ;
      RECT 63.585 1.997 64.225 2.153 ;
      RECT 63.56 2.033 64.235 2.148 ;
      RECT 63.56 2.06 64.24 2.078 ;
      RECT 63.625 1.885 64.2 2.155 ;
      RECT 63.816 1.87 64.2 2.155 ;
      RECT 63.65 1.873 64.2 2.155 ;
      RECT 63.73 1.871 63.816 2.182 ;
      RECT 63.816 1.868 64.195 2.155 ;
      RECT 64 1.845 64.195 2.155 ;
      RECT 63.902 1.866 64.195 2.155 ;
      RECT 63.985 1.86 64 2.168 ;
      RECT 64.135 3.225 64.14 3.425 ;
      RECT 63.6 3.29 63.645 3.425 ;
      RECT 64.17 3.225 64.19 3.398 ;
      RECT 64.14 3.225 64.17 3.413 ;
      RECT 64.075 3.225 64.135 3.45 ;
      RECT 64.06 3.225 64.075 3.48 ;
      RECT 64.045 3.225 64.06 3.493 ;
      RECT 64.025 3.225 64.045 3.508 ;
      RECT 64.02 3.225 64.025 3.517 ;
      RECT 64.01 3.229 64.02 3.522 ;
      RECT 63.995 3.239 64.01 3.533 ;
      RECT 63.97 3.255 63.995 3.543 ;
      RECT 63.96 3.269 63.97 3.545 ;
      RECT 63.94 3.281 63.96 3.542 ;
      RECT 63.91 3.302 63.94 3.536 ;
      RECT 63.9 3.314 63.91 3.531 ;
      RECT 63.89 3.312 63.9 3.528 ;
      RECT 63.875 3.311 63.89 3.523 ;
      RECT 63.87 3.31 63.875 3.518 ;
      RECT 63.835 3.308 63.87 3.508 ;
      RECT 63.815 3.305 63.835 3.49 ;
      RECT 63.805 3.303 63.815 3.485 ;
      RECT 63.795 3.302 63.805 3.48 ;
      RECT 63.76 3.3 63.795 3.468 ;
      RECT 63.705 3.296 63.76 3.448 ;
      RECT 63.695 3.294 63.705 3.433 ;
      RECT 63.69 3.294 63.695 3.428 ;
      RECT 63.645 3.292 63.69 3.425 ;
      RECT 63.55 3.29 63.6 3.429 ;
      RECT 63.54 3.291 63.55 3.434 ;
      RECT 63.48 3.298 63.54 3.448 ;
      RECT 63.455 3.306 63.48 3.468 ;
      RECT 63.445 3.31 63.455 3.48 ;
      RECT 63.44 3.311 63.445 3.485 ;
      RECT 63.425 3.313 63.44 3.488 ;
      RECT 63.41 3.315 63.425 3.493 ;
      RECT 63.405 3.315 63.41 3.496 ;
      RECT 63.36 3.32 63.405 3.507 ;
      RECT 63.355 3.324 63.36 3.519 ;
      RECT 63.33 3.32 63.355 3.523 ;
      RECT 63.32 3.316 63.33 3.527 ;
      RECT 63.31 3.315 63.32 3.531 ;
      RECT 63.295 3.305 63.31 3.537 ;
      RECT 63.29 3.293 63.295 3.541 ;
      RECT 63.285 3.29 63.29 3.542 ;
      RECT 63.28 3.287 63.285 3.544 ;
      RECT 63.265 3.275 63.28 3.543 ;
      RECT 63.25 3.257 63.265 3.54 ;
      RECT 63.23 3.236 63.25 3.533 ;
      RECT 63.165 3.225 63.23 3.505 ;
      RECT 63.161 3.225 63.165 3.484 ;
      RECT 63.075 3.225 63.161 3.454 ;
      RECT 63.06 3.225 63.075 3.41 ;
      RECT 63.635 2.325 63.64 2.56 ;
      RECT 62.765 2.241 62.77 2.445 ;
      RECT 63.345 2.27 63.35 2.425 ;
      RECT 63.265 2.25 63.27 2.425 ;
      RECT 63.935 2.392 63.95 2.745 ;
      RECT 63.861 2.377 63.935 2.745 ;
      RECT 63.775 2.36 63.861 2.745 ;
      RECT 63.765 2.35 63.775 2.743 ;
      RECT 63.76 2.348 63.765 2.738 ;
      RECT 63.745 2.346 63.76 2.724 ;
      RECT 63.675 2.338 63.745 2.664 ;
      RECT 63.655 2.329 63.675 2.598 ;
      RECT 63.65 2.326 63.655 2.578 ;
      RECT 63.64 2.325 63.65 2.568 ;
      RECT 63.63 2.325 63.635 2.552 ;
      RECT 63.62 2.324 63.63 2.542 ;
      RECT 63.61 2.322 63.62 2.53 ;
      RECT 63.595 2.319 63.61 2.51 ;
      RECT 63.585 2.317 63.595 2.495 ;
      RECT 63.565 2.314 63.585 2.483 ;
      RECT 63.56 2.312 63.565 2.473 ;
      RECT 63.535 2.31 63.56 2.46 ;
      RECT 63.505 2.305 63.535 2.445 ;
      RECT 63.425 2.296 63.505 2.436 ;
      RECT 63.38 2.285 63.425 2.429 ;
      RECT 63.36 2.276 63.38 2.426 ;
      RECT 63.35 2.271 63.36 2.425 ;
      RECT 63.305 2.265 63.345 2.425 ;
      RECT 63.29 2.257 63.305 2.425 ;
      RECT 63.27 2.252 63.29 2.425 ;
      RECT 63.25 2.249 63.265 2.425 ;
      RECT 63.167 2.248 63.25 2.424 ;
      RECT 63.081 2.247 63.167 2.42 ;
      RECT 62.995 2.245 63.081 2.417 ;
      RECT 62.942 2.244 62.995 2.419 ;
      RECT 62.856 2.243 62.942 2.428 ;
      RECT 62.77 2.242 62.856 2.44 ;
      RECT 62.75 2.241 62.765 2.448 ;
      RECT 62.67 2.24 62.75 2.46 ;
      RECT 62.645 2.24 62.67 2.473 ;
      RECT 62.62 2.24 62.645 2.488 ;
      RECT 62.615 2.24 62.62 2.51 ;
      RECT 62.61 2.24 62.615 2.528 ;
      RECT 62.605 2.24 62.61 2.545 ;
      RECT 62.6 2.24 62.605 2.558 ;
      RECT 62.595 2.24 62.6 2.568 ;
      RECT 62.555 2.24 62.595 2.653 ;
      RECT 62.54 2.24 62.555 2.738 ;
      RECT 62.53 2.241 62.54 2.75 ;
      RECT 62.495 2.246 62.53 2.755 ;
      RECT 62.455 2.255 62.495 2.755 ;
      RECT 62.44 2.265 62.455 2.755 ;
      RECT 62.435 2.275 62.44 2.755 ;
      RECT 62.415 2.302 62.435 2.755 ;
      RECT 62.365 2.385 62.415 2.755 ;
      RECT 62.36 2.447 62.365 2.755 ;
      RECT 62.35 2.46 62.36 2.755 ;
      RECT 62.34 2.482 62.35 2.755 ;
      RECT 62.33 2.507 62.34 2.75 ;
      RECT 62.325 2.545 62.33 2.743 ;
      RECT 62.315 2.655 62.325 2.738 ;
      RECT 63.71 3.576 63.725 3.835 ;
      RECT 63.71 3.591 63.73 3.834 ;
      RECT 63.626 3.591 63.73 3.832 ;
      RECT 63.626 3.605 63.735 3.831 ;
      RECT 63.54 3.647 63.74 3.828 ;
      RECT 63.535 3.59 63.725 3.823 ;
      RECT 63.535 3.661 63.745 3.82 ;
      RECT 63.53 3.692 63.745 3.818 ;
      RECT 63.535 3.689 63.76 3.808 ;
      RECT 63.53 3.735 63.775 3.793 ;
      RECT 63.53 3.763 63.78 3.778 ;
      RECT 63.54 3.565 63.71 3.828 ;
      RECT 63.3 2.575 63.47 2.745 ;
      RECT 63.265 2.575 63.47 2.74 ;
      RECT 63.255 2.575 63.47 2.733 ;
      RECT 63.25 2.56 63.42 2.73 ;
      RECT 62.08 3.097 62.345 3.54 ;
      RECT 62.075 3.068 62.29 3.538 ;
      RECT 62.07 3.222 62.35 3.533 ;
      RECT 62.075 3.117 62.35 3.533 ;
      RECT 62.075 3.128 62.36 3.52 ;
      RECT 62.075 3.075 62.32 3.538 ;
      RECT 62.08 3.062 62.29 3.54 ;
      RECT 62.08 3.06 62.24 3.54 ;
      RECT 62.181 3.052 62.24 3.54 ;
      RECT 62.095 3.053 62.24 3.54 ;
      RECT 62.181 3.051 62.23 3.54 ;
      RECT 61.985 1.866 62.16 2.165 ;
      RECT 62.035 1.828 62.16 2.165 ;
      RECT 62.02 1.83 62.246 2.157 ;
      RECT 62.02 1.833 62.285 2.144 ;
      RECT 62.02 1.834 62.295 2.13 ;
      RECT 61.975 1.885 62.295 2.12 ;
      RECT 62.02 1.835 62.3 2.115 ;
      RECT 61.975 2.045 62.305 2.105 ;
      RECT 61.96 1.905 62.3 2.045 ;
      RECT 61.955 1.921 62.3 1.985 ;
      RECT 62 1.845 62.3 2.115 ;
      RECT 62.035 1.826 62.121 2.165 ;
      RECT 60.13 1.74 60.3 2.935 ;
      RECT 60.13 1.74 60.595 1.91 ;
      RECT 60.13 6.97 60.595 7.14 ;
      RECT 60.13 5.945 60.3 7.14 ;
      RECT 59.14 1.74 59.31 2.935 ;
      RECT 59.14 1.74 59.605 1.91 ;
      RECT 59.14 6.97 59.605 7.14 ;
      RECT 59.14 5.945 59.31 7.14 ;
      RECT 57.285 2.635 57.455 3.865 ;
      RECT 57.34 0.855 57.51 2.805 ;
      RECT 57.285 0.575 57.455 1.025 ;
      RECT 57.285 7.855 57.455 8.305 ;
      RECT 57.34 6.075 57.51 8.025 ;
      RECT 57.285 5.015 57.455 6.245 ;
      RECT 56.765 0.575 56.935 3.865 ;
      RECT 56.765 2.075 57.17 2.405 ;
      RECT 56.765 1.235 57.17 1.565 ;
      RECT 56.765 5.015 56.935 8.305 ;
      RECT 56.765 7.315 57.17 7.645 ;
      RECT 56.765 6.475 57.17 6.805 ;
      RECT 54.69 3.126 54.695 3.298 ;
      RECT 54.685 3.119 54.69 3.388 ;
      RECT 54.68 3.113 54.685 3.407 ;
      RECT 54.66 3.107 54.68 3.417 ;
      RECT 54.645 3.102 54.66 3.425 ;
      RECT 54.608 3.096 54.645 3.423 ;
      RECT 54.522 3.082 54.608 3.419 ;
      RECT 54.436 3.064 54.522 3.414 ;
      RECT 54.35 3.045 54.436 3.408 ;
      RECT 54.32 3.033 54.35 3.404 ;
      RECT 54.3 3.027 54.32 3.403 ;
      RECT 54.235 3.025 54.3 3.401 ;
      RECT 54.22 3.025 54.235 3.393 ;
      RECT 54.205 3.025 54.22 3.38 ;
      RECT 54.2 3.025 54.205 3.37 ;
      RECT 54.185 3.025 54.2 3.348 ;
      RECT 54.17 3.025 54.185 3.315 ;
      RECT 54.165 3.025 54.17 3.293 ;
      RECT 54.155 3.025 54.165 3.275 ;
      RECT 54.14 3.025 54.155 3.253 ;
      RECT 54.12 3.025 54.14 3.215 ;
      RECT 54.47 2.31 54.505 2.749 ;
      RECT 54.47 2.31 54.51 2.748 ;
      RECT 54.415 2.37 54.51 2.747 ;
      RECT 54.28 2.542 54.51 2.746 ;
      RECT 54.39 2.42 54.51 2.746 ;
      RECT 54.28 2.542 54.535 2.736 ;
      RECT 54.335 2.487 54.615 2.653 ;
      RECT 54.51 2.281 54.515 2.744 ;
      RECT 54.365 2.457 54.655 2.53 ;
      RECT 54.38 2.44 54.51 2.746 ;
      RECT 54.515 2.28 54.685 2.468 ;
      RECT 54.505 2.283 54.685 2.468 ;
      RECT 54.01 2.16 54.18 2.47 ;
      RECT 54.01 2.16 54.185 2.443 ;
      RECT 54.01 2.16 54.19 2.42 ;
      RECT 54.01 2.16 54.2 2.37 ;
      RECT 54.005 2.265 54.2 2.34 ;
      RECT 54.04 1.835 54.21 2.313 ;
      RECT 54.04 1.835 54.225 2.234 ;
      RECT 54.03 2.045 54.225 2.234 ;
      RECT 54.04 1.845 54.235 2.149 ;
      RECT 53.97 2.587 53.975 2.79 ;
      RECT 53.96 2.575 53.97 2.9 ;
      RECT 53.935 2.575 53.96 2.94 ;
      RECT 53.855 2.575 53.935 3.025 ;
      RECT 53.845 2.575 53.855 3.095 ;
      RECT 53.82 2.575 53.845 3.118 ;
      RECT 53.8 2.575 53.82 3.153 ;
      RECT 53.755 2.585 53.8 3.196 ;
      RECT 53.745 2.597 53.755 3.233 ;
      RECT 53.725 2.611 53.745 3.253 ;
      RECT 53.715 2.629 53.725 3.269 ;
      RECT 53.7 2.655 53.715 3.279 ;
      RECT 53.685 2.696 53.7 3.293 ;
      RECT 53.675 2.731 53.685 3.303 ;
      RECT 53.67 2.747 53.675 3.308 ;
      RECT 53.66 2.762 53.67 3.313 ;
      RECT 53.64 2.805 53.66 3.323 ;
      RECT 53.62 2.842 53.64 3.336 ;
      RECT 53.585 2.865 53.62 3.354 ;
      RECT 53.575 2.879 53.585 3.37 ;
      RECT 53.555 2.889 53.575 3.38 ;
      RECT 53.55 2.898 53.555 3.388 ;
      RECT 53.54 2.905 53.55 3.395 ;
      RECT 53.53 2.912 53.54 3.403 ;
      RECT 53.515 2.922 53.53 3.411 ;
      RECT 53.505 2.936 53.515 3.421 ;
      RECT 53.495 2.948 53.505 3.433 ;
      RECT 53.48 2.97 53.495 3.446 ;
      RECT 53.47 2.992 53.48 3.457 ;
      RECT 53.46 3.012 53.47 3.466 ;
      RECT 53.455 3.027 53.46 3.473 ;
      RECT 53.425 3.06 53.455 3.487 ;
      RECT 53.415 3.095 53.425 3.502 ;
      RECT 53.41 3.102 53.415 3.508 ;
      RECT 53.39 3.117 53.41 3.515 ;
      RECT 53.385 3.132 53.39 3.523 ;
      RECT 53.38 3.141 53.385 3.528 ;
      RECT 53.365 3.147 53.38 3.535 ;
      RECT 53.36 3.153 53.365 3.543 ;
      RECT 53.355 3.157 53.36 3.55 ;
      RECT 53.35 3.161 53.355 3.56 ;
      RECT 53.34 3.166 53.35 3.57 ;
      RECT 53.32 3.177 53.34 3.598 ;
      RECT 53.305 3.189 53.32 3.625 ;
      RECT 53.285 3.202 53.305 3.65 ;
      RECT 53.265 3.217 53.285 3.674 ;
      RECT 53.25 3.232 53.265 3.689 ;
      RECT 53.245 3.243 53.25 3.698 ;
      RECT 53.18 3.288 53.245 3.708 ;
      RECT 53.145 3.347 53.18 3.721 ;
      RECT 53.14 3.37 53.145 3.727 ;
      RECT 53.135 3.377 53.14 3.729 ;
      RECT 53.12 3.387 53.135 3.732 ;
      RECT 53.09 3.412 53.12 3.736 ;
      RECT 53.085 3.43 53.09 3.74 ;
      RECT 53.08 3.437 53.085 3.741 ;
      RECT 53.06 3.445 53.08 3.745 ;
      RECT 53.05 3.452 53.06 3.749 ;
      RECT 53.006 3.463 53.05 3.756 ;
      RECT 52.92 3.491 53.006 3.772 ;
      RECT 52.86 3.515 52.92 3.79 ;
      RECT 52.815 3.525 52.86 3.804 ;
      RECT 52.756 3.533 52.815 3.818 ;
      RECT 52.67 3.54 52.756 3.837 ;
      RECT 52.645 3.545 52.67 3.852 ;
      RECT 52.565 3.548 52.645 3.855 ;
      RECT 52.485 3.552 52.565 3.842 ;
      RECT 52.476 3.555 52.485 3.827 ;
      RECT 52.39 3.555 52.476 3.812 ;
      RECT 52.33 3.557 52.39 3.789 ;
      RECT 52.326 3.56 52.33 3.779 ;
      RECT 52.24 3.56 52.326 3.764 ;
      RECT 52.165 3.56 52.24 3.74 ;
      RECT 53.48 2.569 53.49 2.745 ;
      RECT 53.435 2.536 53.48 2.745 ;
      RECT 53.39 2.487 53.435 2.745 ;
      RECT 53.36 2.457 53.39 2.746 ;
      RECT 53.355 2.44 53.36 2.747 ;
      RECT 53.33 2.42 53.355 2.748 ;
      RECT 53.315 2.395 53.33 2.749 ;
      RECT 53.31 2.382 53.315 2.75 ;
      RECT 53.305 2.376 53.31 2.748 ;
      RECT 53.3 2.368 53.305 2.742 ;
      RECT 53.275 2.36 53.3 2.722 ;
      RECT 53.255 2.349 53.275 2.693 ;
      RECT 53.225 2.334 53.255 2.664 ;
      RECT 53.205 2.32 53.225 2.636 ;
      RECT 53.195 2.314 53.205 2.615 ;
      RECT 53.19 2.311 53.195 2.598 ;
      RECT 53.185 2.308 53.19 2.583 ;
      RECT 53.17 2.303 53.185 2.548 ;
      RECT 53.165 2.299 53.17 2.515 ;
      RECT 53.145 2.294 53.165 2.491 ;
      RECT 53.115 2.286 53.145 2.456 ;
      RECT 53.1 2.28 53.115 2.433 ;
      RECT 53.06 2.273 53.1 2.418 ;
      RECT 53.035 2.265 53.06 2.398 ;
      RECT 53.015 2.26 53.035 2.388 ;
      RECT 52.98 2.254 53.015 2.383 ;
      RECT 52.935 2.245 52.98 2.382 ;
      RECT 52.905 2.241 52.935 2.384 ;
      RECT 52.82 2.249 52.905 2.388 ;
      RECT 52.75 2.26 52.82 2.41 ;
      RECT 52.737 2.266 52.75 2.433 ;
      RECT 52.651 2.273 52.737 2.455 ;
      RECT 52.565 2.285 52.651 2.492 ;
      RECT 52.565 2.662 52.575 2.9 ;
      RECT 52.56 2.291 52.565 2.515 ;
      RECT 52.555 2.547 52.565 2.9 ;
      RECT 52.555 2.292 52.56 2.52 ;
      RECT 52.55 2.293 52.555 2.9 ;
      RECT 52.526 2.295 52.55 2.901 ;
      RECT 52.44 2.303 52.526 2.903 ;
      RECT 52.42 2.317 52.44 2.906 ;
      RECT 52.415 2.345 52.42 2.907 ;
      RECT 52.41 2.357 52.415 2.908 ;
      RECT 52.405 2.372 52.41 2.909 ;
      RECT 52.395 2.402 52.405 2.91 ;
      RECT 52.39 2.44 52.395 2.908 ;
      RECT 52.385 2.46 52.39 2.903 ;
      RECT 52.37 2.495 52.385 2.888 ;
      RECT 52.36 2.547 52.37 2.868 ;
      RECT 52.355 2.577 52.36 2.856 ;
      RECT 52.34 2.59 52.355 2.839 ;
      RECT 52.315 2.594 52.34 2.806 ;
      RECT 52.3 2.592 52.315 2.783 ;
      RECT 52.285 2.591 52.3 2.78 ;
      RECT 52.225 2.589 52.285 2.778 ;
      RECT 52.215 2.587 52.225 2.773 ;
      RECT 52.175 2.586 52.215 2.77 ;
      RECT 52.105 2.583 52.175 2.768 ;
      RECT 52.05 2.581 52.105 2.763 ;
      RECT 51.98 2.575 52.05 2.758 ;
      RECT 51.971 2.575 51.98 2.755 ;
      RECT 51.885 2.575 51.971 2.75 ;
      RECT 51.88 2.575 51.885 2.745 ;
      RECT 53.185 1.81 53.36 2.16 ;
      RECT 53.185 1.825 53.37 2.158 ;
      RECT 53.16 1.775 53.305 2.155 ;
      RECT 53.14 1.776 53.305 2.148 ;
      RECT 53.13 1.777 53.315 2.143 ;
      RECT 53.1 1.778 53.315 2.13 ;
      RECT 53.05 1.779 53.315 2.106 ;
      RECT 53.045 1.781 53.315 2.091 ;
      RECT 53.045 1.847 53.375 2.085 ;
      RECT 53.025 1.788 53.33 2.065 ;
      RECT 53.015 1.797 53.34 1.92 ;
      RECT 53.025 1.792 53.34 2.065 ;
      RECT 53.045 1.782 53.33 2.091 ;
      RECT 52.63 3.107 52.8 3.395 ;
      RECT 52.625 3.125 52.81 3.39 ;
      RECT 52.59 3.133 52.875 3.31 ;
      RECT 52.59 3.133 52.961 3.3 ;
      RECT 52.59 3.133 53.015 3.246 ;
      RECT 52.875 3.03 53.045 3.214 ;
      RECT 52.59 3.185 53.05 3.202 ;
      RECT 52.575 3.155 53.045 3.198 ;
      RECT 52.835 3.037 52.875 3.349 ;
      RECT 52.715 3.074 53.045 3.214 ;
      RECT 52.81 3.049 52.835 3.375 ;
      RECT 52.8 3.056 53.045 3.214 ;
      RECT 52.931 2.52 53 2.779 ;
      RECT 52.931 2.575 53.005 2.778 ;
      RECT 52.845 2.575 53.005 2.777 ;
      RECT 52.84 2.575 53.01 2.77 ;
      RECT 52.83 2.52 53 2.765 ;
      RECT 52.21 1.819 52.385 2.12 ;
      RECT 52.195 1.807 52.21 2.105 ;
      RECT 52.165 1.806 52.195 2.058 ;
      RECT 52.165 1.824 52.39 2.053 ;
      RECT 52.15 1.808 52.21 2.018 ;
      RECT 52.145 1.83 52.4 1.918 ;
      RECT 52.145 1.813 52.296 1.918 ;
      RECT 52.145 1.815 52.3 1.918 ;
      RECT 52.15 1.811 52.296 2.018 ;
      RECT 52.255 3.047 52.26 3.395 ;
      RECT 52.245 3.037 52.255 3.401 ;
      RECT 52.21 3.027 52.245 3.403 ;
      RECT 52.172 3.022 52.21 3.407 ;
      RECT 52.086 3.015 52.172 3.414 ;
      RECT 52 3.005 52.086 3.424 ;
      RECT 51.955 3 52 3.432 ;
      RECT 51.951 3 51.955 3.436 ;
      RECT 51.865 3 51.951 3.443 ;
      RECT 51.85 3 51.865 3.443 ;
      RECT 51.84 2.998 51.85 3.415 ;
      RECT 51.83 2.994 51.84 3.358 ;
      RECT 51.81 2.988 51.83 3.29 ;
      RECT 51.805 2.984 51.81 3.238 ;
      RECT 51.795 2.983 51.805 3.205 ;
      RECT 51.745 2.981 51.795 3.19 ;
      RECT 51.72 2.979 51.745 3.185 ;
      RECT 51.677 2.977 51.72 3.181 ;
      RECT 51.591 2.973 51.677 3.169 ;
      RECT 51.505 2.968 51.591 3.153 ;
      RECT 51.475 2.965 51.505 3.14 ;
      RECT 51.45 2.964 51.475 3.128 ;
      RECT 51.445 2.964 51.45 3.118 ;
      RECT 51.405 2.963 51.445 3.11 ;
      RECT 51.39 2.962 51.405 3.103 ;
      RECT 51.34 2.961 51.39 3.095 ;
      RECT 51.338 2.96 51.34 3.09 ;
      RECT 51.252 2.958 51.338 3.09 ;
      RECT 51.166 2.953 51.252 3.09 ;
      RECT 51.08 2.949 51.166 3.09 ;
      RECT 51.031 2.945 51.08 3.088 ;
      RECT 50.945 2.942 51.031 3.083 ;
      RECT 50.922 2.939 50.945 3.079 ;
      RECT 50.836 2.936 50.922 3.074 ;
      RECT 50.75 2.932 50.836 3.065 ;
      RECT 50.725 2.925 50.75 3.06 ;
      RECT 50.665 2.89 50.725 3.057 ;
      RECT 50.645 2.815 50.665 3.054 ;
      RECT 50.64 2.757 50.645 3.053 ;
      RECT 50.615 2.697 50.64 3.052 ;
      RECT 50.54 2.575 50.615 3.048 ;
      RECT 50.53 2.575 50.54 3.04 ;
      RECT 50.515 2.575 50.53 3.03 ;
      RECT 50.5 2.575 50.515 3 ;
      RECT 50.485 2.575 50.5 2.945 ;
      RECT 50.47 2.575 50.485 2.883 ;
      RECT 50.445 2.575 50.47 2.808 ;
      RECT 50.44 2.575 50.445 2.758 ;
      RECT 51.785 2.12 51.805 2.429 ;
      RECT 51.771 2.122 51.82 2.426 ;
      RECT 51.771 2.127 51.84 2.417 ;
      RECT 51.685 2.125 51.82 2.411 ;
      RECT 51.685 2.133 51.875 2.394 ;
      RECT 51.65 2.135 51.875 2.393 ;
      RECT 51.62 2.143 51.875 2.384 ;
      RECT 51.61 2.148 51.895 2.37 ;
      RECT 51.65 2.138 51.895 2.37 ;
      RECT 51.65 2.141 51.905 2.358 ;
      RECT 51.62 2.143 51.915 2.345 ;
      RECT 51.62 2.147 51.925 2.288 ;
      RECT 51.61 2.152 51.93 2.203 ;
      RECT 51.771 2.12 51.805 2.426 ;
      RECT 51.21 2.223 51.215 2.435 ;
      RECT 51.085 2.22 51.1 2.435 ;
      RECT 50.55 2.25 50.62 2.435 ;
      RECT 50.435 2.25 50.47 2.43 ;
      RECT 51.556 2.552 51.575 2.746 ;
      RECT 51.47 2.507 51.556 2.747 ;
      RECT 51.46 2.46 51.47 2.749 ;
      RECT 51.455 2.44 51.46 2.75 ;
      RECT 51.435 2.405 51.455 2.751 ;
      RECT 51.42 2.355 51.435 2.752 ;
      RECT 51.4 2.292 51.42 2.753 ;
      RECT 51.39 2.255 51.4 2.754 ;
      RECT 51.375 2.244 51.39 2.755 ;
      RECT 51.37 2.236 51.375 2.753 ;
      RECT 51.36 2.235 51.37 2.745 ;
      RECT 51.33 2.232 51.36 2.724 ;
      RECT 51.255 2.227 51.33 2.669 ;
      RECT 51.24 2.223 51.255 2.615 ;
      RECT 51.23 2.223 51.24 2.51 ;
      RECT 51.215 2.223 51.23 2.443 ;
      RECT 51.2 2.223 51.21 2.433 ;
      RECT 51.145 2.222 51.2 2.43 ;
      RECT 51.1 2.22 51.145 2.433 ;
      RECT 51.072 2.22 51.085 2.436 ;
      RECT 50.986 2.224 51.072 2.438 ;
      RECT 50.9 2.23 50.986 2.443 ;
      RECT 50.88 2.234 50.9 2.445 ;
      RECT 50.878 2.235 50.88 2.444 ;
      RECT 50.792 2.237 50.878 2.443 ;
      RECT 50.706 2.242 50.792 2.44 ;
      RECT 50.62 2.247 50.706 2.437 ;
      RECT 50.47 2.25 50.55 2.433 ;
      RECT 51.246 3.225 51.295 3.559 ;
      RECT 51.246 3.225 51.3 3.558 ;
      RECT 51.16 3.225 51.3 3.557 ;
      RECT 50.935 3.333 51.305 3.555 ;
      RECT 51.16 3.225 51.33 3.548 ;
      RECT 51.13 3.237 51.335 3.539 ;
      RECT 51.115 3.255 51.34 3.536 ;
      RECT 50.93 3.339 51.34 3.463 ;
      RECT 50.925 3.346 51.34 3.423 ;
      RECT 50.94 3.312 51.34 3.536 ;
      RECT 51.101 3.258 51.305 3.555 ;
      RECT 51.015 3.278 51.34 3.536 ;
      RECT 51.115 3.252 51.335 3.539 ;
      RECT 50.885 2.576 51.075 2.77 ;
      RECT 50.88 2.578 51.075 2.769 ;
      RECT 50.875 2.582 51.09 2.766 ;
      RECT 50.89 2.575 51.09 2.766 ;
      RECT 50.875 2.685 51.095 2.761 ;
      RECT 50.17 3.185 50.261 3.483 ;
      RECT 50.165 3.187 50.34 3.478 ;
      RECT 50.17 3.185 50.34 3.478 ;
      RECT 50.165 3.191 50.36 3.476 ;
      RECT 50.165 3.246 50.4 3.475 ;
      RECT 50.165 3.281 50.415 3.469 ;
      RECT 50.165 3.315 50.425 3.459 ;
      RECT 50.155 3.195 50.36 3.31 ;
      RECT 50.155 3.215 50.375 3.31 ;
      RECT 50.155 3.198 50.365 3.31 ;
      RECT 50.38 1.966 50.385 2.028 ;
      RECT 50.375 1.888 50.38 2.051 ;
      RECT 50.37 1.845 50.375 2.062 ;
      RECT 50.365 1.835 50.37 2.074 ;
      RECT 50.36 1.835 50.365 2.083 ;
      RECT 50.335 1.835 50.36 2.115 ;
      RECT 50.33 1.835 50.335 2.148 ;
      RECT 50.315 1.835 50.33 2.173 ;
      RECT 50.305 1.835 50.315 2.2 ;
      RECT 50.3 1.835 50.305 2.213 ;
      RECT 50.295 1.835 50.3 2.228 ;
      RECT 50.285 1.835 50.295 2.243 ;
      RECT 50.28 1.835 50.285 2.263 ;
      RECT 50.255 1.835 50.28 2.298 ;
      RECT 50.21 1.835 50.255 2.343 ;
      RECT 50.2 1.835 50.21 2.356 ;
      RECT 50.115 1.92 50.2 2.363 ;
      RECT 50.08 2.042 50.115 2.372 ;
      RECT 50.075 2.082 50.08 2.376 ;
      RECT 50.055 2.105 50.075 2.378 ;
      RECT 50.05 2.135 50.055 2.381 ;
      RECT 50.04 2.147 50.05 2.382 ;
      RECT 49.995 2.17 50.04 2.387 ;
      RECT 49.955 2.2 49.995 2.395 ;
      RECT 49.92 2.212 49.955 2.401 ;
      RECT 49.915 2.217 49.92 2.405 ;
      RECT 49.845 2.227 49.915 2.412 ;
      RECT 49.805 2.237 49.845 2.422 ;
      RECT 49.785 2.242 49.805 2.428 ;
      RECT 49.775 2.246 49.785 2.433 ;
      RECT 49.77 2.249 49.775 2.436 ;
      RECT 49.76 2.25 49.77 2.437 ;
      RECT 49.735 2.252 49.76 2.441 ;
      RECT 49.725 2.257 49.735 2.444 ;
      RECT 49.68 2.265 49.725 2.445 ;
      RECT 49.555 2.27 49.68 2.445 ;
      RECT 50.11 2.567 50.13 2.749 ;
      RECT 50.061 2.552 50.11 2.748 ;
      RECT 49.975 2.567 50.13 2.746 ;
      RECT 49.96 2.567 50.13 2.745 ;
      RECT 49.925 2.545 50.095 2.73 ;
      RECT 49.995 3.565 50.01 3.774 ;
      RECT 49.995 3.573 50.015 3.773 ;
      RECT 49.94 3.573 50.015 3.772 ;
      RECT 49.92 3.577 50.02 3.77 ;
      RECT 49.9 3.527 49.94 3.769 ;
      RECT 49.845 3.585 50.025 3.767 ;
      RECT 49.81 3.542 49.94 3.765 ;
      RECT 49.806 3.545 49.995 3.764 ;
      RECT 49.72 3.553 49.995 3.762 ;
      RECT 49.72 3.597 50.03 3.755 ;
      RECT 49.71 3.69 50.03 3.753 ;
      RECT 49.72 3.609 50.035 3.738 ;
      RECT 49.72 3.63 50.05 3.708 ;
      RECT 49.72 3.657 50.055 3.678 ;
      RECT 49.845 3.535 49.94 3.767 ;
      RECT 49.475 2.58 49.48 3.118 ;
      RECT 49.28 2.91 49.285 3.105 ;
      RECT 47.58 2.575 47.595 2.955 ;
      RECT 49.645 2.575 49.65 2.745 ;
      RECT 49.64 2.575 49.645 2.755 ;
      RECT 49.635 2.575 49.64 2.768 ;
      RECT 49.61 2.575 49.635 2.81 ;
      RECT 49.585 2.575 49.61 2.883 ;
      RECT 49.57 2.575 49.585 2.935 ;
      RECT 49.565 2.575 49.57 2.965 ;
      RECT 49.54 2.575 49.565 3.005 ;
      RECT 49.525 2.575 49.54 3.06 ;
      RECT 49.52 2.575 49.525 3.093 ;
      RECT 49.495 2.575 49.52 3.113 ;
      RECT 49.48 2.575 49.495 3.119 ;
      RECT 49.41 2.61 49.475 3.115 ;
      RECT 49.36 2.665 49.41 3.11 ;
      RECT 49.35 2.697 49.36 3.108 ;
      RECT 49.345 2.722 49.35 3.108 ;
      RECT 49.325 2.795 49.345 3.108 ;
      RECT 49.315 2.875 49.325 3.107 ;
      RECT 49.3 2.905 49.315 3.107 ;
      RECT 49.285 2.91 49.3 3.106 ;
      RECT 49.225 2.912 49.28 3.103 ;
      RECT 49.195 2.917 49.225 3.099 ;
      RECT 49.193 2.92 49.195 3.098 ;
      RECT 49.107 2.922 49.193 3.095 ;
      RECT 49.021 2.928 49.107 3.089 ;
      RECT 48.935 2.933 49.021 3.083 ;
      RECT 48.862 2.938 48.935 3.084 ;
      RECT 48.776 2.944 48.862 3.092 ;
      RECT 48.69 2.95 48.776 3.101 ;
      RECT 48.67 2.954 48.69 3.106 ;
      RECT 48.623 2.956 48.67 3.109 ;
      RECT 48.537 2.961 48.623 3.115 ;
      RECT 48.451 2.966 48.537 3.124 ;
      RECT 48.365 2.972 48.451 3.132 ;
      RECT 48.28 2.97 48.365 3.141 ;
      RECT 48.276 2.965 48.28 3.145 ;
      RECT 48.19 2.96 48.276 3.137 ;
      RECT 48.126 2.951 48.19 3.125 ;
      RECT 48.04 2.942 48.126 3.112 ;
      RECT 48.016 2.935 48.04 3.103 ;
      RECT 47.93 2.929 48.016 3.09 ;
      RECT 47.89 2.922 47.93 3.076 ;
      RECT 47.885 2.912 47.89 3.072 ;
      RECT 47.875 2.9 47.885 3.071 ;
      RECT 47.855 2.87 47.875 3.068 ;
      RECT 47.8 2.79 47.855 3.062 ;
      RECT 47.78 2.709 47.8 3.057 ;
      RECT 47.76 2.667 47.78 3.053 ;
      RECT 47.735 2.62 47.76 3.047 ;
      RECT 47.73 2.595 47.735 3.044 ;
      RECT 47.695 2.575 47.73 3.039 ;
      RECT 47.686 2.575 47.695 3.032 ;
      RECT 47.6 2.575 47.686 3.002 ;
      RECT 47.595 2.575 47.6 2.965 ;
      RECT 47.56 2.575 47.58 2.887 ;
      RECT 47.555 2.617 47.56 2.852 ;
      RECT 47.55 2.692 47.555 2.808 ;
      RECT 49 2.497 49.175 2.745 ;
      RECT 49 2.497 49.18 2.743 ;
      RECT 48.995 2.529 49.18 2.703 ;
      RECT 49.025 2.47 49.195 2.69 ;
      RECT 48.99 2.547 49.195 2.623 ;
      RECT 48.3 2.01 48.47 2.185 ;
      RECT 48.3 2.01 48.642 2.177 ;
      RECT 48.3 2.01 48.725 2.171 ;
      RECT 48.3 2.01 48.76 2.167 ;
      RECT 48.3 2.01 48.78 2.166 ;
      RECT 48.3 2.01 48.866 2.162 ;
      RECT 48.76 1.835 48.93 2.157 ;
      RECT 48.335 1.942 48.96 2.155 ;
      RECT 48.325 1.997 48.965 2.153 ;
      RECT 48.3 2.033 48.975 2.148 ;
      RECT 48.3 2.06 48.98 2.078 ;
      RECT 48.365 1.885 48.94 2.155 ;
      RECT 48.556 1.87 48.94 2.155 ;
      RECT 48.39 1.873 48.94 2.155 ;
      RECT 48.47 1.871 48.556 2.182 ;
      RECT 48.556 1.868 48.935 2.155 ;
      RECT 48.74 1.845 48.935 2.155 ;
      RECT 48.642 1.866 48.935 2.155 ;
      RECT 48.725 1.86 48.74 2.168 ;
      RECT 48.875 3.225 48.88 3.425 ;
      RECT 48.34 3.29 48.385 3.425 ;
      RECT 48.91 3.225 48.93 3.398 ;
      RECT 48.88 3.225 48.91 3.413 ;
      RECT 48.815 3.225 48.875 3.45 ;
      RECT 48.8 3.225 48.815 3.48 ;
      RECT 48.785 3.225 48.8 3.493 ;
      RECT 48.765 3.225 48.785 3.508 ;
      RECT 48.76 3.225 48.765 3.517 ;
      RECT 48.75 3.229 48.76 3.522 ;
      RECT 48.735 3.239 48.75 3.533 ;
      RECT 48.71 3.255 48.735 3.543 ;
      RECT 48.7 3.269 48.71 3.545 ;
      RECT 48.68 3.281 48.7 3.542 ;
      RECT 48.65 3.302 48.68 3.536 ;
      RECT 48.64 3.314 48.65 3.531 ;
      RECT 48.63 3.312 48.64 3.528 ;
      RECT 48.615 3.311 48.63 3.523 ;
      RECT 48.61 3.31 48.615 3.518 ;
      RECT 48.575 3.308 48.61 3.508 ;
      RECT 48.555 3.305 48.575 3.49 ;
      RECT 48.545 3.303 48.555 3.485 ;
      RECT 48.535 3.302 48.545 3.48 ;
      RECT 48.5 3.3 48.535 3.468 ;
      RECT 48.445 3.296 48.5 3.448 ;
      RECT 48.435 3.294 48.445 3.433 ;
      RECT 48.43 3.294 48.435 3.428 ;
      RECT 48.385 3.292 48.43 3.425 ;
      RECT 48.29 3.29 48.34 3.429 ;
      RECT 48.28 3.291 48.29 3.434 ;
      RECT 48.22 3.298 48.28 3.448 ;
      RECT 48.195 3.306 48.22 3.468 ;
      RECT 48.185 3.31 48.195 3.48 ;
      RECT 48.18 3.311 48.185 3.485 ;
      RECT 48.165 3.313 48.18 3.488 ;
      RECT 48.15 3.315 48.165 3.493 ;
      RECT 48.145 3.315 48.15 3.496 ;
      RECT 48.1 3.32 48.145 3.507 ;
      RECT 48.095 3.324 48.1 3.519 ;
      RECT 48.07 3.32 48.095 3.523 ;
      RECT 48.06 3.316 48.07 3.527 ;
      RECT 48.05 3.315 48.06 3.531 ;
      RECT 48.035 3.305 48.05 3.537 ;
      RECT 48.03 3.293 48.035 3.541 ;
      RECT 48.025 3.29 48.03 3.542 ;
      RECT 48.02 3.287 48.025 3.544 ;
      RECT 48.005 3.275 48.02 3.543 ;
      RECT 47.99 3.257 48.005 3.54 ;
      RECT 47.97 3.236 47.99 3.533 ;
      RECT 47.905 3.225 47.97 3.505 ;
      RECT 47.901 3.225 47.905 3.484 ;
      RECT 47.815 3.225 47.901 3.454 ;
      RECT 47.8 3.225 47.815 3.41 ;
      RECT 48.375 2.325 48.38 2.56 ;
      RECT 47.505 2.241 47.51 2.445 ;
      RECT 48.085 2.27 48.09 2.425 ;
      RECT 48.005 2.25 48.01 2.425 ;
      RECT 48.675 2.392 48.69 2.745 ;
      RECT 48.601 2.377 48.675 2.745 ;
      RECT 48.515 2.36 48.601 2.745 ;
      RECT 48.505 2.35 48.515 2.743 ;
      RECT 48.5 2.348 48.505 2.738 ;
      RECT 48.485 2.346 48.5 2.724 ;
      RECT 48.415 2.338 48.485 2.664 ;
      RECT 48.395 2.329 48.415 2.598 ;
      RECT 48.39 2.326 48.395 2.578 ;
      RECT 48.38 2.325 48.39 2.568 ;
      RECT 48.37 2.325 48.375 2.552 ;
      RECT 48.36 2.324 48.37 2.542 ;
      RECT 48.35 2.322 48.36 2.53 ;
      RECT 48.335 2.319 48.35 2.51 ;
      RECT 48.325 2.317 48.335 2.495 ;
      RECT 48.305 2.314 48.325 2.483 ;
      RECT 48.3 2.312 48.305 2.473 ;
      RECT 48.275 2.31 48.3 2.46 ;
      RECT 48.245 2.305 48.275 2.445 ;
      RECT 48.165 2.296 48.245 2.436 ;
      RECT 48.12 2.285 48.165 2.429 ;
      RECT 48.1 2.276 48.12 2.426 ;
      RECT 48.09 2.271 48.1 2.425 ;
      RECT 48.045 2.265 48.085 2.425 ;
      RECT 48.03 2.257 48.045 2.425 ;
      RECT 48.01 2.252 48.03 2.425 ;
      RECT 47.99 2.249 48.005 2.425 ;
      RECT 47.907 2.248 47.99 2.424 ;
      RECT 47.821 2.247 47.907 2.42 ;
      RECT 47.735 2.245 47.821 2.417 ;
      RECT 47.682 2.244 47.735 2.419 ;
      RECT 47.596 2.243 47.682 2.428 ;
      RECT 47.51 2.242 47.596 2.44 ;
      RECT 47.49 2.241 47.505 2.448 ;
      RECT 47.41 2.24 47.49 2.46 ;
      RECT 47.385 2.24 47.41 2.473 ;
      RECT 47.36 2.24 47.385 2.488 ;
      RECT 47.355 2.24 47.36 2.51 ;
      RECT 47.35 2.24 47.355 2.528 ;
      RECT 47.345 2.24 47.35 2.545 ;
      RECT 47.34 2.24 47.345 2.558 ;
      RECT 47.335 2.24 47.34 2.568 ;
      RECT 47.295 2.24 47.335 2.653 ;
      RECT 47.28 2.24 47.295 2.738 ;
      RECT 47.27 2.241 47.28 2.75 ;
      RECT 47.235 2.246 47.27 2.755 ;
      RECT 47.195 2.255 47.235 2.755 ;
      RECT 47.18 2.265 47.195 2.755 ;
      RECT 47.175 2.275 47.18 2.755 ;
      RECT 47.155 2.302 47.175 2.755 ;
      RECT 47.105 2.385 47.155 2.755 ;
      RECT 47.1 2.447 47.105 2.755 ;
      RECT 47.09 2.46 47.1 2.755 ;
      RECT 47.08 2.482 47.09 2.755 ;
      RECT 47.07 2.507 47.08 2.75 ;
      RECT 47.065 2.545 47.07 2.743 ;
      RECT 47.055 2.655 47.065 2.738 ;
      RECT 48.45 3.576 48.465 3.835 ;
      RECT 48.45 3.591 48.47 3.834 ;
      RECT 48.366 3.591 48.47 3.832 ;
      RECT 48.366 3.605 48.475 3.831 ;
      RECT 48.28 3.647 48.48 3.828 ;
      RECT 48.275 3.59 48.465 3.823 ;
      RECT 48.275 3.661 48.485 3.82 ;
      RECT 48.27 3.692 48.485 3.818 ;
      RECT 48.275 3.689 48.5 3.808 ;
      RECT 48.27 3.735 48.515 3.793 ;
      RECT 48.27 3.763 48.52 3.778 ;
      RECT 48.28 3.565 48.45 3.828 ;
      RECT 48.04 2.575 48.21 2.745 ;
      RECT 48.005 2.575 48.21 2.74 ;
      RECT 47.995 2.575 48.21 2.733 ;
      RECT 47.99 2.56 48.16 2.73 ;
      RECT 46.82 3.097 47.085 3.54 ;
      RECT 46.815 3.068 47.03 3.538 ;
      RECT 46.81 3.222 47.09 3.533 ;
      RECT 46.815 3.117 47.09 3.533 ;
      RECT 46.815 3.128 47.1 3.52 ;
      RECT 46.815 3.075 47.06 3.538 ;
      RECT 46.82 3.062 47.03 3.54 ;
      RECT 46.82 3.06 46.98 3.54 ;
      RECT 46.921 3.052 46.98 3.54 ;
      RECT 46.835 3.053 46.98 3.54 ;
      RECT 46.921 3.051 46.97 3.54 ;
      RECT 46.725 1.866 46.9 2.165 ;
      RECT 46.775 1.828 46.9 2.165 ;
      RECT 46.76 1.83 46.986 2.157 ;
      RECT 46.76 1.833 47.025 2.144 ;
      RECT 46.76 1.834 47.035 2.13 ;
      RECT 46.715 1.885 47.035 2.12 ;
      RECT 46.76 1.835 47.04 2.115 ;
      RECT 46.715 2.045 47.045 2.105 ;
      RECT 46.7 1.905 47.04 2.045 ;
      RECT 46.695 1.921 47.04 1.985 ;
      RECT 46.74 1.845 47.04 2.115 ;
      RECT 46.775 1.826 46.861 2.165 ;
      RECT 44.87 1.74 45.04 2.935 ;
      RECT 44.87 1.74 45.335 1.91 ;
      RECT 44.87 6.97 45.335 7.14 ;
      RECT 44.87 5.945 45.04 7.14 ;
      RECT 43.88 1.74 44.05 2.935 ;
      RECT 43.88 1.74 44.345 1.91 ;
      RECT 43.88 6.97 44.345 7.14 ;
      RECT 43.88 5.945 44.05 7.14 ;
      RECT 42.025 2.635 42.195 3.865 ;
      RECT 42.08 0.855 42.25 2.805 ;
      RECT 42.025 0.575 42.195 1.025 ;
      RECT 42.025 7.855 42.195 8.305 ;
      RECT 42.08 6.075 42.25 8.025 ;
      RECT 42.025 5.015 42.195 6.245 ;
      RECT 41.505 0.575 41.675 3.865 ;
      RECT 41.505 2.075 41.91 2.405 ;
      RECT 41.505 1.235 41.91 1.565 ;
      RECT 41.505 5.015 41.675 8.305 ;
      RECT 41.505 7.315 41.91 7.645 ;
      RECT 41.505 6.475 41.91 6.805 ;
      RECT 39.43 3.126 39.435 3.298 ;
      RECT 39.425 3.119 39.43 3.388 ;
      RECT 39.42 3.113 39.425 3.407 ;
      RECT 39.4 3.107 39.42 3.417 ;
      RECT 39.385 3.102 39.4 3.425 ;
      RECT 39.348 3.096 39.385 3.423 ;
      RECT 39.262 3.082 39.348 3.419 ;
      RECT 39.176 3.064 39.262 3.414 ;
      RECT 39.09 3.045 39.176 3.408 ;
      RECT 39.06 3.033 39.09 3.404 ;
      RECT 39.04 3.027 39.06 3.403 ;
      RECT 38.975 3.025 39.04 3.401 ;
      RECT 38.96 3.025 38.975 3.393 ;
      RECT 38.945 3.025 38.96 3.38 ;
      RECT 38.94 3.025 38.945 3.37 ;
      RECT 38.925 3.025 38.94 3.348 ;
      RECT 38.91 3.025 38.925 3.315 ;
      RECT 38.905 3.025 38.91 3.293 ;
      RECT 38.895 3.025 38.905 3.275 ;
      RECT 38.88 3.025 38.895 3.253 ;
      RECT 38.86 3.025 38.88 3.215 ;
      RECT 39.21 2.31 39.245 2.749 ;
      RECT 39.21 2.31 39.25 2.748 ;
      RECT 39.155 2.37 39.25 2.747 ;
      RECT 39.02 2.542 39.25 2.746 ;
      RECT 39.13 2.42 39.25 2.746 ;
      RECT 39.02 2.542 39.275 2.736 ;
      RECT 39.075 2.487 39.355 2.653 ;
      RECT 39.25 2.281 39.255 2.744 ;
      RECT 39.105 2.457 39.395 2.53 ;
      RECT 39.12 2.44 39.25 2.746 ;
      RECT 39.255 2.28 39.425 2.468 ;
      RECT 39.245 2.283 39.425 2.468 ;
      RECT 38.75 2.16 38.92 2.47 ;
      RECT 38.75 2.16 38.925 2.443 ;
      RECT 38.75 2.16 38.93 2.42 ;
      RECT 38.75 2.16 38.94 2.37 ;
      RECT 38.745 2.265 38.94 2.34 ;
      RECT 38.78 1.835 38.95 2.313 ;
      RECT 38.78 1.835 38.965 2.234 ;
      RECT 38.77 2.045 38.965 2.234 ;
      RECT 38.78 1.845 38.975 2.149 ;
      RECT 38.71 2.587 38.715 2.79 ;
      RECT 38.7 2.575 38.71 2.9 ;
      RECT 38.675 2.575 38.7 2.94 ;
      RECT 38.595 2.575 38.675 3.025 ;
      RECT 38.585 2.575 38.595 3.095 ;
      RECT 38.56 2.575 38.585 3.118 ;
      RECT 38.54 2.575 38.56 3.153 ;
      RECT 38.495 2.585 38.54 3.196 ;
      RECT 38.485 2.597 38.495 3.233 ;
      RECT 38.465 2.611 38.485 3.253 ;
      RECT 38.455 2.629 38.465 3.269 ;
      RECT 38.44 2.655 38.455 3.279 ;
      RECT 38.425 2.696 38.44 3.293 ;
      RECT 38.415 2.731 38.425 3.303 ;
      RECT 38.41 2.747 38.415 3.308 ;
      RECT 38.4 2.762 38.41 3.313 ;
      RECT 38.38 2.805 38.4 3.323 ;
      RECT 38.36 2.842 38.38 3.336 ;
      RECT 38.325 2.865 38.36 3.354 ;
      RECT 38.315 2.879 38.325 3.37 ;
      RECT 38.295 2.889 38.315 3.38 ;
      RECT 38.29 2.898 38.295 3.388 ;
      RECT 38.28 2.905 38.29 3.395 ;
      RECT 38.27 2.912 38.28 3.403 ;
      RECT 38.255 2.922 38.27 3.411 ;
      RECT 38.245 2.936 38.255 3.421 ;
      RECT 38.235 2.948 38.245 3.433 ;
      RECT 38.22 2.97 38.235 3.446 ;
      RECT 38.21 2.992 38.22 3.457 ;
      RECT 38.2 3.012 38.21 3.466 ;
      RECT 38.195 3.027 38.2 3.473 ;
      RECT 38.165 3.06 38.195 3.487 ;
      RECT 38.155 3.095 38.165 3.502 ;
      RECT 38.15 3.102 38.155 3.508 ;
      RECT 38.13 3.117 38.15 3.515 ;
      RECT 38.125 3.132 38.13 3.523 ;
      RECT 38.12 3.141 38.125 3.528 ;
      RECT 38.105 3.147 38.12 3.535 ;
      RECT 38.1 3.153 38.105 3.543 ;
      RECT 38.095 3.157 38.1 3.55 ;
      RECT 38.09 3.161 38.095 3.56 ;
      RECT 38.08 3.166 38.09 3.57 ;
      RECT 38.06 3.177 38.08 3.598 ;
      RECT 38.045 3.189 38.06 3.625 ;
      RECT 38.025 3.202 38.045 3.65 ;
      RECT 38.005 3.217 38.025 3.674 ;
      RECT 37.99 3.232 38.005 3.689 ;
      RECT 37.985 3.243 37.99 3.698 ;
      RECT 37.92 3.288 37.985 3.708 ;
      RECT 37.885 3.347 37.92 3.721 ;
      RECT 37.88 3.37 37.885 3.727 ;
      RECT 37.875 3.377 37.88 3.729 ;
      RECT 37.86 3.387 37.875 3.732 ;
      RECT 37.83 3.412 37.86 3.736 ;
      RECT 37.825 3.43 37.83 3.74 ;
      RECT 37.82 3.437 37.825 3.741 ;
      RECT 37.8 3.445 37.82 3.745 ;
      RECT 37.79 3.452 37.8 3.749 ;
      RECT 37.746 3.463 37.79 3.756 ;
      RECT 37.66 3.491 37.746 3.772 ;
      RECT 37.6 3.515 37.66 3.79 ;
      RECT 37.555 3.525 37.6 3.804 ;
      RECT 37.496 3.533 37.555 3.818 ;
      RECT 37.41 3.54 37.496 3.837 ;
      RECT 37.385 3.545 37.41 3.852 ;
      RECT 37.305 3.548 37.385 3.855 ;
      RECT 37.225 3.552 37.305 3.842 ;
      RECT 37.216 3.555 37.225 3.827 ;
      RECT 37.13 3.555 37.216 3.812 ;
      RECT 37.07 3.557 37.13 3.789 ;
      RECT 37.066 3.56 37.07 3.779 ;
      RECT 36.98 3.56 37.066 3.764 ;
      RECT 36.905 3.56 36.98 3.74 ;
      RECT 38.22 2.569 38.23 2.745 ;
      RECT 38.175 2.536 38.22 2.745 ;
      RECT 38.13 2.487 38.175 2.745 ;
      RECT 38.1 2.457 38.13 2.746 ;
      RECT 38.095 2.44 38.1 2.747 ;
      RECT 38.07 2.42 38.095 2.748 ;
      RECT 38.055 2.395 38.07 2.749 ;
      RECT 38.05 2.382 38.055 2.75 ;
      RECT 38.045 2.376 38.05 2.748 ;
      RECT 38.04 2.368 38.045 2.742 ;
      RECT 38.015 2.36 38.04 2.722 ;
      RECT 37.995 2.349 38.015 2.693 ;
      RECT 37.965 2.334 37.995 2.664 ;
      RECT 37.945 2.32 37.965 2.636 ;
      RECT 37.935 2.314 37.945 2.615 ;
      RECT 37.93 2.311 37.935 2.598 ;
      RECT 37.925 2.308 37.93 2.583 ;
      RECT 37.91 2.303 37.925 2.548 ;
      RECT 37.905 2.299 37.91 2.515 ;
      RECT 37.885 2.294 37.905 2.491 ;
      RECT 37.855 2.286 37.885 2.456 ;
      RECT 37.84 2.28 37.855 2.433 ;
      RECT 37.8 2.273 37.84 2.418 ;
      RECT 37.775 2.265 37.8 2.398 ;
      RECT 37.755 2.26 37.775 2.388 ;
      RECT 37.72 2.254 37.755 2.383 ;
      RECT 37.675 2.245 37.72 2.382 ;
      RECT 37.645 2.241 37.675 2.384 ;
      RECT 37.56 2.249 37.645 2.388 ;
      RECT 37.49 2.26 37.56 2.41 ;
      RECT 37.477 2.266 37.49 2.433 ;
      RECT 37.391 2.273 37.477 2.455 ;
      RECT 37.305 2.285 37.391 2.492 ;
      RECT 37.305 2.662 37.315 2.9 ;
      RECT 37.3 2.291 37.305 2.515 ;
      RECT 37.295 2.547 37.305 2.9 ;
      RECT 37.295 2.292 37.3 2.52 ;
      RECT 37.29 2.293 37.295 2.9 ;
      RECT 37.266 2.295 37.29 2.901 ;
      RECT 37.18 2.303 37.266 2.903 ;
      RECT 37.16 2.317 37.18 2.906 ;
      RECT 37.155 2.345 37.16 2.907 ;
      RECT 37.15 2.357 37.155 2.908 ;
      RECT 37.145 2.372 37.15 2.909 ;
      RECT 37.135 2.402 37.145 2.91 ;
      RECT 37.13 2.44 37.135 2.908 ;
      RECT 37.125 2.46 37.13 2.903 ;
      RECT 37.11 2.495 37.125 2.888 ;
      RECT 37.1 2.547 37.11 2.868 ;
      RECT 37.095 2.577 37.1 2.856 ;
      RECT 37.08 2.59 37.095 2.839 ;
      RECT 37.055 2.594 37.08 2.806 ;
      RECT 37.04 2.592 37.055 2.783 ;
      RECT 37.025 2.591 37.04 2.78 ;
      RECT 36.965 2.589 37.025 2.778 ;
      RECT 36.955 2.587 36.965 2.773 ;
      RECT 36.915 2.586 36.955 2.77 ;
      RECT 36.845 2.583 36.915 2.768 ;
      RECT 36.79 2.581 36.845 2.763 ;
      RECT 36.72 2.575 36.79 2.758 ;
      RECT 36.711 2.575 36.72 2.755 ;
      RECT 36.625 2.575 36.711 2.75 ;
      RECT 36.62 2.575 36.625 2.745 ;
      RECT 37.925 1.81 38.1 2.16 ;
      RECT 37.925 1.825 38.11 2.158 ;
      RECT 37.9 1.775 38.045 2.155 ;
      RECT 37.88 1.776 38.045 2.148 ;
      RECT 37.87 1.777 38.055 2.143 ;
      RECT 37.84 1.778 38.055 2.13 ;
      RECT 37.79 1.779 38.055 2.106 ;
      RECT 37.785 1.781 38.055 2.091 ;
      RECT 37.785 1.847 38.115 2.085 ;
      RECT 37.765 1.788 38.07 2.065 ;
      RECT 37.755 1.797 38.08 1.92 ;
      RECT 37.765 1.792 38.08 2.065 ;
      RECT 37.785 1.782 38.07 2.091 ;
      RECT 37.37 3.107 37.54 3.395 ;
      RECT 37.365 3.125 37.55 3.39 ;
      RECT 37.33 3.133 37.615 3.31 ;
      RECT 37.33 3.133 37.701 3.3 ;
      RECT 37.33 3.133 37.755 3.246 ;
      RECT 37.615 3.03 37.785 3.214 ;
      RECT 37.33 3.185 37.79 3.202 ;
      RECT 37.315 3.155 37.785 3.198 ;
      RECT 37.575 3.037 37.615 3.349 ;
      RECT 37.455 3.074 37.785 3.214 ;
      RECT 37.55 3.049 37.575 3.375 ;
      RECT 37.54 3.056 37.785 3.214 ;
      RECT 37.671 2.52 37.74 2.779 ;
      RECT 37.671 2.575 37.745 2.778 ;
      RECT 37.585 2.575 37.745 2.777 ;
      RECT 37.58 2.575 37.75 2.77 ;
      RECT 37.57 2.52 37.74 2.765 ;
      RECT 36.95 1.819 37.125 2.12 ;
      RECT 36.935 1.807 36.95 2.105 ;
      RECT 36.905 1.806 36.935 2.058 ;
      RECT 36.905 1.824 37.13 2.053 ;
      RECT 36.89 1.808 36.95 2.018 ;
      RECT 36.885 1.83 37.14 1.918 ;
      RECT 36.885 1.813 37.036 1.918 ;
      RECT 36.885 1.815 37.04 1.918 ;
      RECT 36.89 1.811 37.036 2.018 ;
      RECT 36.995 3.047 37 3.395 ;
      RECT 36.985 3.037 36.995 3.401 ;
      RECT 36.95 3.027 36.985 3.403 ;
      RECT 36.912 3.022 36.95 3.407 ;
      RECT 36.826 3.015 36.912 3.414 ;
      RECT 36.74 3.005 36.826 3.424 ;
      RECT 36.695 3 36.74 3.432 ;
      RECT 36.691 3 36.695 3.436 ;
      RECT 36.605 3 36.691 3.443 ;
      RECT 36.59 3 36.605 3.443 ;
      RECT 36.58 2.998 36.59 3.415 ;
      RECT 36.57 2.994 36.58 3.358 ;
      RECT 36.55 2.988 36.57 3.29 ;
      RECT 36.545 2.984 36.55 3.238 ;
      RECT 36.535 2.983 36.545 3.205 ;
      RECT 36.485 2.981 36.535 3.19 ;
      RECT 36.46 2.979 36.485 3.185 ;
      RECT 36.417 2.977 36.46 3.181 ;
      RECT 36.331 2.973 36.417 3.169 ;
      RECT 36.245 2.968 36.331 3.153 ;
      RECT 36.215 2.965 36.245 3.14 ;
      RECT 36.19 2.964 36.215 3.128 ;
      RECT 36.185 2.964 36.19 3.118 ;
      RECT 36.145 2.963 36.185 3.11 ;
      RECT 36.13 2.962 36.145 3.103 ;
      RECT 36.08 2.961 36.13 3.095 ;
      RECT 36.078 2.96 36.08 3.09 ;
      RECT 35.992 2.958 36.078 3.09 ;
      RECT 35.906 2.953 35.992 3.09 ;
      RECT 35.82 2.949 35.906 3.09 ;
      RECT 35.771 2.945 35.82 3.088 ;
      RECT 35.685 2.942 35.771 3.083 ;
      RECT 35.662 2.939 35.685 3.079 ;
      RECT 35.576 2.936 35.662 3.074 ;
      RECT 35.49 2.932 35.576 3.065 ;
      RECT 35.465 2.925 35.49 3.06 ;
      RECT 35.405 2.89 35.465 3.057 ;
      RECT 35.385 2.815 35.405 3.054 ;
      RECT 35.38 2.757 35.385 3.053 ;
      RECT 35.355 2.697 35.38 3.052 ;
      RECT 35.28 2.575 35.355 3.048 ;
      RECT 35.27 2.575 35.28 3.04 ;
      RECT 35.255 2.575 35.27 3.03 ;
      RECT 35.24 2.575 35.255 3 ;
      RECT 35.225 2.575 35.24 2.945 ;
      RECT 35.21 2.575 35.225 2.883 ;
      RECT 35.185 2.575 35.21 2.808 ;
      RECT 35.18 2.575 35.185 2.758 ;
      RECT 36.525 2.12 36.545 2.429 ;
      RECT 36.511 2.122 36.56 2.426 ;
      RECT 36.511 2.127 36.58 2.417 ;
      RECT 36.425 2.125 36.56 2.411 ;
      RECT 36.425 2.133 36.615 2.394 ;
      RECT 36.39 2.135 36.615 2.393 ;
      RECT 36.36 2.143 36.615 2.384 ;
      RECT 36.35 2.148 36.635 2.37 ;
      RECT 36.39 2.138 36.635 2.37 ;
      RECT 36.39 2.141 36.645 2.358 ;
      RECT 36.36 2.143 36.655 2.345 ;
      RECT 36.36 2.147 36.665 2.288 ;
      RECT 36.35 2.152 36.67 2.203 ;
      RECT 36.511 2.12 36.545 2.426 ;
      RECT 35.95 2.223 35.955 2.435 ;
      RECT 35.825 2.22 35.84 2.435 ;
      RECT 35.29 2.25 35.36 2.435 ;
      RECT 35.175 2.25 35.21 2.43 ;
      RECT 36.296 2.552 36.315 2.746 ;
      RECT 36.21 2.507 36.296 2.747 ;
      RECT 36.2 2.46 36.21 2.749 ;
      RECT 36.195 2.44 36.2 2.75 ;
      RECT 36.175 2.405 36.195 2.751 ;
      RECT 36.16 2.355 36.175 2.752 ;
      RECT 36.14 2.292 36.16 2.753 ;
      RECT 36.13 2.255 36.14 2.754 ;
      RECT 36.115 2.244 36.13 2.755 ;
      RECT 36.11 2.236 36.115 2.753 ;
      RECT 36.1 2.235 36.11 2.745 ;
      RECT 36.07 2.232 36.1 2.724 ;
      RECT 35.995 2.227 36.07 2.669 ;
      RECT 35.98 2.223 35.995 2.615 ;
      RECT 35.97 2.223 35.98 2.51 ;
      RECT 35.955 2.223 35.97 2.443 ;
      RECT 35.94 2.223 35.95 2.433 ;
      RECT 35.885 2.222 35.94 2.43 ;
      RECT 35.84 2.22 35.885 2.433 ;
      RECT 35.812 2.22 35.825 2.436 ;
      RECT 35.726 2.224 35.812 2.438 ;
      RECT 35.64 2.23 35.726 2.443 ;
      RECT 35.62 2.234 35.64 2.445 ;
      RECT 35.618 2.235 35.62 2.444 ;
      RECT 35.532 2.237 35.618 2.443 ;
      RECT 35.446 2.242 35.532 2.44 ;
      RECT 35.36 2.247 35.446 2.437 ;
      RECT 35.21 2.25 35.29 2.433 ;
      RECT 35.986 3.225 36.035 3.559 ;
      RECT 35.986 3.225 36.04 3.558 ;
      RECT 35.9 3.225 36.04 3.557 ;
      RECT 35.675 3.333 36.045 3.555 ;
      RECT 35.9 3.225 36.07 3.548 ;
      RECT 35.87 3.237 36.075 3.539 ;
      RECT 35.855 3.255 36.08 3.536 ;
      RECT 35.67 3.339 36.08 3.463 ;
      RECT 35.665 3.346 36.08 3.423 ;
      RECT 35.68 3.312 36.08 3.536 ;
      RECT 35.841 3.258 36.045 3.555 ;
      RECT 35.755 3.278 36.08 3.536 ;
      RECT 35.855 3.252 36.075 3.539 ;
      RECT 35.625 2.576 35.815 2.77 ;
      RECT 35.62 2.578 35.815 2.769 ;
      RECT 35.615 2.582 35.83 2.766 ;
      RECT 35.63 2.575 35.83 2.766 ;
      RECT 35.615 2.685 35.835 2.761 ;
      RECT 34.91 3.185 35.001 3.483 ;
      RECT 34.905 3.187 35.08 3.478 ;
      RECT 34.91 3.185 35.08 3.478 ;
      RECT 34.905 3.191 35.1 3.476 ;
      RECT 34.905 3.246 35.14 3.475 ;
      RECT 34.905 3.281 35.155 3.469 ;
      RECT 34.905 3.315 35.165 3.459 ;
      RECT 34.895 3.195 35.1 3.31 ;
      RECT 34.895 3.215 35.115 3.31 ;
      RECT 34.895 3.198 35.105 3.31 ;
      RECT 35.12 1.966 35.125 2.028 ;
      RECT 35.115 1.888 35.12 2.051 ;
      RECT 35.11 1.845 35.115 2.062 ;
      RECT 35.105 1.835 35.11 2.074 ;
      RECT 35.1 1.835 35.105 2.083 ;
      RECT 35.075 1.835 35.1 2.115 ;
      RECT 35.07 1.835 35.075 2.148 ;
      RECT 35.055 1.835 35.07 2.173 ;
      RECT 35.045 1.835 35.055 2.2 ;
      RECT 35.04 1.835 35.045 2.213 ;
      RECT 35.035 1.835 35.04 2.228 ;
      RECT 35.025 1.835 35.035 2.243 ;
      RECT 35.02 1.835 35.025 2.263 ;
      RECT 34.995 1.835 35.02 2.298 ;
      RECT 34.95 1.835 34.995 2.343 ;
      RECT 34.94 1.835 34.95 2.356 ;
      RECT 34.855 1.92 34.94 2.363 ;
      RECT 34.82 2.042 34.855 2.372 ;
      RECT 34.815 2.082 34.82 2.376 ;
      RECT 34.795 2.105 34.815 2.378 ;
      RECT 34.79 2.135 34.795 2.381 ;
      RECT 34.78 2.147 34.79 2.382 ;
      RECT 34.735 2.17 34.78 2.387 ;
      RECT 34.695 2.2 34.735 2.395 ;
      RECT 34.66 2.212 34.695 2.401 ;
      RECT 34.655 2.217 34.66 2.405 ;
      RECT 34.585 2.227 34.655 2.412 ;
      RECT 34.545 2.237 34.585 2.422 ;
      RECT 34.525 2.242 34.545 2.428 ;
      RECT 34.515 2.246 34.525 2.433 ;
      RECT 34.51 2.249 34.515 2.436 ;
      RECT 34.5 2.25 34.51 2.437 ;
      RECT 34.475 2.252 34.5 2.441 ;
      RECT 34.465 2.257 34.475 2.444 ;
      RECT 34.42 2.265 34.465 2.445 ;
      RECT 34.295 2.27 34.42 2.445 ;
      RECT 34.85 2.567 34.87 2.749 ;
      RECT 34.801 2.552 34.85 2.748 ;
      RECT 34.715 2.567 34.87 2.746 ;
      RECT 34.7 2.567 34.87 2.745 ;
      RECT 34.665 2.545 34.835 2.73 ;
      RECT 34.735 3.565 34.75 3.774 ;
      RECT 34.735 3.573 34.755 3.773 ;
      RECT 34.68 3.573 34.755 3.772 ;
      RECT 34.66 3.577 34.76 3.77 ;
      RECT 34.64 3.527 34.68 3.769 ;
      RECT 34.585 3.585 34.765 3.767 ;
      RECT 34.55 3.542 34.68 3.765 ;
      RECT 34.546 3.545 34.735 3.764 ;
      RECT 34.46 3.553 34.735 3.762 ;
      RECT 34.46 3.597 34.77 3.755 ;
      RECT 34.45 3.69 34.77 3.753 ;
      RECT 34.46 3.609 34.775 3.738 ;
      RECT 34.46 3.63 34.79 3.708 ;
      RECT 34.46 3.657 34.795 3.678 ;
      RECT 34.585 3.535 34.68 3.767 ;
      RECT 34.215 2.58 34.22 3.118 ;
      RECT 34.02 2.91 34.025 3.105 ;
      RECT 32.32 2.575 32.335 2.955 ;
      RECT 34.385 2.575 34.39 2.745 ;
      RECT 34.38 2.575 34.385 2.755 ;
      RECT 34.375 2.575 34.38 2.768 ;
      RECT 34.35 2.575 34.375 2.81 ;
      RECT 34.325 2.575 34.35 2.883 ;
      RECT 34.31 2.575 34.325 2.935 ;
      RECT 34.305 2.575 34.31 2.965 ;
      RECT 34.28 2.575 34.305 3.005 ;
      RECT 34.265 2.575 34.28 3.06 ;
      RECT 34.26 2.575 34.265 3.093 ;
      RECT 34.235 2.575 34.26 3.113 ;
      RECT 34.22 2.575 34.235 3.119 ;
      RECT 34.15 2.61 34.215 3.115 ;
      RECT 34.1 2.665 34.15 3.11 ;
      RECT 34.09 2.697 34.1 3.108 ;
      RECT 34.085 2.722 34.09 3.108 ;
      RECT 34.065 2.795 34.085 3.108 ;
      RECT 34.055 2.875 34.065 3.107 ;
      RECT 34.04 2.905 34.055 3.107 ;
      RECT 34.025 2.91 34.04 3.106 ;
      RECT 33.965 2.912 34.02 3.103 ;
      RECT 33.935 2.917 33.965 3.099 ;
      RECT 33.933 2.92 33.935 3.098 ;
      RECT 33.847 2.922 33.933 3.095 ;
      RECT 33.761 2.928 33.847 3.089 ;
      RECT 33.675 2.933 33.761 3.083 ;
      RECT 33.602 2.938 33.675 3.084 ;
      RECT 33.516 2.944 33.602 3.092 ;
      RECT 33.43 2.95 33.516 3.101 ;
      RECT 33.41 2.954 33.43 3.106 ;
      RECT 33.363 2.956 33.41 3.109 ;
      RECT 33.277 2.961 33.363 3.115 ;
      RECT 33.191 2.966 33.277 3.124 ;
      RECT 33.105 2.972 33.191 3.132 ;
      RECT 33.02 2.97 33.105 3.141 ;
      RECT 33.016 2.965 33.02 3.145 ;
      RECT 32.93 2.96 33.016 3.137 ;
      RECT 32.866 2.951 32.93 3.125 ;
      RECT 32.78 2.942 32.866 3.112 ;
      RECT 32.756 2.935 32.78 3.103 ;
      RECT 32.67 2.929 32.756 3.09 ;
      RECT 32.63 2.922 32.67 3.076 ;
      RECT 32.625 2.912 32.63 3.072 ;
      RECT 32.615 2.9 32.625 3.071 ;
      RECT 32.595 2.87 32.615 3.068 ;
      RECT 32.54 2.79 32.595 3.062 ;
      RECT 32.52 2.709 32.54 3.057 ;
      RECT 32.5 2.667 32.52 3.053 ;
      RECT 32.475 2.62 32.5 3.047 ;
      RECT 32.47 2.595 32.475 3.044 ;
      RECT 32.435 2.575 32.47 3.039 ;
      RECT 32.426 2.575 32.435 3.032 ;
      RECT 32.34 2.575 32.426 3.002 ;
      RECT 32.335 2.575 32.34 2.965 ;
      RECT 32.3 2.575 32.32 2.887 ;
      RECT 32.295 2.617 32.3 2.852 ;
      RECT 32.29 2.692 32.295 2.808 ;
      RECT 33.74 2.497 33.915 2.745 ;
      RECT 33.74 2.497 33.92 2.743 ;
      RECT 33.735 2.529 33.92 2.703 ;
      RECT 33.765 2.47 33.935 2.69 ;
      RECT 33.73 2.547 33.935 2.623 ;
      RECT 33.04 2.01 33.21 2.185 ;
      RECT 33.04 2.01 33.382 2.177 ;
      RECT 33.04 2.01 33.465 2.171 ;
      RECT 33.04 2.01 33.5 2.167 ;
      RECT 33.04 2.01 33.52 2.166 ;
      RECT 33.04 2.01 33.606 2.162 ;
      RECT 33.5 1.835 33.67 2.157 ;
      RECT 33.075 1.942 33.7 2.155 ;
      RECT 33.065 1.997 33.705 2.153 ;
      RECT 33.04 2.033 33.715 2.148 ;
      RECT 33.04 2.06 33.72 2.078 ;
      RECT 33.105 1.885 33.68 2.155 ;
      RECT 33.296 1.87 33.68 2.155 ;
      RECT 33.13 1.873 33.68 2.155 ;
      RECT 33.21 1.871 33.296 2.182 ;
      RECT 33.296 1.868 33.675 2.155 ;
      RECT 33.48 1.845 33.675 2.155 ;
      RECT 33.382 1.866 33.675 2.155 ;
      RECT 33.465 1.86 33.48 2.168 ;
      RECT 33.615 3.225 33.62 3.425 ;
      RECT 33.08 3.29 33.125 3.425 ;
      RECT 33.65 3.225 33.67 3.398 ;
      RECT 33.62 3.225 33.65 3.413 ;
      RECT 33.555 3.225 33.615 3.45 ;
      RECT 33.54 3.225 33.555 3.48 ;
      RECT 33.525 3.225 33.54 3.493 ;
      RECT 33.505 3.225 33.525 3.508 ;
      RECT 33.5 3.225 33.505 3.517 ;
      RECT 33.49 3.229 33.5 3.522 ;
      RECT 33.475 3.239 33.49 3.533 ;
      RECT 33.45 3.255 33.475 3.543 ;
      RECT 33.44 3.269 33.45 3.545 ;
      RECT 33.42 3.281 33.44 3.542 ;
      RECT 33.39 3.302 33.42 3.536 ;
      RECT 33.38 3.314 33.39 3.531 ;
      RECT 33.37 3.312 33.38 3.528 ;
      RECT 33.355 3.311 33.37 3.523 ;
      RECT 33.35 3.31 33.355 3.518 ;
      RECT 33.315 3.308 33.35 3.508 ;
      RECT 33.295 3.305 33.315 3.49 ;
      RECT 33.285 3.303 33.295 3.485 ;
      RECT 33.275 3.302 33.285 3.48 ;
      RECT 33.24 3.3 33.275 3.468 ;
      RECT 33.185 3.296 33.24 3.448 ;
      RECT 33.175 3.294 33.185 3.433 ;
      RECT 33.17 3.294 33.175 3.428 ;
      RECT 33.125 3.292 33.17 3.425 ;
      RECT 33.03 3.29 33.08 3.429 ;
      RECT 33.02 3.291 33.03 3.434 ;
      RECT 32.96 3.298 33.02 3.448 ;
      RECT 32.935 3.306 32.96 3.468 ;
      RECT 32.925 3.31 32.935 3.48 ;
      RECT 32.92 3.311 32.925 3.485 ;
      RECT 32.905 3.313 32.92 3.488 ;
      RECT 32.89 3.315 32.905 3.493 ;
      RECT 32.885 3.315 32.89 3.496 ;
      RECT 32.84 3.32 32.885 3.507 ;
      RECT 32.835 3.324 32.84 3.519 ;
      RECT 32.81 3.32 32.835 3.523 ;
      RECT 32.8 3.316 32.81 3.527 ;
      RECT 32.79 3.315 32.8 3.531 ;
      RECT 32.775 3.305 32.79 3.537 ;
      RECT 32.77 3.293 32.775 3.541 ;
      RECT 32.765 3.29 32.77 3.542 ;
      RECT 32.76 3.287 32.765 3.544 ;
      RECT 32.745 3.275 32.76 3.543 ;
      RECT 32.73 3.257 32.745 3.54 ;
      RECT 32.71 3.236 32.73 3.533 ;
      RECT 32.645 3.225 32.71 3.505 ;
      RECT 32.641 3.225 32.645 3.484 ;
      RECT 32.555 3.225 32.641 3.454 ;
      RECT 32.54 3.225 32.555 3.41 ;
      RECT 33.115 2.325 33.12 2.56 ;
      RECT 32.245 2.241 32.25 2.445 ;
      RECT 32.825 2.27 32.83 2.425 ;
      RECT 32.745 2.25 32.75 2.425 ;
      RECT 33.415 2.392 33.43 2.745 ;
      RECT 33.341 2.377 33.415 2.745 ;
      RECT 33.255 2.36 33.341 2.745 ;
      RECT 33.245 2.35 33.255 2.743 ;
      RECT 33.24 2.348 33.245 2.738 ;
      RECT 33.225 2.346 33.24 2.724 ;
      RECT 33.155 2.338 33.225 2.664 ;
      RECT 33.135 2.329 33.155 2.598 ;
      RECT 33.13 2.326 33.135 2.578 ;
      RECT 33.12 2.325 33.13 2.568 ;
      RECT 33.11 2.325 33.115 2.552 ;
      RECT 33.1 2.324 33.11 2.542 ;
      RECT 33.09 2.322 33.1 2.53 ;
      RECT 33.075 2.319 33.09 2.51 ;
      RECT 33.065 2.317 33.075 2.495 ;
      RECT 33.045 2.314 33.065 2.483 ;
      RECT 33.04 2.312 33.045 2.473 ;
      RECT 33.015 2.31 33.04 2.46 ;
      RECT 32.985 2.305 33.015 2.445 ;
      RECT 32.905 2.296 32.985 2.436 ;
      RECT 32.86 2.285 32.905 2.429 ;
      RECT 32.84 2.276 32.86 2.426 ;
      RECT 32.83 2.271 32.84 2.425 ;
      RECT 32.785 2.265 32.825 2.425 ;
      RECT 32.77 2.257 32.785 2.425 ;
      RECT 32.75 2.252 32.77 2.425 ;
      RECT 32.73 2.249 32.745 2.425 ;
      RECT 32.647 2.248 32.73 2.424 ;
      RECT 32.561 2.247 32.647 2.42 ;
      RECT 32.475 2.245 32.561 2.417 ;
      RECT 32.422 2.244 32.475 2.419 ;
      RECT 32.336 2.243 32.422 2.428 ;
      RECT 32.25 2.242 32.336 2.44 ;
      RECT 32.23 2.241 32.245 2.448 ;
      RECT 32.15 2.24 32.23 2.46 ;
      RECT 32.125 2.24 32.15 2.473 ;
      RECT 32.1 2.24 32.125 2.488 ;
      RECT 32.095 2.24 32.1 2.51 ;
      RECT 32.09 2.24 32.095 2.528 ;
      RECT 32.085 2.24 32.09 2.545 ;
      RECT 32.08 2.24 32.085 2.558 ;
      RECT 32.075 2.24 32.08 2.568 ;
      RECT 32.035 2.24 32.075 2.653 ;
      RECT 32.02 2.24 32.035 2.738 ;
      RECT 32.01 2.241 32.02 2.75 ;
      RECT 31.975 2.246 32.01 2.755 ;
      RECT 31.935 2.255 31.975 2.755 ;
      RECT 31.92 2.265 31.935 2.755 ;
      RECT 31.915 2.275 31.92 2.755 ;
      RECT 31.895 2.302 31.915 2.755 ;
      RECT 31.845 2.385 31.895 2.755 ;
      RECT 31.84 2.447 31.845 2.755 ;
      RECT 31.83 2.46 31.84 2.755 ;
      RECT 31.82 2.482 31.83 2.755 ;
      RECT 31.81 2.507 31.82 2.75 ;
      RECT 31.805 2.545 31.81 2.743 ;
      RECT 31.795 2.655 31.805 2.738 ;
      RECT 33.19 3.576 33.205 3.835 ;
      RECT 33.19 3.591 33.21 3.834 ;
      RECT 33.106 3.591 33.21 3.832 ;
      RECT 33.106 3.605 33.215 3.831 ;
      RECT 33.02 3.647 33.22 3.828 ;
      RECT 33.015 3.59 33.205 3.823 ;
      RECT 33.015 3.661 33.225 3.82 ;
      RECT 33.01 3.692 33.225 3.818 ;
      RECT 33.015 3.689 33.24 3.808 ;
      RECT 33.01 3.735 33.255 3.793 ;
      RECT 33.01 3.763 33.26 3.778 ;
      RECT 33.02 3.565 33.19 3.828 ;
      RECT 32.78 2.575 32.95 2.745 ;
      RECT 32.745 2.575 32.95 2.74 ;
      RECT 32.735 2.575 32.95 2.733 ;
      RECT 32.73 2.56 32.9 2.73 ;
      RECT 31.56 3.097 31.825 3.54 ;
      RECT 31.555 3.068 31.77 3.538 ;
      RECT 31.55 3.222 31.83 3.533 ;
      RECT 31.555 3.117 31.83 3.533 ;
      RECT 31.555 3.128 31.84 3.52 ;
      RECT 31.555 3.075 31.8 3.538 ;
      RECT 31.56 3.062 31.77 3.54 ;
      RECT 31.56 3.06 31.72 3.54 ;
      RECT 31.661 3.052 31.72 3.54 ;
      RECT 31.575 3.053 31.72 3.54 ;
      RECT 31.661 3.051 31.71 3.54 ;
      RECT 31.465 1.866 31.64 2.165 ;
      RECT 31.515 1.828 31.64 2.165 ;
      RECT 31.5 1.83 31.726 2.157 ;
      RECT 31.5 1.833 31.765 2.144 ;
      RECT 31.5 1.834 31.775 2.13 ;
      RECT 31.455 1.885 31.775 2.12 ;
      RECT 31.5 1.835 31.78 2.115 ;
      RECT 31.455 2.045 31.785 2.105 ;
      RECT 31.44 1.905 31.78 2.045 ;
      RECT 31.435 1.921 31.78 1.985 ;
      RECT 31.48 1.845 31.78 2.115 ;
      RECT 31.515 1.826 31.601 2.165 ;
      RECT 29.61 1.74 29.78 2.935 ;
      RECT 29.61 1.74 30.075 1.91 ;
      RECT 29.61 6.97 30.075 7.14 ;
      RECT 29.61 5.945 29.78 7.14 ;
      RECT 28.62 1.74 28.79 2.935 ;
      RECT 28.62 1.74 29.085 1.91 ;
      RECT 28.62 6.97 29.085 7.14 ;
      RECT 28.62 5.945 28.79 7.14 ;
      RECT 26.765 2.635 26.935 3.865 ;
      RECT 26.82 0.855 26.99 2.805 ;
      RECT 26.765 0.575 26.935 1.025 ;
      RECT 26.765 7.855 26.935 8.305 ;
      RECT 26.82 6.075 26.99 8.025 ;
      RECT 26.765 5.015 26.935 6.245 ;
      RECT 26.245 0.575 26.415 3.865 ;
      RECT 26.245 2.075 26.65 2.405 ;
      RECT 26.245 1.235 26.65 1.565 ;
      RECT 26.245 5.015 26.415 8.305 ;
      RECT 26.245 7.315 26.65 7.645 ;
      RECT 26.245 6.475 26.65 6.805 ;
      RECT 24.17 3.126 24.175 3.298 ;
      RECT 24.165 3.119 24.17 3.388 ;
      RECT 24.16 3.113 24.165 3.407 ;
      RECT 24.14 3.107 24.16 3.417 ;
      RECT 24.125 3.102 24.14 3.425 ;
      RECT 24.088 3.096 24.125 3.423 ;
      RECT 24.002 3.082 24.088 3.419 ;
      RECT 23.916 3.064 24.002 3.414 ;
      RECT 23.83 3.045 23.916 3.408 ;
      RECT 23.8 3.033 23.83 3.404 ;
      RECT 23.78 3.027 23.8 3.403 ;
      RECT 23.715 3.025 23.78 3.401 ;
      RECT 23.7 3.025 23.715 3.393 ;
      RECT 23.685 3.025 23.7 3.38 ;
      RECT 23.68 3.025 23.685 3.37 ;
      RECT 23.665 3.025 23.68 3.348 ;
      RECT 23.65 3.025 23.665 3.315 ;
      RECT 23.645 3.025 23.65 3.293 ;
      RECT 23.635 3.025 23.645 3.275 ;
      RECT 23.62 3.025 23.635 3.253 ;
      RECT 23.6 3.025 23.62 3.215 ;
      RECT 23.95 2.31 23.985 2.749 ;
      RECT 23.95 2.31 23.99 2.748 ;
      RECT 23.895 2.37 23.99 2.747 ;
      RECT 23.76 2.542 23.99 2.746 ;
      RECT 23.87 2.42 23.99 2.746 ;
      RECT 23.76 2.542 24.015 2.736 ;
      RECT 23.815 2.487 24.095 2.653 ;
      RECT 23.99 2.281 23.995 2.744 ;
      RECT 23.845 2.457 24.135 2.53 ;
      RECT 23.86 2.44 23.99 2.746 ;
      RECT 23.995 2.28 24.165 2.468 ;
      RECT 23.985 2.283 24.165 2.468 ;
      RECT 23.49 2.16 23.66 2.47 ;
      RECT 23.49 2.16 23.665 2.443 ;
      RECT 23.49 2.16 23.67 2.42 ;
      RECT 23.49 2.16 23.68 2.37 ;
      RECT 23.485 2.265 23.68 2.34 ;
      RECT 23.52 1.835 23.69 2.313 ;
      RECT 23.52 1.835 23.705 2.234 ;
      RECT 23.51 2.045 23.705 2.234 ;
      RECT 23.52 1.845 23.715 2.149 ;
      RECT 23.45 2.587 23.455 2.79 ;
      RECT 23.44 2.575 23.45 2.9 ;
      RECT 23.415 2.575 23.44 2.94 ;
      RECT 23.335 2.575 23.415 3.025 ;
      RECT 23.325 2.575 23.335 3.095 ;
      RECT 23.3 2.575 23.325 3.118 ;
      RECT 23.28 2.575 23.3 3.153 ;
      RECT 23.235 2.585 23.28 3.196 ;
      RECT 23.225 2.597 23.235 3.233 ;
      RECT 23.205 2.611 23.225 3.253 ;
      RECT 23.195 2.629 23.205 3.269 ;
      RECT 23.18 2.655 23.195 3.279 ;
      RECT 23.165 2.696 23.18 3.293 ;
      RECT 23.155 2.731 23.165 3.303 ;
      RECT 23.15 2.747 23.155 3.308 ;
      RECT 23.14 2.762 23.15 3.313 ;
      RECT 23.12 2.805 23.14 3.323 ;
      RECT 23.1 2.842 23.12 3.336 ;
      RECT 23.065 2.865 23.1 3.354 ;
      RECT 23.055 2.879 23.065 3.37 ;
      RECT 23.035 2.889 23.055 3.38 ;
      RECT 23.03 2.898 23.035 3.388 ;
      RECT 23.02 2.905 23.03 3.395 ;
      RECT 23.01 2.912 23.02 3.403 ;
      RECT 22.995 2.922 23.01 3.411 ;
      RECT 22.985 2.936 22.995 3.421 ;
      RECT 22.975 2.948 22.985 3.433 ;
      RECT 22.96 2.97 22.975 3.446 ;
      RECT 22.95 2.992 22.96 3.457 ;
      RECT 22.94 3.012 22.95 3.466 ;
      RECT 22.935 3.027 22.94 3.473 ;
      RECT 22.905 3.06 22.935 3.487 ;
      RECT 22.895 3.095 22.905 3.502 ;
      RECT 22.89 3.102 22.895 3.508 ;
      RECT 22.87 3.117 22.89 3.515 ;
      RECT 22.865 3.132 22.87 3.523 ;
      RECT 22.86 3.141 22.865 3.528 ;
      RECT 22.845 3.147 22.86 3.535 ;
      RECT 22.84 3.153 22.845 3.543 ;
      RECT 22.835 3.157 22.84 3.55 ;
      RECT 22.83 3.161 22.835 3.56 ;
      RECT 22.82 3.166 22.83 3.57 ;
      RECT 22.8 3.177 22.82 3.598 ;
      RECT 22.785 3.189 22.8 3.625 ;
      RECT 22.765 3.202 22.785 3.65 ;
      RECT 22.745 3.217 22.765 3.674 ;
      RECT 22.73 3.232 22.745 3.689 ;
      RECT 22.725 3.243 22.73 3.698 ;
      RECT 22.66 3.288 22.725 3.708 ;
      RECT 22.625 3.347 22.66 3.721 ;
      RECT 22.62 3.37 22.625 3.727 ;
      RECT 22.615 3.377 22.62 3.729 ;
      RECT 22.6 3.387 22.615 3.732 ;
      RECT 22.57 3.412 22.6 3.736 ;
      RECT 22.565 3.43 22.57 3.74 ;
      RECT 22.56 3.437 22.565 3.741 ;
      RECT 22.54 3.445 22.56 3.745 ;
      RECT 22.53 3.452 22.54 3.749 ;
      RECT 22.486 3.463 22.53 3.756 ;
      RECT 22.4 3.491 22.486 3.772 ;
      RECT 22.34 3.515 22.4 3.79 ;
      RECT 22.295 3.525 22.34 3.804 ;
      RECT 22.236 3.533 22.295 3.818 ;
      RECT 22.15 3.54 22.236 3.837 ;
      RECT 22.125 3.545 22.15 3.852 ;
      RECT 22.045 3.548 22.125 3.855 ;
      RECT 21.965 3.552 22.045 3.842 ;
      RECT 21.956 3.555 21.965 3.827 ;
      RECT 21.87 3.555 21.956 3.812 ;
      RECT 21.81 3.557 21.87 3.789 ;
      RECT 21.806 3.56 21.81 3.779 ;
      RECT 21.72 3.56 21.806 3.764 ;
      RECT 21.645 3.56 21.72 3.74 ;
      RECT 22.96 2.569 22.97 2.745 ;
      RECT 22.915 2.536 22.96 2.745 ;
      RECT 22.87 2.487 22.915 2.745 ;
      RECT 22.84 2.457 22.87 2.746 ;
      RECT 22.835 2.44 22.84 2.747 ;
      RECT 22.81 2.42 22.835 2.748 ;
      RECT 22.795 2.395 22.81 2.749 ;
      RECT 22.79 2.382 22.795 2.75 ;
      RECT 22.785 2.376 22.79 2.748 ;
      RECT 22.78 2.368 22.785 2.742 ;
      RECT 22.755 2.36 22.78 2.722 ;
      RECT 22.735 2.349 22.755 2.693 ;
      RECT 22.705 2.334 22.735 2.664 ;
      RECT 22.685 2.32 22.705 2.636 ;
      RECT 22.675 2.314 22.685 2.615 ;
      RECT 22.67 2.311 22.675 2.598 ;
      RECT 22.665 2.308 22.67 2.583 ;
      RECT 22.65 2.303 22.665 2.548 ;
      RECT 22.645 2.299 22.65 2.515 ;
      RECT 22.625 2.294 22.645 2.491 ;
      RECT 22.595 2.286 22.625 2.456 ;
      RECT 22.58 2.28 22.595 2.433 ;
      RECT 22.54 2.273 22.58 2.418 ;
      RECT 22.515 2.265 22.54 2.398 ;
      RECT 22.495 2.26 22.515 2.388 ;
      RECT 22.46 2.254 22.495 2.383 ;
      RECT 22.415 2.245 22.46 2.382 ;
      RECT 22.385 2.241 22.415 2.384 ;
      RECT 22.3 2.249 22.385 2.388 ;
      RECT 22.23 2.26 22.3 2.41 ;
      RECT 22.217 2.266 22.23 2.433 ;
      RECT 22.131 2.273 22.217 2.455 ;
      RECT 22.045 2.285 22.131 2.492 ;
      RECT 22.045 2.662 22.055 2.9 ;
      RECT 22.04 2.291 22.045 2.515 ;
      RECT 22.035 2.547 22.045 2.9 ;
      RECT 22.035 2.292 22.04 2.52 ;
      RECT 22.03 2.293 22.035 2.9 ;
      RECT 22.006 2.295 22.03 2.901 ;
      RECT 21.92 2.303 22.006 2.903 ;
      RECT 21.9 2.317 21.92 2.906 ;
      RECT 21.895 2.345 21.9 2.907 ;
      RECT 21.89 2.357 21.895 2.908 ;
      RECT 21.885 2.372 21.89 2.909 ;
      RECT 21.875 2.402 21.885 2.91 ;
      RECT 21.87 2.44 21.875 2.908 ;
      RECT 21.865 2.46 21.87 2.903 ;
      RECT 21.85 2.495 21.865 2.888 ;
      RECT 21.84 2.547 21.85 2.868 ;
      RECT 21.835 2.577 21.84 2.856 ;
      RECT 21.82 2.59 21.835 2.839 ;
      RECT 21.795 2.594 21.82 2.806 ;
      RECT 21.78 2.592 21.795 2.783 ;
      RECT 21.765 2.591 21.78 2.78 ;
      RECT 21.705 2.589 21.765 2.778 ;
      RECT 21.695 2.587 21.705 2.773 ;
      RECT 21.655 2.586 21.695 2.77 ;
      RECT 21.585 2.583 21.655 2.768 ;
      RECT 21.53 2.581 21.585 2.763 ;
      RECT 21.46 2.575 21.53 2.758 ;
      RECT 21.451 2.575 21.46 2.755 ;
      RECT 21.365 2.575 21.451 2.75 ;
      RECT 21.36 2.575 21.365 2.745 ;
      RECT 22.665 1.81 22.84 2.16 ;
      RECT 22.665 1.825 22.85 2.158 ;
      RECT 22.64 1.775 22.785 2.155 ;
      RECT 22.62 1.776 22.785 2.148 ;
      RECT 22.61 1.777 22.795 2.143 ;
      RECT 22.58 1.778 22.795 2.13 ;
      RECT 22.53 1.779 22.795 2.106 ;
      RECT 22.525 1.781 22.795 2.091 ;
      RECT 22.525 1.847 22.855 2.085 ;
      RECT 22.505 1.788 22.81 2.065 ;
      RECT 22.495 1.797 22.82 1.92 ;
      RECT 22.505 1.792 22.82 2.065 ;
      RECT 22.525 1.782 22.81 2.091 ;
      RECT 22.11 3.107 22.28 3.395 ;
      RECT 22.105 3.125 22.29 3.39 ;
      RECT 22.07 3.133 22.355 3.31 ;
      RECT 22.07 3.133 22.441 3.3 ;
      RECT 22.07 3.133 22.495 3.246 ;
      RECT 22.355 3.03 22.525 3.214 ;
      RECT 22.07 3.185 22.53 3.202 ;
      RECT 22.055 3.155 22.525 3.198 ;
      RECT 22.315 3.037 22.355 3.349 ;
      RECT 22.195 3.074 22.525 3.214 ;
      RECT 22.29 3.049 22.315 3.375 ;
      RECT 22.28 3.056 22.525 3.214 ;
      RECT 22.411 2.52 22.48 2.779 ;
      RECT 22.411 2.575 22.485 2.778 ;
      RECT 22.325 2.575 22.485 2.777 ;
      RECT 22.32 2.575 22.49 2.77 ;
      RECT 22.31 2.52 22.48 2.765 ;
      RECT 21.69 1.819 21.865 2.12 ;
      RECT 21.675 1.807 21.69 2.105 ;
      RECT 21.645 1.806 21.675 2.058 ;
      RECT 21.645 1.824 21.87 2.053 ;
      RECT 21.63 1.808 21.69 2.018 ;
      RECT 21.625 1.83 21.88 1.918 ;
      RECT 21.625 1.813 21.776 1.918 ;
      RECT 21.625 1.815 21.78 1.918 ;
      RECT 21.63 1.811 21.776 2.018 ;
      RECT 21.735 3.047 21.74 3.395 ;
      RECT 21.725 3.037 21.735 3.401 ;
      RECT 21.69 3.027 21.725 3.403 ;
      RECT 21.652 3.022 21.69 3.407 ;
      RECT 21.566 3.015 21.652 3.414 ;
      RECT 21.48 3.005 21.566 3.424 ;
      RECT 21.435 3 21.48 3.432 ;
      RECT 21.431 3 21.435 3.436 ;
      RECT 21.345 3 21.431 3.443 ;
      RECT 21.33 3 21.345 3.443 ;
      RECT 21.32 2.998 21.33 3.415 ;
      RECT 21.31 2.994 21.32 3.358 ;
      RECT 21.29 2.988 21.31 3.29 ;
      RECT 21.285 2.984 21.29 3.238 ;
      RECT 21.275 2.983 21.285 3.205 ;
      RECT 21.225 2.981 21.275 3.19 ;
      RECT 21.2 2.979 21.225 3.185 ;
      RECT 21.157 2.977 21.2 3.181 ;
      RECT 21.071 2.973 21.157 3.169 ;
      RECT 20.985 2.968 21.071 3.153 ;
      RECT 20.955 2.965 20.985 3.14 ;
      RECT 20.93 2.964 20.955 3.128 ;
      RECT 20.925 2.964 20.93 3.118 ;
      RECT 20.885 2.963 20.925 3.11 ;
      RECT 20.87 2.962 20.885 3.103 ;
      RECT 20.82 2.961 20.87 3.095 ;
      RECT 20.818 2.96 20.82 3.09 ;
      RECT 20.732 2.958 20.818 3.09 ;
      RECT 20.646 2.953 20.732 3.09 ;
      RECT 20.56 2.949 20.646 3.09 ;
      RECT 20.511 2.945 20.56 3.088 ;
      RECT 20.425 2.942 20.511 3.083 ;
      RECT 20.402 2.939 20.425 3.079 ;
      RECT 20.316 2.936 20.402 3.074 ;
      RECT 20.23 2.932 20.316 3.065 ;
      RECT 20.205 2.925 20.23 3.06 ;
      RECT 20.145 2.89 20.205 3.057 ;
      RECT 20.125 2.815 20.145 3.054 ;
      RECT 20.12 2.757 20.125 3.053 ;
      RECT 20.095 2.697 20.12 3.052 ;
      RECT 20.02 2.575 20.095 3.048 ;
      RECT 20.01 2.575 20.02 3.04 ;
      RECT 19.995 2.575 20.01 3.03 ;
      RECT 19.98 2.575 19.995 3 ;
      RECT 19.965 2.575 19.98 2.945 ;
      RECT 19.95 2.575 19.965 2.883 ;
      RECT 19.925 2.575 19.95 2.808 ;
      RECT 19.92 2.575 19.925 2.758 ;
      RECT 21.265 2.12 21.285 2.429 ;
      RECT 21.251 2.122 21.3 2.426 ;
      RECT 21.251 2.127 21.32 2.417 ;
      RECT 21.165 2.125 21.3 2.411 ;
      RECT 21.165 2.133 21.355 2.394 ;
      RECT 21.13 2.135 21.355 2.393 ;
      RECT 21.1 2.143 21.355 2.384 ;
      RECT 21.09 2.148 21.375 2.37 ;
      RECT 21.13 2.138 21.375 2.37 ;
      RECT 21.13 2.141 21.385 2.358 ;
      RECT 21.1 2.143 21.395 2.345 ;
      RECT 21.1 2.147 21.405 2.288 ;
      RECT 21.09 2.152 21.41 2.203 ;
      RECT 21.251 2.12 21.285 2.426 ;
      RECT 20.69 2.223 20.695 2.435 ;
      RECT 20.565 2.22 20.58 2.435 ;
      RECT 20.03 2.25 20.1 2.435 ;
      RECT 19.915 2.25 19.95 2.43 ;
      RECT 21.036 2.552 21.055 2.746 ;
      RECT 20.95 2.507 21.036 2.747 ;
      RECT 20.94 2.46 20.95 2.749 ;
      RECT 20.935 2.44 20.94 2.75 ;
      RECT 20.915 2.405 20.935 2.751 ;
      RECT 20.9 2.355 20.915 2.752 ;
      RECT 20.88 2.292 20.9 2.753 ;
      RECT 20.87 2.255 20.88 2.754 ;
      RECT 20.855 2.244 20.87 2.755 ;
      RECT 20.85 2.236 20.855 2.753 ;
      RECT 20.84 2.235 20.85 2.745 ;
      RECT 20.81 2.232 20.84 2.724 ;
      RECT 20.735 2.227 20.81 2.669 ;
      RECT 20.72 2.223 20.735 2.615 ;
      RECT 20.71 2.223 20.72 2.51 ;
      RECT 20.695 2.223 20.71 2.443 ;
      RECT 20.68 2.223 20.69 2.433 ;
      RECT 20.625 2.222 20.68 2.43 ;
      RECT 20.58 2.22 20.625 2.433 ;
      RECT 20.552 2.22 20.565 2.436 ;
      RECT 20.466 2.224 20.552 2.438 ;
      RECT 20.38 2.23 20.466 2.443 ;
      RECT 20.36 2.234 20.38 2.445 ;
      RECT 20.358 2.235 20.36 2.444 ;
      RECT 20.272 2.237 20.358 2.443 ;
      RECT 20.186 2.242 20.272 2.44 ;
      RECT 20.1 2.247 20.186 2.437 ;
      RECT 19.95 2.25 20.03 2.433 ;
      RECT 20.726 3.225 20.775 3.559 ;
      RECT 20.726 3.225 20.78 3.558 ;
      RECT 20.64 3.225 20.78 3.557 ;
      RECT 20.415 3.333 20.785 3.555 ;
      RECT 20.64 3.225 20.81 3.548 ;
      RECT 20.61 3.237 20.815 3.539 ;
      RECT 20.595 3.255 20.82 3.536 ;
      RECT 20.41 3.339 20.82 3.463 ;
      RECT 20.405 3.346 20.82 3.423 ;
      RECT 20.42 3.312 20.82 3.536 ;
      RECT 20.581 3.258 20.785 3.555 ;
      RECT 20.495 3.278 20.82 3.536 ;
      RECT 20.595 3.252 20.815 3.539 ;
      RECT 20.365 2.576 20.555 2.77 ;
      RECT 20.36 2.578 20.555 2.769 ;
      RECT 20.355 2.582 20.57 2.766 ;
      RECT 20.37 2.575 20.57 2.766 ;
      RECT 20.355 2.685 20.575 2.761 ;
      RECT 19.65 3.185 19.741 3.483 ;
      RECT 19.645 3.187 19.82 3.478 ;
      RECT 19.65 3.185 19.82 3.478 ;
      RECT 19.645 3.191 19.84 3.476 ;
      RECT 19.645 3.246 19.88 3.475 ;
      RECT 19.645 3.281 19.895 3.469 ;
      RECT 19.645 3.315 19.905 3.459 ;
      RECT 19.635 3.195 19.84 3.31 ;
      RECT 19.635 3.215 19.855 3.31 ;
      RECT 19.635 3.198 19.845 3.31 ;
      RECT 19.86 1.966 19.865 2.028 ;
      RECT 19.855 1.888 19.86 2.051 ;
      RECT 19.85 1.845 19.855 2.062 ;
      RECT 19.845 1.835 19.85 2.074 ;
      RECT 19.84 1.835 19.845 2.083 ;
      RECT 19.815 1.835 19.84 2.115 ;
      RECT 19.81 1.835 19.815 2.148 ;
      RECT 19.795 1.835 19.81 2.173 ;
      RECT 19.785 1.835 19.795 2.2 ;
      RECT 19.78 1.835 19.785 2.213 ;
      RECT 19.775 1.835 19.78 2.228 ;
      RECT 19.765 1.835 19.775 2.243 ;
      RECT 19.76 1.835 19.765 2.263 ;
      RECT 19.735 1.835 19.76 2.298 ;
      RECT 19.69 1.835 19.735 2.343 ;
      RECT 19.68 1.835 19.69 2.356 ;
      RECT 19.595 1.92 19.68 2.363 ;
      RECT 19.56 2.042 19.595 2.372 ;
      RECT 19.555 2.082 19.56 2.376 ;
      RECT 19.535 2.105 19.555 2.378 ;
      RECT 19.53 2.135 19.535 2.381 ;
      RECT 19.52 2.147 19.53 2.382 ;
      RECT 19.475 2.17 19.52 2.387 ;
      RECT 19.435 2.2 19.475 2.395 ;
      RECT 19.4 2.212 19.435 2.401 ;
      RECT 19.395 2.217 19.4 2.405 ;
      RECT 19.325 2.227 19.395 2.412 ;
      RECT 19.285 2.237 19.325 2.422 ;
      RECT 19.265 2.242 19.285 2.428 ;
      RECT 19.255 2.246 19.265 2.433 ;
      RECT 19.25 2.249 19.255 2.436 ;
      RECT 19.24 2.25 19.25 2.437 ;
      RECT 19.215 2.252 19.24 2.441 ;
      RECT 19.205 2.257 19.215 2.444 ;
      RECT 19.16 2.265 19.205 2.445 ;
      RECT 19.035 2.27 19.16 2.445 ;
      RECT 19.59 2.567 19.61 2.749 ;
      RECT 19.541 2.552 19.59 2.748 ;
      RECT 19.455 2.567 19.61 2.746 ;
      RECT 19.44 2.567 19.61 2.745 ;
      RECT 19.405 2.545 19.575 2.73 ;
      RECT 19.475 3.565 19.49 3.774 ;
      RECT 19.475 3.573 19.495 3.773 ;
      RECT 19.42 3.573 19.495 3.772 ;
      RECT 19.4 3.577 19.5 3.77 ;
      RECT 19.38 3.527 19.42 3.769 ;
      RECT 19.325 3.585 19.505 3.767 ;
      RECT 19.29 3.542 19.42 3.765 ;
      RECT 19.286 3.545 19.475 3.764 ;
      RECT 19.2 3.553 19.475 3.762 ;
      RECT 19.2 3.597 19.51 3.755 ;
      RECT 19.19 3.69 19.51 3.753 ;
      RECT 19.2 3.609 19.515 3.738 ;
      RECT 19.2 3.63 19.53 3.708 ;
      RECT 19.2 3.657 19.535 3.678 ;
      RECT 19.325 3.535 19.42 3.767 ;
      RECT 18.955 2.58 18.96 3.118 ;
      RECT 18.76 2.91 18.765 3.105 ;
      RECT 17.06 2.575 17.075 2.955 ;
      RECT 19.125 2.575 19.13 2.745 ;
      RECT 19.12 2.575 19.125 2.755 ;
      RECT 19.115 2.575 19.12 2.768 ;
      RECT 19.09 2.575 19.115 2.81 ;
      RECT 19.065 2.575 19.09 2.883 ;
      RECT 19.05 2.575 19.065 2.935 ;
      RECT 19.045 2.575 19.05 2.965 ;
      RECT 19.02 2.575 19.045 3.005 ;
      RECT 19.005 2.575 19.02 3.06 ;
      RECT 19 2.575 19.005 3.093 ;
      RECT 18.975 2.575 19 3.113 ;
      RECT 18.96 2.575 18.975 3.119 ;
      RECT 18.89 2.61 18.955 3.115 ;
      RECT 18.84 2.665 18.89 3.11 ;
      RECT 18.83 2.697 18.84 3.108 ;
      RECT 18.825 2.722 18.83 3.108 ;
      RECT 18.805 2.795 18.825 3.108 ;
      RECT 18.795 2.875 18.805 3.107 ;
      RECT 18.78 2.905 18.795 3.107 ;
      RECT 18.765 2.91 18.78 3.106 ;
      RECT 18.705 2.912 18.76 3.103 ;
      RECT 18.675 2.917 18.705 3.099 ;
      RECT 18.673 2.92 18.675 3.098 ;
      RECT 18.587 2.922 18.673 3.095 ;
      RECT 18.501 2.928 18.587 3.089 ;
      RECT 18.415 2.933 18.501 3.083 ;
      RECT 18.342 2.938 18.415 3.084 ;
      RECT 18.256 2.944 18.342 3.092 ;
      RECT 18.17 2.95 18.256 3.101 ;
      RECT 18.15 2.954 18.17 3.106 ;
      RECT 18.103 2.956 18.15 3.109 ;
      RECT 18.017 2.961 18.103 3.115 ;
      RECT 17.931 2.966 18.017 3.124 ;
      RECT 17.845 2.972 17.931 3.132 ;
      RECT 17.76 2.97 17.845 3.141 ;
      RECT 17.756 2.965 17.76 3.145 ;
      RECT 17.67 2.96 17.756 3.137 ;
      RECT 17.606 2.951 17.67 3.125 ;
      RECT 17.52 2.942 17.606 3.112 ;
      RECT 17.496 2.935 17.52 3.103 ;
      RECT 17.41 2.929 17.496 3.09 ;
      RECT 17.37 2.922 17.41 3.076 ;
      RECT 17.365 2.912 17.37 3.072 ;
      RECT 17.355 2.9 17.365 3.071 ;
      RECT 17.335 2.87 17.355 3.068 ;
      RECT 17.28 2.79 17.335 3.062 ;
      RECT 17.26 2.709 17.28 3.057 ;
      RECT 17.24 2.667 17.26 3.053 ;
      RECT 17.215 2.62 17.24 3.047 ;
      RECT 17.21 2.595 17.215 3.044 ;
      RECT 17.175 2.575 17.21 3.039 ;
      RECT 17.166 2.575 17.175 3.032 ;
      RECT 17.08 2.575 17.166 3.002 ;
      RECT 17.075 2.575 17.08 2.965 ;
      RECT 17.04 2.575 17.06 2.887 ;
      RECT 17.035 2.617 17.04 2.852 ;
      RECT 17.03 2.692 17.035 2.808 ;
      RECT 18.48 2.497 18.655 2.745 ;
      RECT 18.48 2.497 18.66 2.743 ;
      RECT 18.475 2.529 18.66 2.703 ;
      RECT 18.505 2.47 18.675 2.69 ;
      RECT 18.47 2.547 18.675 2.623 ;
      RECT 17.78 2.01 17.95 2.185 ;
      RECT 17.78 2.01 18.122 2.177 ;
      RECT 17.78 2.01 18.205 2.171 ;
      RECT 17.78 2.01 18.24 2.167 ;
      RECT 17.78 2.01 18.26 2.166 ;
      RECT 17.78 2.01 18.346 2.162 ;
      RECT 18.24 1.835 18.41 2.157 ;
      RECT 17.815 1.942 18.44 2.155 ;
      RECT 17.805 1.997 18.445 2.153 ;
      RECT 17.78 2.033 18.455 2.148 ;
      RECT 17.78 2.06 18.46 2.078 ;
      RECT 17.845 1.885 18.42 2.155 ;
      RECT 18.036 1.87 18.42 2.155 ;
      RECT 17.87 1.873 18.42 2.155 ;
      RECT 17.95 1.871 18.036 2.182 ;
      RECT 18.036 1.868 18.415 2.155 ;
      RECT 18.22 1.845 18.415 2.155 ;
      RECT 18.122 1.866 18.415 2.155 ;
      RECT 18.205 1.86 18.22 2.168 ;
      RECT 18.355 3.225 18.36 3.425 ;
      RECT 17.82 3.29 17.865 3.425 ;
      RECT 18.39 3.225 18.41 3.398 ;
      RECT 18.36 3.225 18.39 3.413 ;
      RECT 18.295 3.225 18.355 3.45 ;
      RECT 18.28 3.225 18.295 3.48 ;
      RECT 18.265 3.225 18.28 3.493 ;
      RECT 18.245 3.225 18.265 3.508 ;
      RECT 18.24 3.225 18.245 3.517 ;
      RECT 18.23 3.229 18.24 3.522 ;
      RECT 18.215 3.239 18.23 3.533 ;
      RECT 18.19 3.255 18.215 3.543 ;
      RECT 18.18 3.269 18.19 3.545 ;
      RECT 18.16 3.281 18.18 3.542 ;
      RECT 18.13 3.302 18.16 3.536 ;
      RECT 18.12 3.314 18.13 3.531 ;
      RECT 18.11 3.312 18.12 3.528 ;
      RECT 18.095 3.311 18.11 3.523 ;
      RECT 18.09 3.31 18.095 3.518 ;
      RECT 18.055 3.308 18.09 3.508 ;
      RECT 18.035 3.305 18.055 3.49 ;
      RECT 18.025 3.303 18.035 3.485 ;
      RECT 18.015 3.302 18.025 3.48 ;
      RECT 17.98 3.3 18.015 3.468 ;
      RECT 17.925 3.296 17.98 3.448 ;
      RECT 17.915 3.294 17.925 3.433 ;
      RECT 17.91 3.294 17.915 3.428 ;
      RECT 17.865 3.292 17.91 3.425 ;
      RECT 17.77 3.29 17.82 3.429 ;
      RECT 17.76 3.291 17.77 3.434 ;
      RECT 17.7 3.298 17.76 3.448 ;
      RECT 17.675 3.306 17.7 3.468 ;
      RECT 17.665 3.31 17.675 3.48 ;
      RECT 17.66 3.311 17.665 3.485 ;
      RECT 17.645 3.313 17.66 3.488 ;
      RECT 17.63 3.315 17.645 3.493 ;
      RECT 17.625 3.315 17.63 3.496 ;
      RECT 17.58 3.32 17.625 3.507 ;
      RECT 17.575 3.324 17.58 3.519 ;
      RECT 17.55 3.32 17.575 3.523 ;
      RECT 17.54 3.316 17.55 3.527 ;
      RECT 17.53 3.315 17.54 3.531 ;
      RECT 17.515 3.305 17.53 3.537 ;
      RECT 17.51 3.293 17.515 3.541 ;
      RECT 17.505 3.29 17.51 3.542 ;
      RECT 17.5 3.287 17.505 3.544 ;
      RECT 17.485 3.275 17.5 3.543 ;
      RECT 17.47 3.257 17.485 3.54 ;
      RECT 17.45 3.236 17.47 3.533 ;
      RECT 17.385 3.225 17.45 3.505 ;
      RECT 17.381 3.225 17.385 3.484 ;
      RECT 17.295 3.225 17.381 3.454 ;
      RECT 17.28 3.225 17.295 3.41 ;
      RECT 17.855 2.325 17.86 2.56 ;
      RECT 16.985 2.241 16.99 2.445 ;
      RECT 17.565 2.27 17.57 2.425 ;
      RECT 17.485 2.25 17.49 2.425 ;
      RECT 18.155 2.392 18.17 2.745 ;
      RECT 18.081 2.377 18.155 2.745 ;
      RECT 17.995 2.36 18.081 2.745 ;
      RECT 17.985 2.35 17.995 2.743 ;
      RECT 17.98 2.348 17.985 2.738 ;
      RECT 17.965 2.346 17.98 2.724 ;
      RECT 17.895 2.338 17.965 2.664 ;
      RECT 17.875 2.329 17.895 2.598 ;
      RECT 17.87 2.326 17.875 2.578 ;
      RECT 17.86 2.325 17.87 2.568 ;
      RECT 17.85 2.325 17.855 2.552 ;
      RECT 17.84 2.324 17.85 2.542 ;
      RECT 17.83 2.322 17.84 2.53 ;
      RECT 17.815 2.319 17.83 2.51 ;
      RECT 17.805 2.317 17.815 2.495 ;
      RECT 17.785 2.314 17.805 2.483 ;
      RECT 17.78 2.312 17.785 2.473 ;
      RECT 17.755 2.31 17.78 2.46 ;
      RECT 17.725 2.305 17.755 2.445 ;
      RECT 17.645 2.296 17.725 2.436 ;
      RECT 17.6 2.285 17.645 2.429 ;
      RECT 17.58 2.276 17.6 2.426 ;
      RECT 17.57 2.271 17.58 2.425 ;
      RECT 17.525 2.265 17.565 2.425 ;
      RECT 17.51 2.257 17.525 2.425 ;
      RECT 17.49 2.252 17.51 2.425 ;
      RECT 17.47 2.249 17.485 2.425 ;
      RECT 17.387 2.248 17.47 2.424 ;
      RECT 17.301 2.247 17.387 2.42 ;
      RECT 17.215 2.245 17.301 2.417 ;
      RECT 17.162 2.244 17.215 2.419 ;
      RECT 17.076 2.243 17.162 2.428 ;
      RECT 16.99 2.242 17.076 2.44 ;
      RECT 16.97 2.241 16.985 2.448 ;
      RECT 16.89 2.24 16.97 2.46 ;
      RECT 16.865 2.24 16.89 2.473 ;
      RECT 16.84 2.24 16.865 2.488 ;
      RECT 16.835 2.24 16.84 2.51 ;
      RECT 16.83 2.24 16.835 2.528 ;
      RECT 16.825 2.24 16.83 2.545 ;
      RECT 16.82 2.24 16.825 2.558 ;
      RECT 16.815 2.24 16.82 2.568 ;
      RECT 16.775 2.24 16.815 2.653 ;
      RECT 16.76 2.24 16.775 2.738 ;
      RECT 16.75 2.241 16.76 2.75 ;
      RECT 16.715 2.246 16.75 2.755 ;
      RECT 16.675 2.255 16.715 2.755 ;
      RECT 16.66 2.265 16.675 2.755 ;
      RECT 16.655 2.275 16.66 2.755 ;
      RECT 16.635 2.302 16.655 2.755 ;
      RECT 16.585 2.385 16.635 2.755 ;
      RECT 16.58 2.447 16.585 2.755 ;
      RECT 16.57 2.46 16.58 2.755 ;
      RECT 16.56 2.482 16.57 2.755 ;
      RECT 16.55 2.507 16.56 2.75 ;
      RECT 16.545 2.545 16.55 2.743 ;
      RECT 16.535 2.655 16.545 2.738 ;
      RECT 17.93 3.576 17.945 3.835 ;
      RECT 17.93 3.591 17.95 3.834 ;
      RECT 17.846 3.591 17.95 3.832 ;
      RECT 17.846 3.605 17.955 3.831 ;
      RECT 17.76 3.647 17.96 3.828 ;
      RECT 17.755 3.59 17.945 3.823 ;
      RECT 17.755 3.661 17.965 3.82 ;
      RECT 17.75 3.692 17.965 3.818 ;
      RECT 17.755 3.689 17.98 3.808 ;
      RECT 17.75 3.735 17.995 3.793 ;
      RECT 17.75 3.763 18 3.778 ;
      RECT 17.76 3.565 17.93 3.828 ;
      RECT 17.52 2.575 17.69 2.745 ;
      RECT 17.485 2.575 17.69 2.74 ;
      RECT 17.475 2.575 17.69 2.733 ;
      RECT 17.47 2.56 17.64 2.73 ;
      RECT 16.3 3.097 16.565 3.54 ;
      RECT 16.295 3.068 16.51 3.538 ;
      RECT 16.29 3.222 16.57 3.533 ;
      RECT 16.295 3.117 16.57 3.533 ;
      RECT 16.295 3.128 16.58 3.52 ;
      RECT 16.295 3.075 16.54 3.538 ;
      RECT 16.3 3.062 16.51 3.54 ;
      RECT 16.3 3.06 16.46 3.54 ;
      RECT 16.401 3.052 16.46 3.54 ;
      RECT 16.315 3.053 16.46 3.54 ;
      RECT 16.401 3.051 16.45 3.54 ;
      RECT 16.205 1.866 16.38 2.165 ;
      RECT 16.255 1.828 16.38 2.165 ;
      RECT 16.24 1.83 16.466 2.157 ;
      RECT 16.24 1.833 16.505 2.144 ;
      RECT 16.24 1.834 16.515 2.13 ;
      RECT 16.195 1.885 16.515 2.12 ;
      RECT 16.24 1.835 16.52 2.115 ;
      RECT 16.195 2.045 16.525 2.105 ;
      RECT 16.18 1.905 16.52 2.045 ;
      RECT 16.175 1.921 16.52 1.985 ;
      RECT 16.22 1.845 16.52 2.115 ;
      RECT 16.255 1.826 16.341 2.165 ;
      RECT 14.35 1.74 14.52 2.935 ;
      RECT 14.35 1.74 14.815 1.91 ;
      RECT 14.35 6.97 14.815 7.14 ;
      RECT 14.35 5.945 14.52 7.14 ;
      RECT 13.36 1.74 13.53 2.935 ;
      RECT 13.36 1.74 13.825 1.91 ;
      RECT 13.36 6.97 13.825 7.14 ;
      RECT 13.36 5.945 13.53 7.14 ;
      RECT 11.505 2.635 11.675 3.865 ;
      RECT 11.56 0.855 11.73 2.805 ;
      RECT 11.505 0.575 11.675 1.025 ;
      RECT 11.505 7.855 11.675 8.305 ;
      RECT 11.56 6.075 11.73 8.025 ;
      RECT 11.505 5.015 11.675 6.245 ;
      RECT 10.985 0.575 11.155 3.865 ;
      RECT 10.985 2.075 11.39 2.405 ;
      RECT 10.985 1.235 11.39 1.565 ;
      RECT 10.985 5.015 11.155 8.305 ;
      RECT 10.985 7.315 11.39 7.645 ;
      RECT 10.985 6.475 11.39 6.805 ;
      RECT 8.91 3.126 8.915 3.298 ;
      RECT 8.905 3.119 8.91 3.388 ;
      RECT 8.9 3.113 8.905 3.407 ;
      RECT 8.88 3.107 8.9 3.417 ;
      RECT 8.865 3.102 8.88 3.425 ;
      RECT 8.828 3.096 8.865 3.423 ;
      RECT 8.742 3.082 8.828 3.419 ;
      RECT 8.656 3.064 8.742 3.414 ;
      RECT 8.57 3.045 8.656 3.408 ;
      RECT 8.54 3.033 8.57 3.404 ;
      RECT 8.52 3.027 8.54 3.403 ;
      RECT 8.455 3.025 8.52 3.401 ;
      RECT 8.44 3.025 8.455 3.393 ;
      RECT 8.425 3.025 8.44 3.38 ;
      RECT 8.42 3.025 8.425 3.37 ;
      RECT 8.405 3.025 8.42 3.348 ;
      RECT 8.39 3.025 8.405 3.315 ;
      RECT 8.385 3.025 8.39 3.293 ;
      RECT 8.375 3.025 8.385 3.275 ;
      RECT 8.36 3.025 8.375 3.253 ;
      RECT 8.34 3.025 8.36 3.215 ;
      RECT 8.69 2.31 8.725 2.749 ;
      RECT 8.69 2.31 8.73 2.748 ;
      RECT 8.635 2.37 8.73 2.747 ;
      RECT 8.5 2.542 8.73 2.746 ;
      RECT 8.61 2.42 8.73 2.746 ;
      RECT 8.5 2.542 8.755 2.736 ;
      RECT 8.555 2.487 8.835 2.653 ;
      RECT 8.73 2.281 8.735 2.744 ;
      RECT 8.585 2.457 8.875 2.53 ;
      RECT 8.6 2.44 8.73 2.746 ;
      RECT 8.735 2.28 8.905 2.468 ;
      RECT 8.725 2.283 8.905 2.468 ;
      RECT 8.23 2.16 8.4 2.47 ;
      RECT 8.23 2.16 8.405 2.443 ;
      RECT 8.23 2.16 8.41 2.42 ;
      RECT 8.23 2.16 8.42 2.37 ;
      RECT 8.225 2.265 8.42 2.34 ;
      RECT 8.26 1.835 8.43 2.313 ;
      RECT 8.26 1.835 8.445 2.234 ;
      RECT 8.25 2.045 8.445 2.234 ;
      RECT 8.26 1.845 8.455 2.149 ;
      RECT 8.19 2.587 8.195 2.79 ;
      RECT 8.18 2.575 8.19 2.9 ;
      RECT 8.155 2.575 8.18 2.94 ;
      RECT 8.075 2.575 8.155 3.025 ;
      RECT 8.065 2.575 8.075 3.095 ;
      RECT 8.04 2.575 8.065 3.118 ;
      RECT 8.02 2.575 8.04 3.153 ;
      RECT 7.975 2.585 8.02 3.196 ;
      RECT 7.965 2.597 7.975 3.233 ;
      RECT 7.945 2.611 7.965 3.253 ;
      RECT 7.935 2.629 7.945 3.269 ;
      RECT 7.92 2.655 7.935 3.279 ;
      RECT 7.905 2.696 7.92 3.293 ;
      RECT 7.895 2.731 7.905 3.303 ;
      RECT 7.89 2.747 7.895 3.308 ;
      RECT 7.88 2.762 7.89 3.313 ;
      RECT 7.86 2.805 7.88 3.323 ;
      RECT 7.84 2.842 7.86 3.336 ;
      RECT 7.805 2.865 7.84 3.354 ;
      RECT 7.795 2.879 7.805 3.37 ;
      RECT 7.775 2.889 7.795 3.38 ;
      RECT 7.77 2.898 7.775 3.388 ;
      RECT 7.76 2.905 7.77 3.395 ;
      RECT 7.75 2.912 7.76 3.403 ;
      RECT 7.735 2.922 7.75 3.411 ;
      RECT 7.725 2.936 7.735 3.421 ;
      RECT 7.715 2.948 7.725 3.433 ;
      RECT 7.7 2.97 7.715 3.446 ;
      RECT 7.69 2.992 7.7 3.457 ;
      RECT 7.68 3.012 7.69 3.466 ;
      RECT 7.675 3.027 7.68 3.473 ;
      RECT 7.645 3.06 7.675 3.487 ;
      RECT 7.635 3.095 7.645 3.502 ;
      RECT 7.63 3.102 7.635 3.508 ;
      RECT 7.61 3.117 7.63 3.515 ;
      RECT 7.605 3.132 7.61 3.523 ;
      RECT 7.6 3.141 7.605 3.528 ;
      RECT 7.585 3.147 7.6 3.535 ;
      RECT 7.58 3.153 7.585 3.543 ;
      RECT 7.575 3.157 7.58 3.55 ;
      RECT 7.57 3.161 7.575 3.56 ;
      RECT 7.56 3.166 7.57 3.57 ;
      RECT 7.54 3.177 7.56 3.598 ;
      RECT 7.525 3.189 7.54 3.625 ;
      RECT 7.505 3.202 7.525 3.65 ;
      RECT 7.485 3.217 7.505 3.674 ;
      RECT 7.47 3.232 7.485 3.689 ;
      RECT 7.465 3.243 7.47 3.698 ;
      RECT 7.4 3.288 7.465 3.708 ;
      RECT 7.365 3.347 7.4 3.721 ;
      RECT 7.36 3.37 7.365 3.727 ;
      RECT 7.355 3.377 7.36 3.729 ;
      RECT 7.34 3.387 7.355 3.732 ;
      RECT 7.31 3.412 7.34 3.736 ;
      RECT 7.305 3.43 7.31 3.74 ;
      RECT 7.3 3.437 7.305 3.741 ;
      RECT 7.28 3.445 7.3 3.745 ;
      RECT 7.27 3.452 7.28 3.749 ;
      RECT 7.226 3.463 7.27 3.756 ;
      RECT 7.14 3.491 7.226 3.772 ;
      RECT 7.08 3.515 7.14 3.79 ;
      RECT 7.035 3.525 7.08 3.804 ;
      RECT 6.976 3.533 7.035 3.818 ;
      RECT 6.89 3.54 6.976 3.837 ;
      RECT 6.865 3.545 6.89 3.852 ;
      RECT 6.785 3.548 6.865 3.855 ;
      RECT 6.705 3.552 6.785 3.842 ;
      RECT 6.696 3.555 6.705 3.827 ;
      RECT 6.61 3.555 6.696 3.812 ;
      RECT 6.55 3.557 6.61 3.789 ;
      RECT 6.546 3.56 6.55 3.779 ;
      RECT 6.46 3.56 6.546 3.764 ;
      RECT 6.385 3.56 6.46 3.74 ;
      RECT 7.7 2.569 7.71 2.745 ;
      RECT 7.655 2.536 7.7 2.745 ;
      RECT 7.61 2.487 7.655 2.745 ;
      RECT 7.58 2.457 7.61 2.746 ;
      RECT 7.575 2.44 7.58 2.747 ;
      RECT 7.55 2.42 7.575 2.748 ;
      RECT 7.535 2.395 7.55 2.749 ;
      RECT 7.53 2.382 7.535 2.75 ;
      RECT 7.525 2.376 7.53 2.748 ;
      RECT 7.52 2.368 7.525 2.742 ;
      RECT 7.495 2.36 7.52 2.722 ;
      RECT 7.475 2.349 7.495 2.693 ;
      RECT 7.445 2.334 7.475 2.664 ;
      RECT 7.425 2.32 7.445 2.636 ;
      RECT 7.415 2.314 7.425 2.615 ;
      RECT 7.41 2.311 7.415 2.598 ;
      RECT 7.405 2.308 7.41 2.583 ;
      RECT 7.39 2.303 7.405 2.548 ;
      RECT 7.385 2.299 7.39 2.515 ;
      RECT 7.365 2.294 7.385 2.491 ;
      RECT 7.335 2.286 7.365 2.456 ;
      RECT 7.32 2.28 7.335 2.433 ;
      RECT 7.28 2.273 7.32 2.418 ;
      RECT 7.255 2.265 7.28 2.398 ;
      RECT 7.235 2.26 7.255 2.388 ;
      RECT 7.2 2.254 7.235 2.383 ;
      RECT 7.155 2.245 7.2 2.382 ;
      RECT 7.125 2.241 7.155 2.384 ;
      RECT 7.04 2.249 7.125 2.388 ;
      RECT 6.97 2.26 7.04 2.41 ;
      RECT 6.957 2.266 6.97 2.433 ;
      RECT 6.871 2.273 6.957 2.455 ;
      RECT 6.785 2.285 6.871 2.492 ;
      RECT 6.785 2.662 6.795 2.9 ;
      RECT 6.78 2.291 6.785 2.515 ;
      RECT 6.775 2.547 6.785 2.9 ;
      RECT 6.775 2.292 6.78 2.52 ;
      RECT 6.77 2.293 6.775 2.9 ;
      RECT 6.746 2.295 6.77 2.901 ;
      RECT 6.66 2.303 6.746 2.903 ;
      RECT 6.64 2.317 6.66 2.906 ;
      RECT 6.635 2.345 6.64 2.907 ;
      RECT 6.63 2.357 6.635 2.908 ;
      RECT 6.625 2.372 6.63 2.909 ;
      RECT 6.615 2.402 6.625 2.91 ;
      RECT 6.61 2.44 6.615 2.908 ;
      RECT 6.605 2.46 6.61 2.903 ;
      RECT 6.59 2.495 6.605 2.888 ;
      RECT 6.58 2.547 6.59 2.868 ;
      RECT 6.575 2.577 6.58 2.856 ;
      RECT 6.56 2.59 6.575 2.839 ;
      RECT 6.535 2.594 6.56 2.806 ;
      RECT 6.52 2.592 6.535 2.783 ;
      RECT 6.505 2.591 6.52 2.78 ;
      RECT 6.445 2.589 6.505 2.778 ;
      RECT 6.435 2.587 6.445 2.773 ;
      RECT 6.395 2.586 6.435 2.77 ;
      RECT 6.325 2.583 6.395 2.768 ;
      RECT 6.27 2.581 6.325 2.763 ;
      RECT 6.2 2.575 6.27 2.758 ;
      RECT 6.191 2.575 6.2 2.755 ;
      RECT 6.105 2.575 6.191 2.75 ;
      RECT 6.1 2.575 6.105 2.745 ;
      RECT 7.405 1.81 7.58 2.16 ;
      RECT 7.405 1.825 7.59 2.158 ;
      RECT 7.38 1.775 7.525 2.155 ;
      RECT 7.36 1.776 7.525 2.148 ;
      RECT 7.35 1.777 7.535 2.143 ;
      RECT 7.32 1.778 7.535 2.13 ;
      RECT 7.27 1.779 7.535 2.106 ;
      RECT 7.265 1.781 7.535 2.091 ;
      RECT 7.265 1.847 7.595 2.085 ;
      RECT 7.245 1.788 7.55 2.065 ;
      RECT 7.235 1.797 7.56 1.92 ;
      RECT 7.245 1.792 7.56 2.065 ;
      RECT 7.265 1.782 7.55 2.091 ;
      RECT 6.85 3.107 7.02 3.395 ;
      RECT 6.845 3.125 7.03 3.39 ;
      RECT 6.81 3.133 7.095 3.31 ;
      RECT 6.81 3.133 7.181 3.3 ;
      RECT 6.81 3.133 7.235 3.246 ;
      RECT 7.095 3.03 7.265 3.214 ;
      RECT 6.81 3.185 7.27 3.202 ;
      RECT 6.795 3.155 7.265 3.198 ;
      RECT 7.055 3.037 7.095 3.349 ;
      RECT 6.935 3.074 7.265 3.214 ;
      RECT 7.03 3.049 7.055 3.375 ;
      RECT 7.02 3.056 7.265 3.214 ;
      RECT 7.151 2.52 7.22 2.779 ;
      RECT 7.151 2.575 7.225 2.778 ;
      RECT 7.065 2.575 7.225 2.777 ;
      RECT 7.06 2.575 7.23 2.77 ;
      RECT 7.05 2.52 7.22 2.765 ;
      RECT 6.43 1.819 6.605 2.12 ;
      RECT 6.415 1.807 6.43 2.105 ;
      RECT 6.385 1.806 6.415 2.058 ;
      RECT 6.385 1.824 6.61 2.053 ;
      RECT 6.37 1.808 6.43 2.018 ;
      RECT 6.365 1.83 6.62 1.918 ;
      RECT 6.365 1.813 6.516 1.918 ;
      RECT 6.365 1.815 6.52 1.918 ;
      RECT 6.37 1.811 6.516 2.018 ;
      RECT 6.475 3.047 6.48 3.395 ;
      RECT 6.465 3.037 6.475 3.401 ;
      RECT 6.43 3.027 6.465 3.403 ;
      RECT 6.392 3.022 6.43 3.407 ;
      RECT 6.306 3.015 6.392 3.414 ;
      RECT 6.22 3.005 6.306 3.424 ;
      RECT 6.175 3 6.22 3.432 ;
      RECT 6.171 3 6.175 3.436 ;
      RECT 6.085 3 6.171 3.443 ;
      RECT 6.07 3 6.085 3.443 ;
      RECT 6.06 2.998 6.07 3.415 ;
      RECT 6.05 2.994 6.06 3.358 ;
      RECT 6.03 2.988 6.05 3.29 ;
      RECT 6.025 2.984 6.03 3.238 ;
      RECT 6.015 2.983 6.025 3.205 ;
      RECT 5.965 2.981 6.015 3.19 ;
      RECT 5.94 2.979 5.965 3.185 ;
      RECT 5.897 2.977 5.94 3.181 ;
      RECT 5.811 2.973 5.897 3.169 ;
      RECT 5.725 2.968 5.811 3.153 ;
      RECT 5.695 2.965 5.725 3.14 ;
      RECT 5.67 2.964 5.695 3.128 ;
      RECT 5.665 2.964 5.67 3.118 ;
      RECT 5.625 2.963 5.665 3.11 ;
      RECT 5.61 2.962 5.625 3.103 ;
      RECT 5.56 2.961 5.61 3.095 ;
      RECT 5.558 2.96 5.56 3.09 ;
      RECT 5.472 2.958 5.558 3.09 ;
      RECT 5.386 2.953 5.472 3.09 ;
      RECT 5.3 2.949 5.386 3.09 ;
      RECT 5.251 2.945 5.3 3.088 ;
      RECT 5.165 2.942 5.251 3.083 ;
      RECT 5.142 2.939 5.165 3.079 ;
      RECT 5.056 2.936 5.142 3.074 ;
      RECT 4.97 2.932 5.056 3.065 ;
      RECT 4.945 2.925 4.97 3.06 ;
      RECT 4.885 2.89 4.945 3.057 ;
      RECT 4.865 2.815 4.885 3.054 ;
      RECT 4.86 2.757 4.865 3.053 ;
      RECT 4.835 2.697 4.86 3.052 ;
      RECT 4.76 2.575 4.835 3.048 ;
      RECT 4.75 2.575 4.76 3.04 ;
      RECT 4.735 2.575 4.75 3.03 ;
      RECT 4.72 2.575 4.735 3 ;
      RECT 4.705 2.575 4.72 2.945 ;
      RECT 4.69 2.575 4.705 2.883 ;
      RECT 4.665 2.575 4.69 2.808 ;
      RECT 4.66 2.575 4.665 2.758 ;
      RECT 6.005 2.12 6.025 2.429 ;
      RECT 5.991 2.122 6.04 2.426 ;
      RECT 5.991 2.127 6.06 2.417 ;
      RECT 5.905 2.125 6.04 2.411 ;
      RECT 5.905 2.133 6.095 2.394 ;
      RECT 5.87 2.135 6.095 2.393 ;
      RECT 5.84 2.143 6.095 2.384 ;
      RECT 5.83 2.148 6.115 2.37 ;
      RECT 5.87 2.138 6.115 2.37 ;
      RECT 5.87 2.141 6.125 2.358 ;
      RECT 5.84 2.143 6.135 2.345 ;
      RECT 5.84 2.147 6.145 2.288 ;
      RECT 5.83 2.152 6.15 2.203 ;
      RECT 5.991 2.12 6.025 2.426 ;
      RECT 5.43 2.223 5.435 2.435 ;
      RECT 5.305 2.22 5.32 2.435 ;
      RECT 4.77 2.25 4.84 2.435 ;
      RECT 4.655 2.25 4.69 2.43 ;
      RECT 5.776 2.552 5.795 2.746 ;
      RECT 5.69 2.507 5.776 2.747 ;
      RECT 5.68 2.46 5.69 2.749 ;
      RECT 5.675 2.44 5.68 2.75 ;
      RECT 5.655 2.405 5.675 2.751 ;
      RECT 5.64 2.355 5.655 2.752 ;
      RECT 5.62 2.292 5.64 2.753 ;
      RECT 5.61 2.255 5.62 2.754 ;
      RECT 5.595 2.244 5.61 2.755 ;
      RECT 5.59 2.236 5.595 2.753 ;
      RECT 5.58 2.235 5.59 2.745 ;
      RECT 5.55 2.232 5.58 2.724 ;
      RECT 5.475 2.227 5.55 2.669 ;
      RECT 5.46 2.223 5.475 2.615 ;
      RECT 5.45 2.223 5.46 2.51 ;
      RECT 5.435 2.223 5.45 2.443 ;
      RECT 5.42 2.223 5.43 2.433 ;
      RECT 5.365 2.222 5.42 2.43 ;
      RECT 5.32 2.22 5.365 2.433 ;
      RECT 5.292 2.22 5.305 2.436 ;
      RECT 5.206 2.224 5.292 2.438 ;
      RECT 5.12 2.23 5.206 2.443 ;
      RECT 5.1 2.234 5.12 2.445 ;
      RECT 5.098 2.235 5.1 2.444 ;
      RECT 5.012 2.237 5.098 2.443 ;
      RECT 4.926 2.242 5.012 2.44 ;
      RECT 4.84 2.247 4.926 2.437 ;
      RECT 4.69 2.25 4.77 2.433 ;
      RECT 5.466 3.225 5.515 3.559 ;
      RECT 5.466 3.225 5.52 3.558 ;
      RECT 5.38 3.225 5.52 3.557 ;
      RECT 5.155 3.333 5.525 3.555 ;
      RECT 5.38 3.225 5.55 3.548 ;
      RECT 5.35 3.237 5.555 3.539 ;
      RECT 5.335 3.255 5.56 3.536 ;
      RECT 5.15 3.339 5.56 3.463 ;
      RECT 5.145 3.346 5.56 3.423 ;
      RECT 5.16 3.312 5.56 3.536 ;
      RECT 5.321 3.258 5.525 3.555 ;
      RECT 5.235 3.278 5.56 3.536 ;
      RECT 5.335 3.252 5.555 3.539 ;
      RECT 5.105 2.576 5.295 2.77 ;
      RECT 5.1 2.578 5.295 2.769 ;
      RECT 5.095 2.582 5.31 2.766 ;
      RECT 5.11 2.575 5.31 2.766 ;
      RECT 5.095 2.685 5.315 2.761 ;
      RECT 4.39 3.185 4.481 3.483 ;
      RECT 4.385 3.187 4.56 3.478 ;
      RECT 4.39 3.185 4.56 3.478 ;
      RECT 4.385 3.191 4.58 3.476 ;
      RECT 4.385 3.246 4.62 3.475 ;
      RECT 4.385 3.281 4.635 3.469 ;
      RECT 4.385 3.315 4.645 3.459 ;
      RECT 4.375 3.195 4.58 3.31 ;
      RECT 4.375 3.215 4.595 3.31 ;
      RECT 4.375 3.198 4.585 3.31 ;
      RECT 4.6 1.966 4.605 2.028 ;
      RECT 4.595 1.888 4.6 2.051 ;
      RECT 4.59 1.845 4.595 2.062 ;
      RECT 4.585 1.835 4.59 2.074 ;
      RECT 4.58 1.835 4.585 2.083 ;
      RECT 4.555 1.835 4.58 2.115 ;
      RECT 4.55 1.835 4.555 2.148 ;
      RECT 4.535 1.835 4.55 2.173 ;
      RECT 4.525 1.835 4.535 2.2 ;
      RECT 4.52 1.835 4.525 2.213 ;
      RECT 4.515 1.835 4.52 2.228 ;
      RECT 4.505 1.835 4.515 2.243 ;
      RECT 4.5 1.835 4.505 2.263 ;
      RECT 4.475 1.835 4.5 2.298 ;
      RECT 4.43 1.835 4.475 2.343 ;
      RECT 4.42 1.835 4.43 2.356 ;
      RECT 4.335 1.92 4.42 2.363 ;
      RECT 4.3 2.042 4.335 2.372 ;
      RECT 4.295 2.082 4.3 2.376 ;
      RECT 4.275 2.105 4.295 2.378 ;
      RECT 4.27 2.135 4.275 2.381 ;
      RECT 4.26 2.147 4.27 2.382 ;
      RECT 4.215 2.17 4.26 2.387 ;
      RECT 4.175 2.2 4.215 2.395 ;
      RECT 4.14 2.212 4.175 2.401 ;
      RECT 4.135 2.217 4.14 2.405 ;
      RECT 4.065 2.227 4.135 2.412 ;
      RECT 4.025 2.237 4.065 2.422 ;
      RECT 4.005 2.242 4.025 2.428 ;
      RECT 3.995 2.246 4.005 2.433 ;
      RECT 3.99 2.249 3.995 2.436 ;
      RECT 3.98 2.25 3.99 2.437 ;
      RECT 3.955 2.252 3.98 2.441 ;
      RECT 3.945 2.257 3.955 2.444 ;
      RECT 3.9 2.265 3.945 2.445 ;
      RECT 3.775 2.27 3.9 2.445 ;
      RECT 4.33 2.567 4.35 2.749 ;
      RECT 4.281 2.552 4.33 2.748 ;
      RECT 4.195 2.567 4.35 2.746 ;
      RECT 4.18 2.567 4.35 2.745 ;
      RECT 4.145 2.545 4.315 2.73 ;
      RECT 4.215 3.565 4.23 3.774 ;
      RECT 4.215 3.573 4.235 3.773 ;
      RECT 4.16 3.573 4.235 3.772 ;
      RECT 4.14 3.577 4.24 3.77 ;
      RECT 4.12 3.527 4.16 3.769 ;
      RECT 4.065 3.585 4.245 3.767 ;
      RECT 4.03 3.542 4.16 3.765 ;
      RECT 4.026 3.545 4.215 3.764 ;
      RECT 3.94 3.553 4.215 3.762 ;
      RECT 3.94 3.597 4.25 3.755 ;
      RECT 3.93 3.69 4.25 3.753 ;
      RECT 3.94 3.609 4.255 3.738 ;
      RECT 3.94 3.63 4.27 3.708 ;
      RECT 3.94 3.657 4.275 3.678 ;
      RECT 4.065 3.535 4.16 3.767 ;
      RECT 3.695 2.58 3.7 3.118 ;
      RECT 3.5 2.91 3.505 3.105 ;
      RECT 1.8 2.575 1.815 2.955 ;
      RECT 3.865 2.575 3.87 2.745 ;
      RECT 3.86 2.575 3.865 2.755 ;
      RECT 3.855 2.575 3.86 2.768 ;
      RECT 3.83 2.575 3.855 2.81 ;
      RECT 3.805 2.575 3.83 2.883 ;
      RECT 3.79 2.575 3.805 2.935 ;
      RECT 3.785 2.575 3.79 2.965 ;
      RECT 3.76 2.575 3.785 3.005 ;
      RECT 3.745 2.575 3.76 3.06 ;
      RECT 3.74 2.575 3.745 3.093 ;
      RECT 3.715 2.575 3.74 3.113 ;
      RECT 3.7 2.575 3.715 3.119 ;
      RECT 3.63 2.61 3.695 3.115 ;
      RECT 3.58 2.665 3.63 3.11 ;
      RECT 3.57 2.697 3.58 3.108 ;
      RECT 3.565 2.722 3.57 3.108 ;
      RECT 3.545 2.795 3.565 3.108 ;
      RECT 3.535 2.875 3.545 3.107 ;
      RECT 3.52 2.905 3.535 3.107 ;
      RECT 3.505 2.91 3.52 3.106 ;
      RECT 3.445 2.912 3.5 3.103 ;
      RECT 3.415 2.917 3.445 3.099 ;
      RECT 3.413 2.92 3.415 3.098 ;
      RECT 3.327 2.922 3.413 3.095 ;
      RECT 3.241 2.928 3.327 3.089 ;
      RECT 3.155 2.933 3.241 3.083 ;
      RECT 3.082 2.938 3.155 3.084 ;
      RECT 2.996 2.944 3.082 3.092 ;
      RECT 2.91 2.95 2.996 3.101 ;
      RECT 2.89 2.954 2.91 3.106 ;
      RECT 2.843 2.956 2.89 3.109 ;
      RECT 2.757 2.961 2.843 3.115 ;
      RECT 2.671 2.966 2.757 3.124 ;
      RECT 2.585 2.972 2.671 3.132 ;
      RECT 2.5 2.97 2.585 3.141 ;
      RECT 2.496 2.965 2.5 3.145 ;
      RECT 2.41 2.96 2.496 3.137 ;
      RECT 2.346 2.951 2.41 3.125 ;
      RECT 2.26 2.942 2.346 3.112 ;
      RECT 2.236 2.935 2.26 3.103 ;
      RECT 2.15 2.929 2.236 3.09 ;
      RECT 2.11 2.922 2.15 3.076 ;
      RECT 2.105 2.912 2.11 3.072 ;
      RECT 2.095 2.9 2.105 3.071 ;
      RECT 2.075 2.87 2.095 3.068 ;
      RECT 2.02 2.79 2.075 3.062 ;
      RECT 2 2.709 2.02 3.057 ;
      RECT 1.98 2.667 2 3.053 ;
      RECT 1.955 2.62 1.98 3.047 ;
      RECT 1.95 2.595 1.955 3.044 ;
      RECT 1.915 2.575 1.95 3.039 ;
      RECT 1.906 2.575 1.915 3.032 ;
      RECT 1.82 2.575 1.906 3.002 ;
      RECT 1.815 2.575 1.82 2.965 ;
      RECT 1.78 2.575 1.8 2.887 ;
      RECT 1.775 2.617 1.78 2.852 ;
      RECT 1.77 2.692 1.775 2.808 ;
      RECT 3.22 2.497 3.395 2.745 ;
      RECT 3.22 2.497 3.4 2.743 ;
      RECT 3.215 2.529 3.4 2.703 ;
      RECT 3.245 2.47 3.415 2.69 ;
      RECT 3.21 2.547 3.415 2.623 ;
      RECT 2.52 2.01 2.69 2.185 ;
      RECT 2.52 2.01 2.862 2.177 ;
      RECT 2.52 2.01 2.945 2.171 ;
      RECT 2.52 2.01 2.98 2.167 ;
      RECT 2.52 2.01 3 2.166 ;
      RECT 2.52 2.01 3.086 2.162 ;
      RECT 2.98 1.835 3.15 2.157 ;
      RECT 2.555 1.942 3.18 2.155 ;
      RECT 2.545 1.997 3.185 2.153 ;
      RECT 2.52 2.033 3.195 2.148 ;
      RECT 2.52 2.06 3.2 2.078 ;
      RECT 2.585 1.885 3.16 2.155 ;
      RECT 2.776 1.87 3.16 2.155 ;
      RECT 2.61 1.873 3.16 2.155 ;
      RECT 2.69 1.871 2.776 2.182 ;
      RECT 2.776 1.868 3.155 2.155 ;
      RECT 2.96 1.845 3.155 2.155 ;
      RECT 2.862 1.866 3.155 2.155 ;
      RECT 2.945 1.86 2.96 2.168 ;
      RECT 3.095 3.225 3.1 3.425 ;
      RECT 2.56 3.29 2.605 3.425 ;
      RECT 3.13 3.225 3.15 3.398 ;
      RECT 3.1 3.225 3.13 3.413 ;
      RECT 3.035 3.225 3.095 3.45 ;
      RECT 3.02 3.225 3.035 3.48 ;
      RECT 3.005 3.225 3.02 3.493 ;
      RECT 2.985 3.225 3.005 3.508 ;
      RECT 2.98 3.225 2.985 3.517 ;
      RECT 2.97 3.229 2.98 3.522 ;
      RECT 2.955 3.239 2.97 3.533 ;
      RECT 2.93 3.255 2.955 3.543 ;
      RECT 2.92 3.269 2.93 3.545 ;
      RECT 2.9 3.281 2.92 3.542 ;
      RECT 2.87 3.302 2.9 3.536 ;
      RECT 2.86 3.314 2.87 3.531 ;
      RECT 2.85 3.312 2.86 3.528 ;
      RECT 2.835 3.311 2.85 3.523 ;
      RECT 2.83 3.31 2.835 3.518 ;
      RECT 2.795 3.308 2.83 3.508 ;
      RECT 2.775 3.305 2.795 3.49 ;
      RECT 2.765 3.303 2.775 3.485 ;
      RECT 2.755 3.302 2.765 3.48 ;
      RECT 2.72 3.3 2.755 3.468 ;
      RECT 2.665 3.296 2.72 3.448 ;
      RECT 2.655 3.294 2.665 3.433 ;
      RECT 2.65 3.294 2.655 3.428 ;
      RECT 2.605 3.292 2.65 3.425 ;
      RECT 2.51 3.29 2.56 3.429 ;
      RECT 2.5 3.291 2.51 3.434 ;
      RECT 2.44 3.298 2.5 3.448 ;
      RECT 2.415 3.306 2.44 3.468 ;
      RECT 2.405 3.31 2.415 3.48 ;
      RECT 2.4 3.311 2.405 3.485 ;
      RECT 2.385 3.313 2.4 3.488 ;
      RECT 2.37 3.315 2.385 3.493 ;
      RECT 2.365 3.315 2.37 3.496 ;
      RECT 2.32 3.32 2.365 3.507 ;
      RECT 2.315 3.324 2.32 3.519 ;
      RECT 2.29 3.32 2.315 3.523 ;
      RECT 2.28 3.316 2.29 3.527 ;
      RECT 2.27 3.315 2.28 3.531 ;
      RECT 2.255 3.305 2.27 3.537 ;
      RECT 2.25 3.293 2.255 3.541 ;
      RECT 2.245 3.29 2.25 3.542 ;
      RECT 2.24 3.287 2.245 3.544 ;
      RECT 2.225 3.275 2.24 3.543 ;
      RECT 2.21 3.257 2.225 3.54 ;
      RECT 2.19 3.236 2.21 3.533 ;
      RECT 2.125 3.225 2.19 3.505 ;
      RECT 2.121 3.225 2.125 3.484 ;
      RECT 2.035 3.225 2.121 3.454 ;
      RECT 2.02 3.225 2.035 3.41 ;
      RECT 2.595 2.325 2.6 2.56 ;
      RECT 1.725 2.241 1.73 2.445 ;
      RECT 2.305 2.27 2.31 2.425 ;
      RECT 2.225 2.25 2.23 2.425 ;
      RECT 2.895 2.392 2.91 2.745 ;
      RECT 2.821 2.377 2.895 2.745 ;
      RECT 2.735 2.36 2.821 2.745 ;
      RECT 2.725 2.35 2.735 2.743 ;
      RECT 2.72 2.348 2.725 2.738 ;
      RECT 2.705 2.346 2.72 2.724 ;
      RECT 2.635 2.338 2.705 2.664 ;
      RECT 2.615 2.329 2.635 2.598 ;
      RECT 2.61 2.326 2.615 2.578 ;
      RECT 2.6 2.325 2.61 2.568 ;
      RECT 2.59 2.325 2.595 2.552 ;
      RECT 2.58 2.324 2.59 2.542 ;
      RECT 2.57 2.322 2.58 2.53 ;
      RECT 2.555 2.319 2.57 2.51 ;
      RECT 2.545 2.317 2.555 2.495 ;
      RECT 2.525 2.314 2.545 2.483 ;
      RECT 2.52 2.312 2.525 2.473 ;
      RECT 2.495 2.31 2.52 2.46 ;
      RECT 2.465 2.305 2.495 2.445 ;
      RECT 2.385 2.296 2.465 2.436 ;
      RECT 2.34 2.285 2.385 2.429 ;
      RECT 2.32 2.276 2.34 2.426 ;
      RECT 2.31 2.271 2.32 2.425 ;
      RECT 2.265 2.265 2.305 2.425 ;
      RECT 2.25 2.257 2.265 2.425 ;
      RECT 2.23 2.252 2.25 2.425 ;
      RECT 2.21 2.249 2.225 2.425 ;
      RECT 2.127 2.248 2.21 2.424 ;
      RECT 2.041 2.247 2.127 2.42 ;
      RECT 1.955 2.245 2.041 2.417 ;
      RECT 1.902 2.244 1.955 2.419 ;
      RECT 1.816 2.243 1.902 2.428 ;
      RECT 1.73 2.242 1.816 2.44 ;
      RECT 1.71 2.241 1.725 2.448 ;
      RECT 1.63 2.24 1.71 2.46 ;
      RECT 1.605 2.24 1.63 2.473 ;
      RECT 1.58 2.24 1.605 2.488 ;
      RECT 1.575 2.24 1.58 2.51 ;
      RECT 1.57 2.24 1.575 2.528 ;
      RECT 1.565 2.24 1.57 2.545 ;
      RECT 1.56 2.24 1.565 2.558 ;
      RECT 1.555 2.24 1.56 2.568 ;
      RECT 1.515 2.24 1.555 2.653 ;
      RECT 1.5 2.24 1.515 2.738 ;
      RECT 1.49 2.241 1.5 2.75 ;
      RECT 1.455 2.246 1.49 2.755 ;
      RECT 1.415 2.255 1.455 2.755 ;
      RECT 1.4 2.265 1.415 2.755 ;
      RECT 1.395 2.275 1.4 2.755 ;
      RECT 1.375 2.302 1.395 2.755 ;
      RECT 1.325 2.385 1.375 2.755 ;
      RECT 1.32 2.447 1.325 2.755 ;
      RECT 1.31 2.46 1.32 2.755 ;
      RECT 1.3 2.482 1.31 2.755 ;
      RECT 1.29 2.507 1.3 2.75 ;
      RECT 1.285 2.545 1.29 2.743 ;
      RECT 1.275 2.655 1.285 2.738 ;
      RECT 2.67 3.576 2.685 3.835 ;
      RECT 2.67 3.591 2.69 3.834 ;
      RECT 2.586 3.591 2.69 3.832 ;
      RECT 2.586 3.605 2.695 3.831 ;
      RECT 2.5 3.647 2.7 3.828 ;
      RECT 2.495 3.59 2.685 3.823 ;
      RECT 2.495 3.661 2.705 3.82 ;
      RECT 2.49 3.692 2.705 3.818 ;
      RECT 2.495 3.689 2.72 3.808 ;
      RECT 2.49 3.735 2.735 3.793 ;
      RECT 2.49 3.763 2.74 3.778 ;
      RECT 2.5 3.565 2.67 3.828 ;
      RECT 2.26 2.575 2.43 2.745 ;
      RECT 2.225 2.575 2.43 2.74 ;
      RECT 2.215 2.575 2.43 2.733 ;
      RECT 2.21 2.56 2.38 2.73 ;
      RECT 1.04 3.097 1.305 3.54 ;
      RECT 1.035 3.068 1.25 3.538 ;
      RECT 1.03 3.222 1.31 3.533 ;
      RECT 1.035 3.117 1.31 3.533 ;
      RECT 1.035 3.128 1.32 3.52 ;
      RECT 1.035 3.075 1.28 3.538 ;
      RECT 1.04 3.062 1.25 3.54 ;
      RECT 1.04 3.06 1.2 3.54 ;
      RECT 1.141 3.052 1.2 3.54 ;
      RECT 1.055 3.053 1.2 3.54 ;
      RECT 1.141 3.051 1.19 3.54 ;
      RECT 0.945 1.866 1.12 2.165 ;
      RECT 0.995 1.828 1.12 2.165 ;
      RECT 0.98 1.83 1.206 2.157 ;
      RECT 0.98 1.833 1.245 2.144 ;
      RECT 0.98 1.834 1.255 2.13 ;
      RECT 0.935 1.885 1.255 2.12 ;
      RECT 0.98 1.835 1.26 2.115 ;
      RECT 0.935 2.045 1.265 2.105 ;
      RECT 0.92 1.905 1.26 2.045 ;
      RECT 0.915 1.921 1.26 1.985 ;
      RECT 0.96 1.845 1.26 2.115 ;
      RECT 0.995 1.826 1.081 2.165 ;
      RECT 75.76 0.575 75.93 1.085 ;
      RECT 75.76 2.395 75.93 3.865 ;
      RECT 75.76 5.015 75.93 6.485 ;
      RECT 75.76 7.795 75.93 8.305 ;
      RECT 74.77 0.575 74.94 1.085 ;
      RECT 74.77 2.395 74.94 3.865 ;
      RECT 74.77 5.015 74.94 6.485 ;
      RECT 74.77 7.795 74.94 8.305 ;
      RECT 73.405 0.575 73.575 3.865 ;
      RECT 73.405 5.015 73.575 8.305 ;
      RECT 72.975 0.575 73.145 1.085 ;
      RECT 72.975 1.655 73.145 3.865 ;
      RECT 72.975 5.015 73.145 7.225 ;
      RECT 72.975 7.795 73.145 8.305 ;
      RECT 71.605 1.66 71.775 2.935 ;
      RECT 71.605 5.945 71.775 7.22 ;
      RECT 60.5 0.575 60.67 1.085 ;
      RECT 60.5 2.395 60.67 3.865 ;
      RECT 60.5 5.015 60.67 6.485 ;
      RECT 60.5 7.795 60.67 8.305 ;
      RECT 59.51 0.575 59.68 1.085 ;
      RECT 59.51 2.395 59.68 3.865 ;
      RECT 59.51 5.015 59.68 6.485 ;
      RECT 59.51 7.795 59.68 8.305 ;
      RECT 58.145 0.575 58.315 3.865 ;
      RECT 58.145 5.015 58.315 8.305 ;
      RECT 57.715 0.575 57.885 1.085 ;
      RECT 57.715 1.655 57.885 3.865 ;
      RECT 57.715 5.015 57.885 7.225 ;
      RECT 57.715 7.795 57.885 8.305 ;
      RECT 56.345 1.66 56.515 2.935 ;
      RECT 56.345 5.945 56.515 7.22 ;
      RECT 45.24 0.575 45.41 1.085 ;
      RECT 45.24 2.395 45.41 3.865 ;
      RECT 45.24 5.015 45.41 6.485 ;
      RECT 45.24 7.795 45.41 8.305 ;
      RECT 44.25 0.575 44.42 1.085 ;
      RECT 44.25 2.395 44.42 3.865 ;
      RECT 44.25 5.015 44.42 6.485 ;
      RECT 44.25 7.795 44.42 8.305 ;
      RECT 42.885 0.575 43.055 3.865 ;
      RECT 42.885 5.015 43.055 8.305 ;
      RECT 42.455 0.575 42.625 1.085 ;
      RECT 42.455 1.655 42.625 3.865 ;
      RECT 42.455 5.015 42.625 7.225 ;
      RECT 42.455 7.795 42.625 8.305 ;
      RECT 41.085 1.66 41.255 2.935 ;
      RECT 41.085 5.945 41.255 7.22 ;
      RECT 29.98 0.575 30.15 1.085 ;
      RECT 29.98 2.395 30.15 3.865 ;
      RECT 29.98 5.015 30.15 6.485 ;
      RECT 29.98 7.795 30.15 8.305 ;
      RECT 28.99 0.575 29.16 1.085 ;
      RECT 28.99 2.395 29.16 3.865 ;
      RECT 28.99 5.015 29.16 6.485 ;
      RECT 28.99 7.795 29.16 8.305 ;
      RECT 27.625 0.575 27.795 3.865 ;
      RECT 27.625 5.015 27.795 8.305 ;
      RECT 27.195 0.575 27.365 1.085 ;
      RECT 27.195 1.655 27.365 3.865 ;
      RECT 27.195 5.015 27.365 7.225 ;
      RECT 27.195 7.795 27.365 8.305 ;
      RECT 25.825 1.66 25.995 2.935 ;
      RECT 25.825 5.945 25.995 7.22 ;
      RECT 14.72 0.575 14.89 1.085 ;
      RECT 14.72 2.395 14.89 3.865 ;
      RECT 14.72 5.015 14.89 6.485 ;
      RECT 14.72 7.795 14.89 8.305 ;
      RECT 13.73 0.575 13.9 1.085 ;
      RECT 13.73 2.395 13.9 3.865 ;
      RECT 13.73 5.015 13.9 6.485 ;
      RECT 13.73 7.795 13.9 8.305 ;
      RECT 12.365 0.575 12.535 3.865 ;
      RECT 12.365 5.015 12.535 8.305 ;
      RECT 11.935 0.575 12.105 1.085 ;
      RECT 11.935 1.655 12.105 3.865 ;
      RECT 11.935 5.015 12.105 7.225 ;
      RECT 11.935 7.795 12.105 8.305 ;
      RECT 10.565 1.66 10.735 2.935 ;
      RECT 10.565 5.945 10.735 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2ya_8

MACRO sky130_osu_sc_12T_hs__fill_1
  CLASS CORE ;
  ORIGIN 0.07 0 ;
  FOREIGN sky130_osu_sc_12T_hs__fill_1 -0.07 0 ;
  SIZE 0.275 BY 4.485 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met1 ;
      RECT 0 0 0.11 0.305 ;
      RECT 0 4.135 0.11 4.44 ;
    LAYER li ;
      RECT 0 0 0.11 0.305 ;
      RECT 0 4.135 0.11 4.44 ;
  END
END sky130_osu_sc_12T_hs__fill_1

MACRO sky130_osu_sc_12T_hs__fill_16
  CLASS CORE ;
  ORIGIN 0.045 0 ;
  FOREIGN sky130_osu_sc_12T_hs__fill_16 -0.045 0 ;
  SIZE 1.82 BY 4.485 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met1 ;
      RECT 0 0 1.76 0.305 ;
      RECT 0 4.135 1.76 4.44 ;
    LAYER li ;
      RECT 0 0 1.76 0.305 ;
      RECT 0 4.135 1.76 4.44 ;
  END
END sky130_osu_sc_12T_hs__fill_16

MACRO sky130_osu_sc_12T_hs__fill_2
  CLASS CORE ;
  ORIGIN 0.035 0 ;
  FOREIGN sky130_osu_sc_12T_hs__fill_2 -0.035 0 ;
  SIZE 0.285 BY 4.485 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met1 ;
      RECT 0 0 0.22 0.305 ;
      RECT 0 4.135 0.22 4.44 ;
    LAYER li ;
      RECT 0 0 0.22 0.305 ;
      RECT 0 4.135 0.22 4.44 ;
  END
END sky130_osu_sc_12T_hs__fill_2

MACRO sky130_osu_sc_12T_hs__fill_32
  CLASS CORE ;
  ORIGIN 0.045 0 ;
  FOREIGN sky130_osu_sc_12T_hs__fill_32 -0.045 0 ;
  SIZE 3.58 BY 4.485 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met1 ;
      RECT 0 0 3.52 0.305 ;
      RECT 0 4.135 3.52 4.44 ;
    LAYER li ;
      RECT 0 0 3.52 0.305 ;
      RECT 0 4.135 3.52 4.44 ;
  END
END sky130_osu_sc_12T_hs__fill_32

MACRO sky130_osu_sc_12T_hs__fill_4
  CLASS CORE ;
  ORIGIN 0.045 0 ;
  FOREIGN sky130_osu_sc_12T_hs__fill_4 -0.045 0 ;
  SIZE 0.525 BY 4.485 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met1 ;
      RECT 0 0 0.44 0.305 ;
      RECT 0 4.135 0.44 4.44 ;
    LAYER li ;
      RECT 0 0 0.44 0.305 ;
      RECT 0 4.135 0.44 4.44 ;
  END
END sky130_osu_sc_12T_hs__fill_4

MACRO sky130_osu_sc_12T_hs__fill_8
  CLASS CORE ;
  ORIGIN 0.045 0 ;
  FOREIGN sky130_osu_sc_12T_hs__fill_8 -0.045 0 ;
  SIZE 0.94 BY 4.485 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met1 ;
      RECT 0 0 0.88 0.305 ;
      RECT 0 4.135 0.88 4.44 ;
    LAYER li ;
      RECT 0 0 0.88 0.305 ;
      RECT 0 4.135 0.88 4.44 ;
  END
END sky130_osu_sc_12T_hs__fill_8

MACRO sky130_osu_sc_12T_hs__inv_1
  CLASS CORE ;
  ORIGIN 0.045 0 ;
  FOREIGN sky130_osu_sc_12T_hs__inv_1 -0.045 0 ;
  SIZE 1.04 BY 4.485 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met1 ;
      RECT 0.545 2.365 0.835 2.595 ;
      RECT 0.605 0.885 0.775 2.595 ;
      RECT 0.545 0.885 0.835 1.115 ;
      RECT 0.175 2.735 0.465 2.965 ;
      RECT 0.175 2.765 0.635 2.935 ;
      RECT 0 0 0.99 0.305 ;
      RECT 0 4.135 0.99 4.44 ;
    LAYER mcon ;
      RECT 0.605 0.915 0.775 1.085 ;
      RECT 0.605 2.395 0.775 2.565 ;
      RECT 0.255 0.105 0.425 0.275 ;
      RECT 0.255 4.165 0.425 4.335 ;
      RECT 0.235 2.765 0.405 2.935 ;
    LAYER li ;
      RECT 0.175 0 0.345 0.935 ;
      RECT 0 0 0.99 0.305 ;
      RECT 0 4.135 0.99 4.44 ;
      RECT 0.175 3.405 0.345 4.44 ;
      RECT 0.235 1.74 0.405 2.935 ;
      RECT 0.235 1.74 0.7 1.91 ;
      RECT 0.605 0.575 0.775 1.085 ;
      RECT 0.605 2.395 0.775 3.865 ;
  END
END sky130_osu_sc_12T_hs__inv_1

MACRO sky130_osu_sc_12T_hs__mux2_1
  CLASS CORE ;
  ORIGIN 0.045 0 ;
  FOREIGN sky130_osu_sc_12T_hs__mux2_1 -0.045 0 ;
  SIZE 2.81 BY 4.485 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met1 ;
      RECT 1.925 1.995 2.215 2.225 ;
      RECT 1.755 2.025 2.215 2.195 ;
      RECT 1.495 1.625 1.785 1.855 ;
      RECT 1.555 0.885 1.725 1.855 ;
      RECT 1.495 0.885 1.785 1.115 ;
      RECT 1.12 2.365 1.41 2.595 ;
      RECT 0.95 2.395 1.41 2.565 ;
      RECT 0.125 2.735 0.415 2.965 ;
      RECT 0.125 2.765 0.585 2.935 ;
      RECT 0 0 2.75 0.305 ;
      RECT 0 4.135 2.75 4.44 ;
    LAYER mcon ;
      RECT 2.295 0.105 2.465 0.275 ;
      RECT 2.295 4.165 2.465 4.335 ;
      RECT 1.985 2.025 2.155 2.195 ;
      RECT 1.615 0.105 1.785 0.275 ;
      RECT 1.555 0.915 1.725 1.085 ;
      RECT 1.555 1.655 1.725 1.825 ;
      RECT 1.18 2.395 1.35 2.565 ;
      RECT 0.935 0.105 1.105 0.275 ;
      RECT 0.255 0.105 0.425 0.275 ;
      RECT 0.185 2.765 0.355 2.935 ;
    LAYER li ;
      RECT 0.175 0 0.345 0.935 ;
      RECT 0 0 2.75 0.305 ;
      RECT 0 4.135 2.75 4.44 ;
      RECT 0.175 3.405 0.345 4.44 ;
      RECT 1.125 2.635 1.295 3.865 ;
      RECT 1.18 0.855 1.35 2.805 ;
      RECT 1.125 0.575 1.295 1.025 ;
      RECT 0.605 0.575 0.775 3.865 ;
      RECT 0.605 2.075 1.01 2.405 ;
      RECT 0.605 1.235 1.01 1.565 ;
      RECT 1.985 0.575 2.155 3.865 ;
      RECT 1.555 0.575 1.725 1.085 ;
      RECT 1.555 1.655 1.725 3.865 ;
      RECT 0.185 1.66 0.355 2.935 ;
  END
END sky130_osu_sc_12T_hs__mux2_1

MACRO sky130_osu_single_mpr2aa_8
  CLASS CORE ;
  ORIGIN 9.415 0 ;
  FOREIGN sky130_osu_single_mpr2aa_8 -9.415 0 ;
  SIZE 15.85 BY 8.88 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT -0.75 1.85 -0.42 2.58 ;
      RECT -0.79 1.735 -0.61 2.385 ;
      RECT -4.29 3.535 -3.96 3.865 ;
      RECT -5.495 3.55 -3.96 3.85 ;
      RECT -5.495 2.43 -5.195 3.85 ;
      RECT -5.75 2.415 -5.42 2.745 ;
      RECT -0.27 2.975 0.06 3.705 ;
      RECT -2.35 2.575 -2.02 3.305 ;
      RECT -3.91 2.015 -3.58 2.745 ;
      RECT -4.79 2.015 -4.46 2.745 ;
      RECT -6.47 2.415 -6.14 3.145 ;
      RECT -7.47 1.855 -7.14 2.585 ;
      RECT -8.91 2.575 -8.58 3.305 ;
    LAYER via2 ;
      RECT -0.205 3.04 -0.005 3.24 ;
      RECT -0.685 2.315 -0.485 2.515 ;
      RECT -2.285 3.04 -2.085 3.24 ;
      RECT -3.845 2.48 -3.645 2.68 ;
      RECT -4.225 3.6 -4.025 3.8 ;
      RECT -4.725 2.48 -4.525 2.68 ;
      RECT -5.685 2.48 -5.485 2.68 ;
      RECT -6.405 2.48 -6.205 2.68 ;
      RECT -7.405 1.92 -7.205 2.12 ;
      RECT -8.845 3.04 -8.645 3.24 ;
    LAYER met2 ;
      RECT 2.705 6.28 3.025 6.605 ;
      RECT 2.735 5.695 2.905 6.605 ;
      RECT 2.735 5.695 2.91 6.045 ;
      RECT 2.735 5.695 3.71 5.87 ;
      RECT 3.535 1.965 3.71 5.87 ;
      RECT -0.245 2.84 0.035 3.28 ;
      RECT -0.245 2.84 0.04 3.238 ;
      RECT -0.245 2.84 0.045 3.135 ;
      RECT -0.245 2.84 0.047 3.015 ;
      RECT -0.245 2.84 0.68 3.01 ;
      RECT 0.51 2.025 0.68 3.01 ;
      RECT -0.245 2.805 0.015 3.28 ;
      RECT 3.48 1.965 3.83 2.315 ;
      RECT 0.51 2.025 3.83 2.195 ;
      RECT 3.505 6.655 3.83 6.98 ;
      RECT 2.39 6.745 3.83 6.915 ;
      RECT 2.39 2.395 2.55 6.915 ;
      RECT 2.705 2.365 3.025 2.685 ;
      RECT 2.39 2.395 3.025 2.565 ;
      RECT 1.655 5.855 2.005 6.205 ;
      RECT 1.725 2.705 1.9 6.205 ;
      RECT 1.65 2.705 2 3.055 ;
      RECT -8.885 3 -8.605 3.28 ;
      RECT -8.915 3 -8.605 3.265 ;
      RECT -8.92 2.963 -8.66 3.263 ;
      RECT -8.925 2.964 -8.66 3.257 ;
      RECT -8.93 2.967 -8.66 3.25 ;
      RECT -8.935 3 -8.605 3.243 ;
      RECT -8.965 2.97 -8.66 3.23 ;
      RECT -8.965 2.997 -8.64 3.23 ;
      RECT -8.965 2.987 -8.645 3.23 ;
      RECT -8.965 2.972 -8.65 3.23 ;
      RECT -8.865 2.962 -8.66 3.28 ;
      RECT -8.865 2.957 -8.67 3.28 ;
      RECT -8.865 2.955 -8.685 3.28 ;
      RECT -8.865 1.42 -8.69 3.28 ;
      RECT 1.045 1.34 1.395 1.69 ;
      RECT -8.865 1.42 1.395 1.595 ;
      RECT -3.175 2.455 -2.94 2.715 ;
      RECT -0.03 2.235 0.135 2.495 ;
      RECT -0.125 2.225 -0.11 2.495 ;
      RECT -1.525 1.795 -1.485 1.935 ;
      RECT -0.11 2.23 -0.03 2.495 ;
      RECT -0.165 2.225 -0.125 2.461 ;
      RECT -0.179 2.225 -0.165 2.461 ;
      RECT -0.265 2.23 -0.179 2.463 ;
      RECT -0.31 2.237 -0.265 2.465 ;
      RECT -0.34 2.237 -0.31 2.467 ;
      RECT -0.365 2.232 -0.34 2.469 ;
      RECT -0.395 2.228 -0.365 2.478 ;
      RECT -0.405 2.225 -0.395 2.49 ;
      RECT -0.41 2.225 -0.405 2.498 ;
      RECT -0.415 2.225 -0.41 2.503 ;
      RECT -0.425 2.224 -0.415 2.513 ;
      RECT -0.43 2.223 -0.425 2.523 ;
      RECT -0.445 2.222 -0.43 2.528 ;
      RECT -0.473 2.219 -0.445 2.555 ;
      RECT -0.559 2.211 -0.473 2.555 ;
      RECT -0.645 2.2 -0.559 2.555 ;
      RECT -0.685 2.185 -0.645 2.555 ;
      RECT -0.725 2.159 -0.685 2.555 ;
      RECT -0.73 2.141 -0.725 2.367 ;
      RECT -0.74 2.137 -0.73 2.357 ;
      RECT -0.755 2.127 -0.74 2.344 ;
      RECT -0.775 2.111 -0.755 2.329 ;
      RECT -0.79 2.096 -0.775 2.314 ;
      RECT -0.8 2.085 -0.79 2.304 ;
      RECT -0.825 2.069 -0.8 2.293 ;
      RECT -0.83 2.056 -0.825 2.283 ;
      RECT -0.835 2.052 -0.83 2.278 ;
      RECT -0.89 2.038 -0.835 2.256 ;
      RECT -0.929 2.019 -0.89 2.22 ;
      RECT -1.015 1.993 -0.929 2.173 ;
      RECT -1.019 1.975 -1.015 2.139 ;
      RECT -1.105 1.956 -1.019 2.117 ;
      RECT -1.11 1.938 -1.105 2.095 ;
      RECT -1.115 1.936 -1.11 2.093 ;
      RECT -1.125 1.935 -1.115 2.088 ;
      RECT -1.185 1.922 -1.125 2.074 ;
      RECT -1.23 1.9 -1.185 2.053 ;
      RECT -1.29 1.877 -1.23 2.032 ;
      RECT -1.354 1.852 -1.29 2.007 ;
      RECT -1.44 1.822 -1.354 1.976 ;
      RECT -1.455 1.802 -1.44 1.955 ;
      RECT -1.485 1.797 -1.455 1.946 ;
      RECT -1.538 1.795 -1.525 1.935 ;
      RECT -1.624 1.795 -1.538 1.937 ;
      RECT -1.71 1.795 -1.624 1.939 ;
      RECT -1.73 1.795 -1.71 1.943 ;
      RECT -1.775 1.797 -1.73 1.954 ;
      RECT -1.815 1.807 -1.775 1.97 ;
      RECT -1.819 1.816 -1.815 1.978 ;
      RECT -1.905 1.836 -1.819 1.994 ;
      RECT -1.915 1.855 -1.905 2.012 ;
      RECT -1.92 1.857 -1.915 2.015 ;
      RECT -1.93 1.861 -1.92 2.018 ;
      RECT -1.95 1.866 -1.93 2.028 ;
      RECT -1.98 1.876 -1.95 2.048 ;
      RECT -1.985 1.883 -1.98 2.062 ;
      RECT -1.995 1.887 -1.985 2.069 ;
      RECT -2.01 1.895 -1.995 2.08 ;
      RECT -2.02 1.905 -2.01 2.091 ;
      RECT -2.03 1.912 -2.02 2.099 ;
      RECT -2.055 1.925 -2.03 2.114 ;
      RECT -2.119 1.961 -2.055 2.153 ;
      RECT -2.205 2.024 -2.119 2.217 ;
      RECT -2.24 2.075 -2.205 2.27 ;
      RECT -2.245 2.092 -2.24 2.287 ;
      RECT -2.26 2.101 -2.245 2.294 ;
      RECT -2.28 2.116 -2.26 2.308 ;
      RECT -2.285 2.127 -2.28 2.318 ;
      RECT -2.305 2.14 -2.285 2.328 ;
      RECT -2.31 2.15 -2.305 2.338 ;
      RECT -2.325 2.155 -2.31 2.347 ;
      RECT -2.335 2.165 -2.325 2.358 ;
      RECT -2.365 2.182 -2.335 2.375 ;
      RECT -2.375 2.2 -2.365 2.393 ;
      RECT -2.39 2.211 -2.375 2.404 ;
      RECT -2.43 2.235 -2.39 2.42 ;
      RECT -2.465 2.269 -2.43 2.437 ;
      RECT -2.495 2.292 -2.465 2.449 ;
      RECT -2.51 2.302 -2.495 2.458 ;
      RECT -2.55 2.312 -2.51 2.469 ;
      RECT -2.57 2.323 -2.55 2.481 ;
      RECT -2.575 2.327 -2.57 2.488 ;
      RECT -2.59 2.331 -2.575 2.493 ;
      RECT -2.6 2.336 -2.59 2.498 ;
      RECT -2.605 2.339 -2.6 2.501 ;
      RECT -2.635 2.345 -2.605 2.508 ;
      RECT -2.67 2.355 -2.635 2.522 ;
      RECT -2.73 2.37 -2.67 2.542 ;
      RECT -2.785 2.39 -2.73 2.566 ;
      RECT -2.814 2.405 -2.785 2.584 ;
      RECT -2.9 2.425 -2.814 2.609 ;
      RECT -2.905 2.44 -2.9 2.629 ;
      RECT -2.915 2.443 -2.905 2.63 ;
      RECT -2.94 2.45 -2.915 2.715 ;
      RECT -2.525 3.685 -2.515 3.875 ;
      RECT -4.265 3.56 -3.985 3.84 ;
      RECT -1.22 2.5 -1.215 2.985 ;
      RECT -1.325 2.5 -1.265 2.76 ;
      RECT -1 3.47 -0.995 3.545 ;
      RECT -1.01 3.337 -1 3.58 ;
      RECT -1.02 3.172 -1.01 3.601 ;
      RECT -1.025 3.042 -1.02 3.617 ;
      RECT -1.035 2.932 -1.025 3.633 ;
      RECT -1.04 2.831 -1.035 3.65 ;
      RECT -1.045 2.813 -1.04 3.66 ;
      RECT -1.05 2.795 -1.045 3.67 ;
      RECT -1.06 2.77 -1.05 3.685 ;
      RECT -1.065 2.75 -1.06 3.7 ;
      RECT -1.085 2.5 -1.065 3.725 ;
      RECT -1.1 2.5 -1.085 3.758 ;
      RECT -1.13 2.5 -1.1 3.78 ;
      RECT -1.15 2.5 -1.13 3.794 ;
      RECT -1.17 2.5 -1.15 3.31 ;
      RECT -1.155 3.377 -1.15 3.799 ;
      RECT -1.16 3.407 -1.155 3.801 ;
      RECT -1.165 3.42 -1.16 3.804 ;
      RECT -1.17 3.43 -1.165 3.808 ;
      RECT -1.175 2.5 -1.17 3.228 ;
      RECT -1.175 3.44 -1.17 3.81 ;
      RECT -1.18 2.5 -1.175 3.205 ;
      RECT -1.19 3.462 -1.175 3.81 ;
      RECT -1.195 2.5 -1.18 3.15 ;
      RECT -1.2 3.487 -1.19 3.81 ;
      RECT -1.2 2.5 -1.195 3.095 ;
      RECT -1.21 2.5 -1.2 3.043 ;
      RECT -1.205 3.5 -1.2 3.811 ;
      RECT -1.21 3.512 -1.205 3.812 ;
      RECT -1.215 2.5 -1.21 3.003 ;
      RECT -1.215 3.525 -1.21 3.813 ;
      RECT -1.23 3.54 -1.215 3.814 ;
      RECT -1.225 2.5 -1.22 2.965 ;
      RECT -1.23 2.5 -1.225 2.93 ;
      RECT -1.235 2.5 -1.23 2.905 ;
      RECT -1.24 3.567 -1.23 3.816 ;
      RECT -1.245 2.5 -1.235 2.863 ;
      RECT -1.245 3.585 -1.24 3.817 ;
      RECT -1.25 2.5 -1.245 2.823 ;
      RECT -1.25 3.592 -1.245 3.818 ;
      RECT -1.255 2.5 -1.25 2.795 ;
      RECT -1.26 3.61 -1.25 3.819 ;
      RECT -1.265 2.5 -1.255 2.775 ;
      RECT -1.27 3.63 -1.26 3.821 ;
      RECT -1.28 3.647 -1.27 3.822 ;
      RECT -1.315 3.67 -1.28 3.825 ;
      RECT -1.37 3.688 -1.315 3.831 ;
      RECT -1.456 3.696 -1.37 3.84 ;
      RECT -1.542 3.707 -1.456 3.851 ;
      RECT -1.628 3.717 -1.542 3.862 ;
      RECT -1.714 3.727 -1.628 3.874 ;
      RECT -1.8 3.737 -1.714 3.885 ;
      RECT -1.82 3.743 -1.8 3.891 ;
      RECT -1.9 3.745 -1.82 3.895 ;
      RECT -1.905 3.744 -1.9 3.9 ;
      RECT -1.913 3.743 -1.905 3.9 ;
      RECT -1.999 3.739 -1.913 3.898 ;
      RECT -2.085 3.731 -1.999 3.895 ;
      RECT -2.171 3.722 -2.085 3.891 ;
      RECT -2.257 3.714 -2.171 3.888 ;
      RECT -2.343 3.706 -2.257 3.884 ;
      RECT -2.429 3.697 -2.343 3.881 ;
      RECT -2.515 3.689 -2.429 3.877 ;
      RECT -2.57 3.682 -2.525 3.875 ;
      RECT -2.655 3.675 -2.57 3.873 ;
      RECT -2.729 3.667 -2.655 3.869 ;
      RECT -2.815 3.659 -2.729 3.866 ;
      RECT -2.818 3.655 -2.815 3.864 ;
      RECT -2.904 3.651 -2.818 3.863 ;
      RECT -2.99 3.643 -2.904 3.86 ;
      RECT -3.075 3.638 -2.99 3.857 ;
      RECT -3.161 3.635 -3.075 3.854 ;
      RECT -3.247 3.633 -3.161 3.851 ;
      RECT -3.333 3.63 -3.247 3.848 ;
      RECT -3.419 3.627 -3.333 3.845 ;
      RECT -3.505 3.624 -3.419 3.842 ;
      RECT -3.581 3.622 -3.505 3.839 ;
      RECT -3.667 3.619 -3.581 3.836 ;
      RECT -3.753 3.616 -3.667 3.834 ;
      RECT -3.839 3.614 -3.753 3.831 ;
      RECT -3.925 3.611 -3.839 3.828 ;
      RECT -3.985 3.602 -3.925 3.826 ;
      RECT -1.475 3.22 -1.4 3.48 ;
      RECT -1.495 3.2 -1.49 3.48 ;
      RECT -2.175 2.985 -2.07 3.28 ;
      RECT -7.73 2.96 -7.66 3.22 ;
      RECT -1.835 2.835 -1.83 3.206 ;
      RECT -1.845 2.89 -1.84 3.206 ;
      RECT -1.54 2.06 -1.48 2.32 ;
      RECT -1.485 3.215 -1.475 3.48 ;
      RECT -1.49 3.205 -1.485 3.48 ;
      RECT -1.57 3.152 -1.495 3.48 ;
      RECT -1.545 2.06 -1.54 2.34 ;
      RECT -1.555 2.06 -1.545 2.36 ;
      RECT -1.57 2.06 -1.555 2.39 ;
      RECT -1.585 2.06 -1.57 2.433 ;
      RECT -1.59 3.095 -1.57 3.48 ;
      RECT -1.6 2.06 -1.585 2.47 ;
      RECT -1.605 3.075 -1.59 3.48 ;
      RECT -1.605 2.06 -1.6 2.493 ;
      RECT -1.615 2.06 -1.605 2.518 ;
      RECT -1.645 3.042 -1.605 3.48 ;
      RECT -1.64 2.06 -1.615 2.568 ;
      RECT -1.645 2.06 -1.64 2.623 ;
      RECT -1.65 2.06 -1.645 2.665 ;
      RECT -1.66 3.005 -1.645 3.48 ;
      RECT -1.655 2.06 -1.65 2.708 ;
      RECT -1.66 2.06 -1.655 2.773 ;
      RECT -1.665 2.06 -1.66 2.795 ;
      RECT -1.665 2.993 -1.66 3.345 ;
      RECT -1.67 2.06 -1.665 2.863 ;
      RECT -1.67 2.985 -1.665 3.328 ;
      RECT -1.675 2.06 -1.67 2.908 ;
      RECT -1.68 2.967 -1.67 3.305 ;
      RECT -1.68 2.06 -1.675 2.945 ;
      RECT -1.69 2.06 -1.68 3.285 ;
      RECT -1.695 2.06 -1.69 3.268 ;
      RECT -1.7 2.06 -1.695 3.253 ;
      RECT -1.705 2.06 -1.7 3.238 ;
      RECT -1.725 2.06 -1.705 3.228 ;
      RECT -1.73 2.06 -1.725 3.218 ;
      RECT -1.74 2.06 -1.73 3.214 ;
      RECT -1.745 2.337 -1.74 3.213 ;
      RECT -1.75 2.36 -1.745 3.212 ;
      RECT -1.755 2.39 -1.75 3.211 ;
      RECT -1.76 2.417 -1.755 3.21 ;
      RECT -1.765 2.445 -1.76 3.21 ;
      RECT -1.77 2.472 -1.765 3.21 ;
      RECT -1.775 2.492 -1.77 3.21 ;
      RECT -1.78 2.52 -1.775 3.21 ;
      RECT -1.79 2.562 -1.78 3.21 ;
      RECT -1.8 2.607 -1.79 3.209 ;
      RECT -1.805 2.66 -1.8 3.208 ;
      RECT -1.81 2.692 -1.805 3.207 ;
      RECT -1.815 2.712 -1.81 3.206 ;
      RECT -1.82 2.75 -1.815 3.206 ;
      RECT -1.825 2.772 -1.82 3.206 ;
      RECT -1.83 2.797 -1.825 3.206 ;
      RECT -1.84 2.862 -1.835 3.206 ;
      RECT -1.855 2.922 -1.845 3.206 ;
      RECT -1.87 2.932 -1.855 3.206 ;
      RECT -1.89 2.942 -1.87 3.206 ;
      RECT -1.92 2.947 -1.89 3.203 ;
      RECT -1.98 2.957 -1.92 3.2 ;
      RECT -2 2.966 -1.98 3.205 ;
      RECT -2.025 2.972 -2 3.218 ;
      RECT -2.045 2.977 -2.025 3.233 ;
      RECT -2.07 2.982 -2.045 3.28 ;
      RECT -2.199 2.984 -2.175 3.28 ;
      RECT -2.285 2.979 -2.199 3.28 ;
      RECT -2.325 2.976 -2.285 3.28 ;
      RECT -2.375 2.978 -2.325 3.26 ;
      RECT -2.405 2.982 -2.375 3.26 ;
      RECT -2.484 2.992 -2.405 3.26 ;
      RECT -2.57 3.007 -2.484 3.261 ;
      RECT -2.62 3.017 -2.57 3.262 ;
      RECT -2.628 3.02 -2.62 3.262 ;
      RECT -2.714 3.022 -2.628 3.263 ;
      RECT -2.8 3.026 -2.714 3.263 ;
      RECT -2.886 3.03 -2.8 3.264 ;
      RECT -2.972 3.033 -2.886 3.265 ;
      RECT -3.058 3.037 -2.972 3.265 ;
      RECT -3.144 3.041 -3.058 3.266 ;
      RECT -3.23 3.044 -3.144 3.267 ;
      RECT -3.316 3.048 -3.23 3.267 ;
      RECT -3.402 3.052 -3.316 3.268 ;
      RECT -3.488 3.056 -3.402 3.269 ;
      RECT -3.574 3.059 -3.488 3.269 ;
      RECT -3.66 3.063 -3.574 3.27 ;
      RECT -3.69 3.065 -3.66 3.27 ;
      RECT -3.776 3.068 -3.69 3.271 ;
      RECT -3.862 3.072 -3.776 3.272 ;
      RECT -3.948 3.076 -3.862 3.273 ;
      RECT -4.034 3.079 -3.948 3.273 ;
      RECT -4.12 3.083 -4.034 3.274 ;
      RECT -4.155 3.088 -4.12 3.275 ;
      RECT -4.21 3.098 -4.155 3.282 ;
      RECT -4.235 3.11 -4.21 3.292 ;
      RECT -4.27 3.123 -4.235 3.3 ;
      RECT -4.31 3.14 -4.27 3.323 ;
      RECT -4.33 3.153 -4.31 3.35 ;
      RECT -4.36 3.165 -4.33 3.378 ;
      RECT -4.365 3.173 -4.36 3.398 ;
      RECT -4.37 3.176 -4.365 3.408 ;
      RECT -4.42 3.188 -4.37 3.442 ;
      RECT -4.43 3.203 -4.42 3.475 ;
      RECT -4.44 3.209 -4.43 3.488 ;
      RECT -4.45 3.216 -4.44 3.5 ;
      RECT -4.475 3.229 -4.45 3.518 ;
      RECT -4.49 3.244 -4.475 3.54 ;
      RECT -4.5 3.252 -4.49 3.556 ;
      RECT -4.515 3.261 -4.5 3.571 ;
      RECT -4.525 3.271 -4.515 3.585 ;
      RECT -4.544 3.284 -4.525 3.602 ;
      RECT -4.63 3.329 -4.544 3.667 ;
      RECT -4.645 3.374 -4.63 3.725 ;
      RECT -4.65 3.383 -4.645 3.738 ;
      RECT -4.66 3.39 -4.65 3.743 ;
      RECT -4.665 3.395 -4.66 3.747 ;
      RECT -4.685 3.405 -4.665 3.754 ;
      RECT -4.71 3.425 -4.685 3.768 ;
      RECT -4.745 3.45 -4.71 3.788 ;
      RECT -4.76 3.473 -4.745 3.803 ;
      RECT -4.77 3.483 -4.76 3.808 ;
      RECT -4.78 3.491 -4.77 3.815 ;
      RECT -4.79 3.5 -4.78 3.821 ;
      RECT -4.81 3.512 -4.79 3.823 ;
      RECT -4.82 3.525 -4.81 3.825 ;
      RECT -4.845 3.54 -4.82 3.828 ;
      RECT -4.865 3.557 -4.845 3.832 ;
      RECT -4.905 3.585 -4.865 3.838 ;
      RECT -4.97 3.632 -4.905 3.847 ;
      RECT -4.985 3.665 -4.97 3.855 ;
      RECT -4.99 3.672 -4.985 3.857 ;
      RECT -5.04 3.697 -4.99 3.862 ;
      RECT -5.055 3.721 -5.04 3.869 ;
      RECT -5.105 3.726 -5.055 3.87 ;
      RECT -5.191 3.73 -5.105 3.87 ;
      RECT -5.277 3.73 -5.191 3.87 ;
      RECT -5.363 3.73 -5.277 3.871 ;
      RECT -5.449 3.73 -5.363 3.871 ;
      RECT -5.535 3.73 -5.449 3.871 ;
      RECT -5.601 3.73 -5.535 3.871 ;
      RECT -5.687 3.73 -5.601 3.872 ;
      RECT -5.773 3.73 -5.687 3.872 ;
      RECT -5.859 3.731 -5.773 3.873 ;
      RECT -5.945 3.731 -5.859 3.873 ;
      RECT -6.031 3.731 -5.945 3.873 ;
      RECT -6.117 3.731 -6.031 3.874 ;
      RECT -6.203 3.731 -6.117 3.874 ;
      RECT -6.289 3.732 -6.203 3.875 ;
      RECT -6.375 3.732 -6.289 3.875 ;
      RECT -6.395 3.732 -6.375 3.875 ;
      RECT -6.481 3.732 -6.395 3.875 ;
      RECT -6.567 3.732 -6.481 3.875 ;
      RECT -6.653 3.733 -6.567 3.875 ;
      RECT -6.739 3.733 -6.653 3.875 ;
      RECT -6.825 3.733 -6.739 3.875 ;
      RECT -6.911 3.734 -6.825 3.875 ;
      RECT -6.997 3.734 -6.911 3.875 ;
      RECT -7.083 3.734 -6.997 3.875 ;
      RECT -7.169 3.734 -7.083 3.875 ;
      RECT -7.255 3.735 -7.169 3.875 ;
      RECT -7.305 3.732 -7.255 3.875 ;
      RECT -7.315 3.73 -7.305 3.874 ;
      RECT -7.319 3.73 -7.315 3.873 ;
      RECT -7.405 3.725 -7.319 3.868 ;
      RECT -7.427 3.718 -7.405 3.862 ;
      RECT -7.513 3.709 -7.427 3.856 ;
      RECT -7.599 3.696 -7.513 3.847 ;
      RECT -7.685 3.682 -7.599 3.837 ;
      RECT -7.73 3.672 -7.685 3.83 ;
      RECT -7.75 2.96 -7.73 3.238 ;
      RECT -7.75 3.665 -7.73 3.826 ;
      RECT -7.78 2.96 -7.75 3.26 ;
      RECT -7.79 3.632 -7.75 3.823 ;
      RECT -7.795 2.96 -7.78 3.28 ;
      RECT -7.795 3.597 -7.79 3.821 ;
      RECT -7.8 2.96 -7.795 3.405 ;
      RECT -7.8 3.557 -7.795 3.821 ;
      RECT -7.81 2.96 -7.8 3.821 ;
      RECT -7.885 2.96 -7.81 3.815 ;
      RECT -7.915 2.96 -7.885 3.805 ;
      RECT -7.92 2.96 -7.915 3.797 ;
      RECT -7.925 3.002 -7.92 3.79 ;
      RECT -7.935 3.071 -7.925 3.781 ;
      RECT -7.94 3.141 -7.935 3.733 ;
      RECT -7.945 3.205 -7.94 3.63 ;
      RECT -7.95 3.24 -7.945 3.585 ;
      RECT -7.952 3.277 -7.95 3.477 ;
      RECT -7.955 3.285 -7.952 3.47 ;
      RECT -7.96 3.35 -7.955 3.413 ;
      RECT -3.885 2.44 -3.605 2.72 ;
      RECT -3.895 2.44 -3.605 2.583 ;
      RECT -3.94 2.305 -3.68 2.565 ;
      RECT -3.94 2.42 -3.625 2.565 ;
      RECT -3.94 2.39 -3.63 2.565 ;
      RECT -3.94 2.377 -3.64 2.565 ;
      RECT -3.94 2.367 -3.645 2.565 ;
      RECT -7.965 2.35 -7.705 2.61 ;
      RECT -4.195 1.9 -3.935 2.16 ;
      RECT -4.205 1.925 -3.935 2.12 ;
      RECT -4.21 1.925 -4.205 2.119 ;
      RECT -4.28 1.92 -4.21 2.111 ;
      RECT -4.365 1.907 -4.28 2.094 ;
      RECT -4.369 1.899 -4.365 2.084 ;
      RECT -4.455 1.892 -4.369 2.074 ;
      RECT -4.464 1.884 -4.455 2.064 ;
      RECT -4.55 1.877 -4.464 2.052 ;
      RECT -4.57 1.868 -4.55 2.038 ;
      RECT -4.625 1.863 -4.57 2.03 ;
      RECT -4.635 1.857 -4.625 2.024 ;
      RECT -4.655 1.855 -4.635 2.02 ;
      RECT -4.663 1.854 -4.655 2.016 ;
      RECT -4.749 1.846 -4.663 2.005 ;
      RECT -4.835 1.832 -4.749 1.985 ;
      RECT -4.895 1.82 -4.835 1.97 ;
      RECT -4.905 1.815 -4.895 1.965 ;
      RECT -4.955 1.815 -4.905 1.967 ;
      RECT -5.002 1.817 -4.955 1.971 ;
      RECT -5.088 1.824 -5.002 1.976 ;
      RECT -5.174 1.832 -5.088 1.982 ;
      RECT -5.26 1.841 -5.174 1.988 ;
      RECT -5.319 1.847 -5.26 1.993 ;
      RECT -5.405 1.852 -5.319 1.999 ;
      RECT -5.48 1.857 -5.405 2.005 ;
      RECT -5.519 1.859 -5.48 2.01 ;
      RECT -5.605 1.856 -5.519 2.015 ;
      RECT -5.69 1.854 -5.605 2.022 ;
      RECT -5.722 1.853 -5.69 2.025 ;
      RECT -5.808 1.852 -5.722 2.026 ;
      RECT -5.894 1.851 -5.808 2.027 ;
      RECT -5.98 1.85 -5.894 2.027 ;
      RECT -6.066 1.849 -5.98 2.028 ;
      RECT -6.152 1.848 -6.066 2.029 ;
      RECT -6.238 1.847 -6.152 2.03 ;
      RECT -6.324 1.846 -6.238 2.03 ;
      RECT -6.41 1.845 -6.324 2.031 ;
      RECT -6.46 1.845 -6.41 2.032 ;
      RECT -6.474 1.846 -6.46 2.032 ;
      RECT -6.56 1.853 -6.474 2.033 ;
      RECT -6.634 1.864 -6.56 2.034 ;
      RECT -6.72 1.873 -6.634 2.035 ;
      RECT -6.755 1.88 -6.72 2.05 ;
      RECT -6.78 1.883 -6.755 2.08 ;
      RECT -6.805 1.892 -6.78 2.109 ;
      RECT -6.815 1.903 -6.805 2.129 ;
      RECT -6.825 1.911 -6.815 2.143 ;
      RECT -6.83 1.917 -6.825 2.153 ;
      RECT -6.855 1.934 -6.83 2.17 ;
      RECT -6.87 1.956 -6.855 2.198 ;
      RECT -6.9 1.982 -6.87 2.228 ;
      RECT -6.92 2.011 -6.9 2.258 ;
      RECT -6.925 2.026 -6.92 2.275 ;
      RECT -6.945 2.041 -6.925 2.29 ;
      RECT -6.955 2.059 -6.945 2.308 ;
      RECT -6.965 2.07 -6.955 2.323 ;
      RECT -7.015 2.102 -6.965 2.349 ;
      RECT -7.02 2.132 -7.015 2.369 ;
      RECT -7.03 2.145 -7.02 2.375 ;
      RECT -7.039 2.155 -7.03 2.383 ;
      RECT -7.05 2.166 -7.039 2.391 ;
      RECT -7.055 2.176 -7.05 2.397 ;
      RECT -7.07 2.197 -7.055 2.404 ;
      RECT -7.085 2.227 -7.07 2.412 ;
      RECT -7.12 2.257 -7.085 2.418 ;
      RECT -7.145 2.275 -7.12 2.425 ;
      RECT -7.195 2.283 -7.145 2.434 ;
      RECT -7.22 2.288 -7.195 2.443 ;
      RECT -7.275 2.294 -7.22 2.453 ;
      RECT -7.28 2.299 -7.275 2.461 ;
      RECT -7.294 2.302 -7.28 2.463 ;
      RECT -7.38 2.314 -7.294 2.475 ;
      RECT -7.39 2.326 -7.38 2.488 ;
      RECT -7.475 2.339 -7.39 2.5 ;
      RECT -7.519 2.356 -7.475 2.514 ;
      RECT -7.605 2.373 -7.519 2.53 ;
      RECT -7.635 2.387 -7.605 2.544 ;
      RECT -7.645 2.392 -7.635 2.549 ;
      RECT -7.705 2.395 -7.645 2.558 ;
      RECT -4.815 2.665 -4.555 2.925 ;
      RECT -4.815 2.665 -4.535 2.778 ;
      RECT -4.815 2.665 -4.51 2.745 ;
      RECT -4.815 2.665 -4.505 2.725 ;
      RECT -4.765 2.44 -4.485 2.72 ;
      RECT -5.21 3.175 -4.95 3.435 ;
      RECT -5.22 3.032 -5.025 3.373 ;
      RECT -5.225 3.14 -5.01 3.365 ;
      RECT -5.23 3.19 -4.95 3.355 ;
      RECT -5.24 3.267 -4.95 3.34 ;
      RECT -5.22 3.115 -5.01 3.373 ;
      RECT -5.21 2.99 -5.025 3.435 ;
      RECT -5.21 2.885 -5.045 3.435 ;
      RECT -5.2 2.872 -5.045 3.435 ;
      RECT -5.2 2.83 -5.055 3.435 ;
      RECT -5.195 2.755 -5.055 3.435 ;
      RECT -5.165 2.405 -5.055 3.435 ;
      RECT -5.16 2.135 -5.035 2.758 ;
      RECT -5.19 2.71 -5.035 2.758 ;
      RECT -5.175 2.512 -5.055 3.435 ;
      RECT -5.185 2.622 -5.035 2.758 ;
      RECT -5.16 2.135 -5.02 2.615 ;
      RECT -5.16 2.135 -5 2.49 ;
      RECT -5.195 2.135 -4.935 2.395 ;
      RECT -5.725 2.44 -5.445 2.72 ;
      RECT -5.74 2.44 -5.445 2.7 ;
      RECT -7.685 3.305 -7.425 3.565 ;
      RECT -5.9 3.16 -5.64 3.42 ;
      RECT -5.92 3.18 -5.64 3.395 ;
      RECT -5.963 3.18 -5.92 3.394 ;
      RECT -6.049 3.181 -5.963 3.391 ;
      RECT -6.135 3.182 -6.049 3.387 ;
      RECT -6.21 3.184 -6.135 3.384 ;
      RECT -6.233 3.185 -6.21 3.382 ;
      RECT -6.319 3.186 -6.233 3.38 ;
      RECT -6.405 3.187 -6.319 3.377 ;
      RECT -6.429 3.188 -6.405 3.375 ;
      RECT -6.515 3.19 -6.429 3.372 ;
      RECT -6.6 3.192 -6.515 3.373 ;
      RECT -6.657 3.193 -6.6 3.379 ;
      RECT -6.743 3.195 -6.657 3.389 ;
      RECT -6.829 3.198 -6.743 3.402 ;
      RECT -6.915 3.2 -6.829 3.414 ;
      RECT -6.929 3.201 -6.915 3.421 ;
      RECT -7.015 3.202 -6.929 3.429 ;
      RECT -7.055 3.204 -7.015 3.438 ;
      RECT -7.064 3.205 -7.055 3.441 ;
      RECT -7.15 3.213 -7.064 3.447 ;
      RECT -7.17 3.222 -7.15 3.455 ;
      RECT -7.255 3.237 -7.17 3.463 ;
      RECT -7.315 3.26 -7.255 3.474 ;
      RECT -7.325 3.272 -7.315 3.479 ;
      RECT -7.365 3.282 -7.325 3.483 ;
      RECT -7.42 3.299 -7.365 3.491 ;
      RECT -7.425 3.309 -7.42 3.495 ;
      RECT -6.359 2.44 -6.3 2.837 ;
      RECT -6.445 2.44 -6.24 2.828 ;
      RECT -6.45 2.47 -6.24 2.823 ;
      RECT -6.484 2.47 -6.24 2.821 ;
      RECT -6.57 2.47 -6.24 2.815 ;
      RECT -6.615 2.47 -6.22 2.793 ;
      RECT -6.615 2.47 -6.2 2.748 ;
      RECT -6.655 2.47 -6.2 2.738 ;
      RECT -6.445 2.44 -6.165 2.72 ;
      RECT -6.71 2.44 -6.45 2.7 ;
      RECT -7.525 1.92 -7.265 2.18 ;
      RECT -7.47 1.88 -7.165 2.16 ;
      RECT -7.47 1.855 -7.295 2.18 ;
    LAYER via1 ;
      RECT 3.595 6.74 3.745 6.89 ;
      RECT 3.58 2.065 3.73 2.215 ;
      RECT 2.79 2.45 2.94 2.6 ;
      RECT 2.79 6.37 2.94 6.52 ;
      RECT 1.755 5.955 1.905 6.105 ;
      RECT 1.75 2.805 1.9 2.955 ;
      RECT 1.145 1.44 1.295 1.59 ;
      RECT -0.07 2.29 0.08 2.44 ;
      RECT -0.19 2.86 -0.04 3.01 ;
      RECT -1.27 2.555 -1.12 2.705 ;
      RECT -1.605 3.275 -1.455 3.425 ;
      RECT -1.685 2.115 -1.535 2.265 ;
      RECT -3.12 2.51 -2.97 2.66 ;
      RECT -3.885 2.36 -3.735 2.51 ;
      RECT -4.14 1.955 -3.99 2.105 ;
      RECT -4.76 2.72 -4.61 2.87 ;
      RECT -5.14 2.19 -4.99 2.34 ;
      RECT -5.155 3.23 -5.005 3.38 ;
      RECT -5.685 2.495 -5.535 2.645 ;
      RECT -5.845 3.215 -5.695 3.365 ;
      RECT -6.655 2.495 -6.505 2.645 ;
      RECT -7.47 1.975 -7.32 2.125 ;
      RECT -7.63 3.36 -7.48 3.51 ;
      RECT -7.865 3.015 -7.715 3.165 ;
      RECT -7.91 2.405 -7.76 2.555 ;
      RECT -8.91 3.025 -8.76 3.175 ;
    LAYER met1 ;
      RECT -9.16 1.26 0.5 1.74 ;
      RECT -9.16 1.26 0.555 1.59 ;
      RECT -9.045 0 0.67 1.585 ;
      RECT -9.415 0 6.435 0.305 ;
      RECT -9.41 4.305 6.435 4.745 ;
      RECT -9.16 4.135 6.435 4.745 ;
      RECT -9.16 3.98 0.5 4.745 ;
      RECT 5.835 2.365 6.125 2.595 ;
      RECT 5.895 0.885 6.065 2.595 ;
      RECT 5.835 0.885 6.125 1.115 ;
      RECT 5.835 7.765 6.125 7.995 ;
      RECT 5.895 6.285 6.065 7.995 ;
      RECT 5.835 6.285 6.125 6.515 ;
      RECT 5.425 2.735 5.755 2.965 ;
      RECT 5.425 2.765 5.925 2.935 ;
      RECT 5.425 2.395 5.615 2.965 ;
      RECT 4.845 2.365 5.135 2.595 ;
      RECT 4.845 2.395 5.615 2.565 ;
      RECT 4.905 0.885 5.075 2.595 ;
      RECT 4.845 0.885 5.135 1.115 ;
      RECT 4.845 7.765 5.135 7.995 ;
      RECT 4.905 6.285 5.075 7.995 ;
      RECT 4.845 6.285 5.135 6.515 ;
      RECT 4.845 6.325 5.695 6.485 ;
      RECT 5.525 5.915 5.695 6.485 ;
      RECT 4.845 6.32 5.235 6.485 ;
      RECT 5.465 5.915 5.755 6.145 ;
      RECT 5.465 5.945 5.925 6.115 ;
      RECT 4.475 2.735 4.765 2.965 ;
      RECT 4.475 2.765 4.935 2.935 ;
      RECT 4.535 1.655 4.7 2.965 ;
      RECT 3.05 1.625 3.34 1.855 ;
      RECT 3.05 1.655 4.7 1.825 ;
      RECT 3.11 0.885 3.28 1.855 ;
      RECT 3.05 0.885 3.34 1.115 ;
      RECT 3.05 7.765 3.34 7.995 ;
      RECT 3.11 7.025 3.28 7.995 ;
      RECT 3.11 7.12 4.7 7.29 ;
      RECT 4.53 5.915 4.7 7.29 ;
      RECT 3.05 7.025 3.34 7.255 ;
      RECT 4.475 5.915 4.765 6.145 ;
      RECT 4.475 5.945 4.935 6.115 ;
      RECT 3.48 1.965 3.83 2.315 ;
      RECT 3.31 2.025 3.83 2.195 ;
      RECT 3.505 6.655 3.83 6.98 ;
      RECT 3.48 6.655 3.83 6.885 ;
      RECT 3.31 6.685 3.83 6.855 ;
      RECT 2.705 2.365 3.025 2.685 ;
      RECT 2.675 2.365 3.025 2.595 ;
      RECT 1.145 2.395 3.025 2.565 ;
      RECT 1.145 1.34 1.315 2.565 ;
      RECT 1.045 1.34 1.395 1.69 ;
      RECT 2.705 6.28 3.025 6.605 ;
      RECT 2.675 6.285 3.025 6.515 ;
      RECT 2.505 6.315 3.025 6.485 ;
      RECT 1.65 2.705 2 3.055 ;
      RECT 1.65 2.765 2.14 2.935 ;
      RECT 1.655 5.855 2.005 6.205 ;
      RECT 1.655 5.945 2.14 6.115 ;
      RECT -0.66 2.465 -0.475 2.675 ;
      RECT -0.67 2.47 -0.46 2.668 ;
      RECT -0.67 2.47 -0.374 2.645 ;
      RECT -0.67 2.47 -0.315 2.62 ;
      RECT -0.67 2.47 -0.26 2.6 ;
      RECT -0.67 2.47 -0.25 2.588 ;
      RECT -0.67 2.47 -0.055 2.527 ;
      RECT -0.67 2.47 -0.025 2.51 ;
      RECT -0.67 2.47 -0.005 2.5 ;
      RECT -0.125 2.235 0.135 2.495 ;
      RECT -0.14 2.325 -0.125 2.542 ;
      RECT -0.605 2.457 0.135 2.495 ;
      RECT -0.154 2.336 -0.14 2.548 ;
      RECT -0.565 2.45 0.135 2.495 ;
      RECT -0.24 2.376 -0.154 2.567 ;
      RECT -0.315 2.437 0.135 2.495 ;
      RECT -0.245 2.412 -0.24 2.584 ;
      RECT -0.26 2.422 0.135 2.495 ;
      RECT -0.25 2.417 -0.245 2.586 ;
      RECT 0.045 2.922 0.05 3.014 ;
      RECT 0.04 2.9 0.045 3.031 ;
      RECT 0.035 2.89 0.04 3.043 ;
      RECT 0.025 2.881 0.035 3.053 ;
      RECT 0.02 2.876 0.025 3.061 ;
      RECT 0.015 2.735 0.02 3.064 ;
      RECT -0.019 2.735 0.015 3.075 ;
      RECT -0.105 2.735 -0.019 3.11 ;
      RECT -0.185 2.735 -0.105 3.158 ;
      RECT -0.214 2.735 -0.185 3.182 ;
      RECT -0.3 2.735 -0.214 3.188 ;
      RECT -0.305 2.919 -0.3 3.193 ;
      RECT -0.34 2.93 -0.305 3.196 ;
      RECT -0.365 2.945 -0.34 3.2 ;
      RECT -0.379 2.954 -0.365 3.202 ;
      RECT -0.465 2.981 -0.379 3.208 ;
      RECT -0.53 3.022 -0.465 3.217 ;
      RECT -0.545 3.042 -0.53 3.222 ;
      RECT -0.575 3.052 -0.545 3.225 ;
      RECT -0.58 3.062 -0.575 3.228 ;
      RECT -0.61 3.067 -0.58 3.23 ;
      RECT -0.63 3.072 -0.61 3.234 ;
      RECT -0.715 3.075 -0.63 3.241 ;
      RECT -0.73 3.072 -0.715 3.247 ;
      RECT -0.74 3.069 -0.73 3.249 ;
      RECT -0.76 3.066 -0.74 3.251 ;
      RECT -0.78 3.062 -0.76 3.252 ;
      RECT -0.795 3.058 -0.78 3.254 ;
      RECT -0.805 3.055 -0.795 3.255 ;
      RECT -0.845 3.049 -0.805 3.253 ;
      RECT -0.855 3.044 -0.845 3.251 ;
      RECT -0.87 3.041 -0.855 3.247 ;
      RECT -0.895 3.036 -0.87 3.24 ;
      RECT -0.945 3.027 -0.895 3.228 ;
      RECT -1.015 3.013 -0.945 3.21 ;
      RECT -1.073 2.998 -1.015 3.192 ;
      RECT -1.159 2.981 -1.073 3.172 ;
      RECT -1.245 2.96 -1.159 3.147 ;
      RECT -1.295 2.945 -1.245 3.128 ;
      RECT -1.299 2.939 -1.295 3.12 ;
      RECT -1.385 2.929 -1.299 3.107 ;
      RECT -1.42 2.914 -1.385 3.09 ;
      RECT -1.435 2.907 -1.42 3.083 ;
      RECT -1.495 2.895 -1.435 3.071 ;
      RECT -1.515 2.882 -1.495 3.059 ;
      RECT -1.555 2.873 -1.515 3.051 ;
      RECT -1.56 2.865 -1.555 3.044 ;
      RECT -1.64 2.855 -1.56 3.03 ;
      RECT -1.655 2.842 -1.64 3.015 ;
      RECT -1.66 2.84 -1.655 3.013 ;
      RECT -1.739 2.828 -1.66 3 ;
      RECT -1.825 2.803 -1.739 2.975 ;
      RECT -1.84 2.772 -1.825 2.96 ;
      RECT -1.855 2.747 -1.84 2.956 ;
      RECT -1.87 2.74 -1.855 2.952 ;
      RECT -2.045 2.745 -2.04 2.948 ;
      RECT -2.05 2.75 -2.045 2.943 ;
      RECT -2.04 2.74 -1.87 2.95 ;
      RECT -1.325 2.5 -1.22 2.76 ;
      RECT -0.51 2.025 -0.505 2.25 ;
      RECT -0.38 2.025 -0.325 2.235 ;
      RECT -0.325 2.03 -0.315 2.228 ;
      RECT -0.419 2.025 -0.38 2.238 ;
      RECT -0.505 2.025 -0.419 2.245 ;
      RECT -0.525 2.03 -0.51 2.251 ;
      RECT -0.535 2.07 -0.525 2.253 ;
      RECT -0.565 2.08 -0.535 2.255 ;
      RECT -0.57 2.085 -0.565 2.257 ;
      RECT -0.595 2.09 -0.57 2.259 ;
      RECT -0.61 2.095 -0.595 2.261 ;
      RECT -0.625 2.097 -0.61 2.263 ;
      RECT -0.63 2.102 -0.625 2.265 ;
      RECT -0.68 2.11 -0.63 2.268 ;
      RECT -0.705 2.119 -0.68 2.273 ;
      RECT -0.715 2.126 -0.705 2.278 ;
      RECT -0.72 2.129 -0.715 2.282 ;
      RECT -0.74 2.132 -0.72 2.291 ;
      RECT -0.77 2.14 -0.74 2.311 ;
      RECT -0.799 2.153 -0.77 2.333 ;
      RECT -0.885 2.187 -0.799 2.377 ;
      RECT -0.89 2.213 -0.885 2.415 ;
      RECT -0.895 2.217 -0.89 2.424 ;
      RECT -0.93 2.23 -0.895 2.457 ;
      RECT -0.94 2.244 -0.93 2.495 ;
      RECT -0.945 2.248 -0.94 2.508 ;
      RECT -0.95 2.252 -0.945 2.513 ;
      RECT -0.96 2.26 -0.95 2.525 ;
      RECT -0.965 2.267 -0.96 2.54 ;
      RECT -0.99 2.28 -0.965 2.565 ;
      RECT -1.03 2.309 -0.99 2.62 ;
      RECT -1.045 2.334 -1.03 2.675 ;
      RECT -1.055 2.345 -1.045 2.698 ;
      RECT -1.06 2.352 -1.055 2.71 ;
      RECT -1.065 2.356 -1.06 2.718 ;
      RECT -1.12 2.384 -1.065 2.76 ;
      RECT -1.14 2.42 -1.12 2.76 ;
      RECT -1.155 2.435 -1.14 2.76 ;
      RECT -1.21 2.467 -1.155 2.76 ;
      RECT -1.22 2.497 -1.21 2.76 ;
      RECT -1.61 2.112 -1.425 2.35 ;
      RECT -1.625 2.114 -1.415 2.345 ;
      RECT -1.74 2.06 -1.48 2.32 ;
      RECT -1.745 2.097 -1.48 2.274 ;
      RECT -1.75 2.107 -1.48 2.271 ;
      RECT -1.755 2.147 -1.415 2.265 ;
      RECT -1.76 2.18 -1.415 2.255 ;
      RECT -1.75 2.122 -1.4 2.193 ;
      RECT -1.453 3.22 -1.44 3.75 ;
      RECT -1.539 3.22 -1.44 3.749 ;
      RECT -1.539 3.22 -1.435 3.748 ;
      RECT -1.625 3.22 -1.435 3.746 ;
      RECT -1.63 3.22 -1.435 3.743 ;
      RECT -1.63 3.22 -1.425 3.741 ;
      RECT -1.635 3.512 -1.425 3.738 ;
      RECT -1.635 3.522 -1.42 3.735 ;
      RECT -1.635 3.59 -1.415 3.731 ;
      RECT -1.645 3.595 -1.415 3.73 ;
      RECT -1.645 3.687 -1.41 3.727 ;
      RECT -1.66 3.22 -1.4 3.48 ;
      RECT -2.43 2.21 -2.385 3.745 ;
      RECT -2.23 2.21 -2.2 2.425 ;
      RECT -3.855 1.95 -3.735 2.16 ;
      RECT -4.195 1.9 -3.935 2.16 ;
      RECT -4.195 1.945 -3.9 2.15 ;
      RECT -2.19 2.226 -2.185 2.28 ;
      RECT -2.195 2.219 -2.19 2.413 ;
      RECT -2.2 2.213 -2.195 2.42 ;
      RECT -2.245 2.21 -2.23 2.433 ;
      RECT -2.25 2.21 -2.245 2.455 ;
      RECT -2.255 2.21 -2.25 2.503 ;
      RECT -2.26 2.21 -2.255 2.523 ;
      RECT -2.27 2.21 -2.26 2.63 ;
      RECT -2.275 2.21 -2.27 2.693 ;
      RECT -2.28 2.21 -2.275 2.75 ;
      RECT -2.285 2.21 -2.28 2.758 ;
      RECT -2.3 2.21 -2.285 2.865 ;
      RECT -2.31 2.21 -2.3 3 ;
      RECT -2.32 2.21 -2.31 3.11 ;
      RECT -2.33 2.21 -2.32 3.167 ;
      RECT -2.335 2.21 -2.33 3.207 ;
      RECT -2.34 2.21 -2.335 3.243 ;
      RECT -2.35 2.21 -2.34 3.283 ;
      RECT -2.355 2.21 -2.35 3.325 ;
      RECT -2.375 2.21 -2.355 3.39 ;
      RECT -2.37 3.535 -2.365 3.715 ;
      RECT -2.375 3.517 -2.37 3.723 ;
      RECT -2.38 2.21 -2.375 3.453 ;
      RECT -2.38 3.497 -2.375 3.73 ;
      RECT -2.385 2.21 -2.38 3.74 ;
      RECT -2.44 2.21 -2.43 2.51 ;
      RECT -2.435 2.757 -2.43 3.745 ;
      RECT -2.44 2.822 -2.435 3.745 ;
      RECT -2.445 2.211 -2.44 2.5 ;
      RECT -2.45 2.887 -2.44 3.745 ;
      RECT -2.455 2.212 -2.445 2.49 ;
      RECT -2.465 3 -2.45 3.745 ;
      RECT -2.46 2.213 -2.455 2.48 ;
      RECT -2.48 2.214 -2.46 2.458 ;
      RECT -2.475 3.097 -2.465 3.745 ;
      RECT -2.48 3.172 -2.475 3.745 ;
      RECT -2.49 2.213 -2.48 2.435 ;
      RECT -2.485 3.215 -2.48 3.745 ;
      RECT -2.49 3.242 -2.485 3.745 ;
      RECT -2.5 2.211 -2.49 2.423 ;
      RECT -2.495 3.285 -2.49 3.745 ;
      RECT -2.5 3.312 -2.495 3.745 ;
      RECT -2.51 2.21 -2.5 2.41 ;
      RECT -2.505 3.327 -2.5 3.745 ;
      RECT -2.545 3.385 -2.505 3.745 ;
      RECT -2.515 2.209 -2.51 2.395 ;
      RECT -2.52 2.207 -2.515 2.388 ;
      RECT -2.53 2.204 -2.52 2.378 ;
      RECT -2.535 2.201 -2.53 2.363 ;
      RECT -2.55 2.197 -2.535 2.356 ;
      RECT -2.555 3.44 -2.545 3.745 ;
      RECT -2.555 2.194 -2.55 2.351 ;
      RECT -2.57 2.19 -2.555 2.345 ;
      RECT -2.56 3.457 -2.555 3.745 ;
      RECT -2.57 3.52 -2.56 3.745 ;
      RECT -2.65 2.175 -2.57 2.325 ;
      RECT -2.575 3.527 -2.57 3.74 ;
      RECT -2.58 3.535 -2.575 3.73 ;
      RECT -2.66 2.161 -2.65 2.309 ;
      RECT -2.675 2.157 -2.66 2.307 ;
      RECT -2.685 2.152 -2.675 2.303 ;
      RECT -2.71 2.145 -2.685 2.295 ;
      RECT -2.715 2.14 -2.71 2.29 ;
      RECT -2.725 2.14 -2.715 2.288 ;
      RECT -2.735 2.138 -2.725 2.286 ;
      RECT -2.765 2.13 -2.735 2.28 ;
      RECT -2.78 2.122 -2.765 2.273 ;
      RECT -2.8 2.117 -2.78 2.266 ;
      RECT -2.805 2.113 -2.8 2.261 ;
      RECT -2.835 2.106 -2.805 2.255 ;
      RECT -2.86 2.097 -2.835 2.245 ;
      RECT -2.89 2.09 -2.86 2.237 ;
      RECT -2.915 2.08 -2.89 2.228 ;
      RECT -2.93 2.072 -2.915 2.222 ;
      RECT -2.955 2.067 -2.93 2.217 ;
      RECT -2.965 2.063 -2.955 2.212 ;
      RECT -2.985 2.058 -2.965 2.207 ;
      RECT -3.02 2.053 -2.985 2.2 ;
      RECT -3.08 2.048 -3.02 2.193 ;
      RECT -3.093 2.044 -3.08 2.191 ;
      RECT -3.179 2.039 -3.093 2.188 ;
      RECT -3.265 2.029 -3.179 2.184 ;
      RECT -3.306 2.022 -3.265 2.181 ;
      RECT -3.392 2.015 -3.306 2.178 ;
      RECT -3.478 2.005 -3.392 2.174 ;
      RECT -3.564 1.995 -3.478 2.169 ;
      RECT -3.65 1.985 -3.564 2.165 ;
      RECT -3.66 1.97 -3.65 2.163 ;
      RECT -3.67 1.955 -3.66 2.163 ;
      RECT -3.735 1.95 -3.67 2.162 ;
      RECT -3.9 1.947 -3.855 2.155 ;
      RECT -2.655 2.852 -2.65 3.043 ;
      RECT -2.66 2.847 -2.655 3.05 ;
      RECT -2.674 2.845 -2.66 3.056 ;
      RECT -2.76 2.845 -2.674 3.058 ;
      RECT -2.764 2.845 -2.76 3.061 ;
      RECT -2.85 2.845 -2.764 3.079 ;
      RECT -2.86 2.85 -2.85 3.098 ;
      RECT -2.87 2.905 -2.86 3.102 ;
      RECT -2.895 2.92 -2.87 3.109 ;
      RECT -2.935 2.94 -2.895 3.122 ;
      RECT -2.94 2.952 -2.935 3.132 ;
      RECT -2.955 2.958 -2.94 3.137 ;
      RECT -2.96 2.963 -2.955 3.141 ;
      RECT -2.98 2.97 -2.96 3.146 ;
      RECT -3.05 2.995 -2.98 3.163 ;
      RECT -3.09 3.023 -3.05 3.183 ;
      RECT -3.095 3.033 -3.09 3.191 ;
      RECT -3.115 3.04 -3.095 3.193 ;
      RECT -3.12 3.047 -3.115 3.196 ;
      RECT -3.15 3.055 -3.12 3.199 ;
      RECT -3.155 3.06 -3.15 3.203 ;
      RECT -3.229 3.064 -3.155 3.211 ;
      RECT -3.315 3.073 -3.229 3.227 ;
      RECT -3.319 3.078 -3.315 3.236 ;
      RECT -3.405 3.083 -3.319 3.246 ;
      RECT -3.445 3.091 -3.405 3.258 ;
      RECT -3.495 3.097 -3.445 3.265 ;
      RECT -3.58 3.106 -3.495 3.28 ;
      RECT -3.655 3.117 -3.58 3.298 ;
      RECT -3.69 3.124 -3.655 3.308 ;
      RECT -3.765 3.132 -3.69 3.313 ;
      RECT -3.82 3.141 -3.765 3.313 ;
      RECT -3.845 3.146 -3.82 3.311 ;
      RECT -3.855 3.149 -3.845 3.309 ;
      RECT -3.89 3.151 -3.855 3.307 ;
      RECT -3.92 3.153 -3.89 3.303 ;
      RECT -3.965 3.152 -3.92 3.299 ;
      RECT -3.985 3.147 -3.965 3.296 ;
      RECT -4.035 3.132 -3.985 3.293 ;
      RECT -4.045 3.117 -4.035 3.288 ;
      RECT -4.095 3.102 -4.045 3.278 ;
      RECT -4.145 3.077 -4.095 3.258 ;
      RECT -4.155 3.062 -4.145 3.24 ;
      RECT -4.16 3.06 -4.155 3.234 ;
      RECT -4.18 3.055 -4.16 3.229 ;
      RECT -4.185 3.047 -4.18 3.223 ;
      RECT -4.2 3.041 -4.185 3.216 ;
      RECT -4.205 3.036 -4.2 3.208 ;
      RECT -4.225 3.031 -4.205 3.2 ;
      RECT -4.24 3.024 -4.225 3.193 ;
      RECT -4.255 3.018 -4.24 3.184 ;
      RECT -4.26 3.012 -4.255 3.177 ;
      RECT -4.305 2.987 -4.26 3.163 ;
      RECT -4.32 2.957 -4.305 3.145 ;
      RECT -4.335 2.94 -4.32 3.136 ;
      RECT -4.36 2.92 -4.335 3.124 ;
      RECT -4.4 2.89 -4.36 3.104 ;
      RECT -4.41 2.86 -4.4 3.089 ;
      RECT -4.425 2.85 -4.41 3.082 ;
      RECT -4.48 2.815 -4.425 3.061 ;
      RECT -4.495 2.778 -4.48 3.04 ;
      RECT -4.505 2.765 -4.495 3.032 ;
      RECT -4.555 2.735 -4.505 3.014 ;
      RECT -4.57 2.665 -4.555 2.995 ;
      RECT -4.615 2.665 -4.57 2.978 ;
      RECT -4.64 2.665 -4.615 2.96 ;
      RECT -4.65 2.665 -4.64 2.953 ;
      RECT -4.729 2.665 -4.65 2.946 ;
      RECT -4.815 2.665 -4.729 2.938 ;
      RECT -4.83 2.697 -4.815 2.933 ;
      RECT -4.905 2.707 -4.83 2.929 ;
      RECT -4.925 2.717 -4.905 2.924 ;
      RECT -4.95 2.717 -4.925 2.921 ;
      RECT -4.96 2.707 -4.95 2.92 ;
      RECT -4.97 2.68 -4.96 2.919 ;
      RECT -5.01 2.675 -4.97 2.917 ;
      RECT -5.055 2.675 -5.01 2.913 ;
      RECT -5.08 2.675 -5.055 2.908 ;
      RECT -5.13 2.675 -5.08 2.895 ;
      RECT -5.17 2.68 -5.16 2.88 ;
      RECT -5.16 2.675 -5.13 2.885 ;
      RECT -3.175 2.455 -2.915 2.715 ;
      RECT -3.18 2.477 -2.915 2.673 ;
      RECT -3.94 2.305 -3.72 2.67 ;
      RECT -3.958 2.392 -3.72 2.669 ;
      RECT -3.975 2.397 -3.72 2.666 ;
      RECT -3.975 2.397 -3.7 2.665 ;
      RECT -4.005 2.407 -3.7 2.663 ;
      RECT -4.01 2.422 -3.7 2.659 ;
      RECT -4.01 2.422 -3.695 2.658 ;
      RECT -4.015 2.48 -3.695 2.656 ;
      RECT -4.015 2.48 -3.685 2.653 ;
      RECT -4.02 2.545 -3.685 2.648 ;
      RECT -3.94 2.305 -3.68 2.565 ;
      RECT -5.195 2.135 -4.935 2.395 ;
      RECT -5.195 2.178 -4.849 2.369 ;
      RECT -5.195 2.178 -4.805 2.368 ;
      RECT -5.195 2.178 -4.785 2.366 ;
      RECT -5.195 2.178 -4.685 2.365 ;
      RECT -5.195 2.178 -4.665 2.363 ;
      RECT -5.195 2.178 -4.655 2.358 ;
      RECT -4.785 2.145 -4.595 2.355 ;
      RECT -4.785 2.147 -4.59 2.353 ;
      RECT -4.795 2.152 -4.585 2.345 ;
      RECT -4.849 2.176 -4.585 2.345 ;
      RECT -4.805 2.17 -4.795 2.367 ;
      RECT -4.795 2.15 -4.59 2.353 ;
      RECT -5.84 3.21 -5.635 3.44 ;
      RECT -5.9 3.16 -5.845 3.42 ;
      RECT -5.84 3.16 -5.64 3.44 ;
      RECT -4.87 3.475 -4.865 3.502 ;
      RECT -4.88 3.385 -4.87 3.507 ;
      RECT -4.885 3.307 -4.88 3.513 ;
      RECT -4.895 3.297 -4.885 3.52 ;
      RECT -4.9 3.287 -4.895 3.526 ;
      RECT -4.91 3.282 -4.9 3.528 ;
      RECT -4.925 3.274 -4.91 3.536 ;
      RECT -4.94 3.265 -4.925 3.548 ;
      RECT -4.95 3.257 -4.94 3.558 ;
      RECT -4.985 3.175 -4.95 3.576 ;
      RECT -5.02 3.175 -4.985 3.595 ;
      RECT -5.035 3.175 -5.02 3.603 ;
      RECT -5.09 3.175 -5.035 3.603 ;
      RECT -5.124 3.175 -5.09 3.594 ;
      RECT -5.21 3.175 -5.124 3.57 ;
      RECT -5.22 3.235 -5.21 3.552 ;
      RECT -5.26 3.237 -5.22 3.543 ;
      RECT -5.265 3.239 -5.26 3.533 ;
      RECT -5.285 3.241 -5.265 3.528 ;
      RECT -5.295 3.244 -5.285 3.523 ;
      RECT -5.305 3.245 -5.295 3.518 ;
      RECT -5.329 3.246 -5.305 3.51 ;
      RECT -5.415 3.251 -5.329 3.488 ;
      RECT -5.47 3.25 -5.415 3.461 ;
      RECT -5.485 3.243 -5.47 3.448 ;
      RECT -5.52 3.238 -5.485 3.444 ;
      RECT -5.575 3.23 -5.52 3.443 ;
      RECT -5.635 3.217 -5.575 3.441 ;
      RECT -5.845 3.16 -5.84 3.428 ;
      RECT -5.77 2.53 -5.585 2.74 ;
      RECT -5.78 2.535 -5.57 2.733 ;
      RECT -5.74 2.44 -5.48 2.7 ;
      RECT -5.785 2.597 -5.48 2.623 ;
      RECT -6.44 2.39 -6.435 3.19 ;
      RECT -6.495 2.44 -6.465 3.19 ;
      RECT -6.505 2.44 -6.5 2.75 ;
      RECT -6.52 2.44 -6.515 2.745 ;
      RECT -6.975 2.485 -6.96 2.7 ;
      RECT -7.045 2.485 -6.96 2.695 ;
      RECT -5.78 2.065 -5.71 2.275 ;
      RECT -5.71 2.072 -5.7 2.27 ;
      RECT -5.814 2.065 -5.78 2.282 ;
      RECT -5.9 2.065 -5.814 2.306 ;
      RECT -5.91 2.07 -5.9 2.325 ;
      RECT -5.915 2.082 -5.91 2.328 ;
      RECT -5.93 2.097 -5.915 2.332 ;
      RECT -5.935 2.115 -5.93 2.336 ;
      RECT -5.975 2.125 -5.935 2.345 ;
      RECT -5.99 2.132 -5.975 2.357 ;
      RECT -6.005 2.137 -5.99 2.362 ;
      RECT -6.02 2.14 -6.005 2.367 ;
      RECT -6.03 2.142 -6.02 2.371 ;
      RECT -6.065 2.149 -6.03 2.379 ;
      RECT -6.1 2.157 -6.065 2.393 ;
      RECT -6.11 2.163 -6.1 2.402 ;
      RECT -6.115 2.165 -6.11 2.404 ;
      RECT -6.135 2.168 -6.115 2.41 ;
      RECT -6.165 2.175 -6.135 2.421 ;
      RECT -6.175 2.181 -6.165 2.428 ;
      RECT -6.2 2.184 -6.175 2.435 ;
      RECT -6.21 2.188 -6.2 2.443 ;
      RECT -6.215 2.189 -6.21 2.465 ;
      RECT -6.22 2.19 -6.215 2.48 ;
      RECT -6.225 2.191 -6.22 2.495 ;
      RECT -6.23 2.192 -6.225 2.51 ;
      RECT -6.235 2.193 -6.23 2.54 ;
      RECT -6.245 2.195 -6.235 2.573 ;
      RECT -6.26 2.199 -6.245 2.62 ;
      RECT -6.27 2.202 -6.26 2.665 ;
      RECT -6.275 2.205 -6.27 2.693 ;
      RECT -6.285 2.207 -6.275 2.72 ;
      RECT -6.29 2.21 -6.285 2.755 ;
      RECT -6.32 2.215 -6.29 2.813 ;
      RECT -6.325 2.22 -6.32 2.898 ;
      RECT -6.33 2.222 -6.325 2.933 ;
      RECT -6.335 2.224 -6.33 3.015 ;
      RECT -6.34 2.226 -6.335 3.103 ;
      RECT -6.35 2.228 -6.34 3.185 ;
      RECT -6.365 2.242 -6.35 3.19 ;
      RECT -6.4 2.287 -6.365 3.19 ;
      RECT -6.41 2.327 -6.4 3.19 ;
      RECT -6.425 2.355 -6.41 3.19 ;
      RECT -6.43 2.372 -6.425 3.19 ;
      RECT -6.435 2.38 -6.43 3.19 ;
      RECT -6.445 2.395 -6.44 3.19 ;
      RECT -6.45 2.402 -6.445 3.19 ;
      RECT -6.46 2.422 -6.45 3.19 ;
      RECT -6.465 2.435 -6.46 3.19 ;
      RECT -6.5 2.44 -6.495 2.775 ;
      RECT -6.515 2.83 -6.495 3.19 ;
      RECT -6.515 2.44 -6.505 2.748 ;
      RECT -6.52 2.87 -6.515 3.19 ;
      RECT -6.57 2.44 -6.52 2.743 ;
      RECT -6.525 2.907 -6.52 3.19 ;
      RECT -6.535 2.93 -6.525 3.19 ;
      RECT -6.54 2.975 -6.535 3.19 ;
      RECT -6.55 2.985 -6.54 3.183 ;
      RECT -6.624 2.44 -6.57 2.737 ;
      RECT -6.71 2.44 -6.624 2.73 ;
      RECT -6.759 2.487 -6.71 2.723 ;
      RECT -6.845 2.495 -6.759 2.716 ;
      RECT -6.86 2.492 -6.845 2.711 ;
      RECT -6.874 2.485 -6.86 2.71 ;
      RECT -6.96 2.485 -6.874 2.705 ;
      RECT -7.055 2.49 -7.045 2.69 ;
      RECT -7.465 1.92 -7.45 2.32 ;
      RECT -7.27 1.92 -7.265 2.18 ;
      RECT -7.525 1.92 -7.48 2.18 ;
      RECT -7.07 3.225 -7.065 3.43 ;
      RECT -7.075 3.215 -7.07 3.435 ;
      RECT -7.08 3.202 -7.075 3.44 ;
      RECT -7.085 3.182 -7.08 3.44 ;
      RECT -7.11 3.135 -7.085 3.44 ;
      RECT -7.145 3.05 -7.11 3.44 ;
      RECT -7.15 2.987 -7.145 3.44 ;
      RECT -7.155 2.972 -7.15 3.44 ;
      RECT -7.17 2.932 -7.155 3.44 ;
      RECT -7.175 2.907 -7.17 3.44 ;
      RECT -7.185 2.89 -7.175 3.44 ;
      RECT -7.22 2.812 -7.185 3.44 ;
      RECT -7.225 2.755 -7.22 3.44 ;
      RECT -7.23 2.742 -7.225 3.44 ;
      RECT -7.24 2.72 -7.23 3.44 ;
      RECT -7.25 2.685 -7.24 3.44 ;
      RECT -7.26 2.655 -7.25 3.44 ;
      RECT -7.27 2.57 -7.26 3.083 ;
      RECT -7.263 3.215 -7.26 3.44 ;
      RECT -7.265 3.225 -7.263 3.44 ;
      RECT -7.275 3.235 -7.265 3.435 ;
      RECT -7.28 1.92 -7.27 2.315 ;
      RECT -7.275 2.447 -7.27 3.058 ;
      RECT -7.28 2.345 -7.275 3.041 ;
      RECT -7.29 1.92 -7.28 3.017 ;
      RECT -7.295 1.92 -7.29 2.988 ;
      RECT -7.3 1.92 -7.295 2.978 ;
      RECT -7.32 1.92 -7.3 2.94 ;
      RECT -7.325 1.92 -7.32 2.898 ;
      RECT -7.33 1.92 -7.325 2.878 ;
      RECT -7.36 1.92 -7.33 2.828 ;
      RECT -7.37 1.92 -7.36 2.775 ;
      RECT -7.375 1.92 -7.37 2.748 ;
      RECT -7.38 1.92 -7.375 2.733 ;
      RECT -7.39 1.92 -7.38 2.71 ;
      RECT -7.4 1.92 -7.39 2.685 ;
      RECT -7.405 1.92 -7.4 2.625 ;
      RECT -7.415 1.92 -7.405 2.563 ;
      RECT -7.42 1.92 -7.415 2.483 ;
      RECT -7.425 1.92 -7.42 2.448 ;
      RECT -7.43 1.92 -7.425 2.423 ;
      RECT -7.435 1.92 -7.43 2.408 ;
      RECT -7.44 1.92 -7.435 2.378 ;
      RECT -7.445 1.92 -7.44 2.355 ;
      RECT -7.45 1.92 -7.445 2.328 ;
      RECT -7.48 1.92 -7.465 2.315 ;
      RECT -8.325 3.455 -8.14 3.665 ;
      RECT -8.335 3.46 -8.125 3.658 ;
      RECT -8.335 3.46 -8.105 3.63 ;
      RECT -8.335 3.46 -8.09 3.609 ;
      RECT -8.335 3.46 -8.075 3.607 ;
      RECT -8.335 3.46 -8.065 3.606 ;
      RECT -8.335 3.46 -8.035 3.603 ;
      RECT -7.685 3.305 -7.425 3.565 ;
      RECT -7.725 3.352 -7.425 3.548 ;
      RECT -7.734 3.36 -7.725 3.551 ;
      RECT -8.14 3.453 -7.425 3.548 ;
      RECT -7.82 3.378 -7.734 3.558 ;
      RECT -8.125 3.45 -7.425 3.548 ;
      RECT -7.879 3.4 -7.82 3.57 ;
      RECT -8.105 3.446 -7.425 3.548 ;
      RECT -7.965 3.412 -7.879 3.581 ;
      RECT -8.09 3.442 -7.425 3.548 ;
      RECT -8.02 3.425 -7.965 3.593 ;
      RECT -8.075 3.44 -7.425 3.548 ;
      RECT -8.035 3.431 -8.02 3.599 ;
      RECT -8.065 3.436 -7.425 3.548 ;
      RECT -7.92 2.96 -7.66 3.22 ;
      RECT -7.92 2.98 -7.55 3.19 ;
      RECT -7.92 2.985 -7.54 3.185 ;
      RECT -7.729 2.399 -7.65 2.63 ;
      RECT -7.815 2.402 -7.6 2.625 ;
      RECT -7.82 2.402 -7.6 2.62 ;
      RECT -7.82 2.407 -7.59 2.618 ;
      RECT -7.845 2.407 -7.59 2.615 ;
      RECT -7.845 2.415 -7.58 2.613 ;
      RECT -7.965 2.35 -7.705 2.61 ;
      RECT -7.965 2.397 -7.655 2.61 ;
      RECT -8.71 2.97 -8.705 3.23 ;
      RECT -8.88 2.74 -8.875 3.23 ;
      RECT -8.995 2.98 -8.99 3.205 ;
      RECT -8.285 2.075 -8.28 2.285 ;
      RECT -8.28 2.08 -8.265 2.28 ;
      RECT -8.345 2.075 -8.285 2.293 ;
      RECT -8.36 2.075 -8.345 2.303 ;
      RECT -8.41 2.075 -8.36 2.32 ;
      RECT -8.43 2.075 -8.41 2.343 ;
      RECT -8.445 2.075 -8.43 2.355 ;
      RECT -8.465 2.075 -8.445 2.365 ;
      RECT -8.475 2.08 -8.465 2.374 ;
      RECT -8.48 2.09 -8.475 2.379 ;
      RECT -8.485 2.102 -8.48 2.383 ;
      RECT -8.495 2.125 -8.485 2.388 ;
      RECT -8.5 2.14 -8.495 2.392 ;
      RECT -8.505 2.157 -8.5 2.395 ;
      RECT -8.51 2.165 -8.505 2.398 ;
      RECT -8.52 2.17 -8.51 2.402 ;
      RECT -8.525 2.177 -8.52 2.407 ;
      RECT -8.535 2.182 -8.525 2.411 ;
      RECT -8.56 2.194 -8.535 2.422 ;
      RECT -8.58 2.211 -8.56 2.438 ;
      RECT -8.605 2.228 -8.58 2.46 ;
      RECT -8.64 2.251 -8.605 2.518 ;
      RECT -8.66 2.273 -8.64 2.58 ;
      RECT -8.665 2.283 -8.66 2.615 ;
      RECT -8.675 2.29 -8.665 2.653 ;
      RECT -8.68 2.297 -8.675 2.673 ;
      RECT -8.685 2.308 -8.68 2.71 ;
      RECT -8.69 2.316 -8.685 2.775 ;
      RECT -8.7 2.327 -8.69 2.828 ;
      RECT -8.705 2.345 -8.7 2.898 ;
      RECT -8.71 2.355 -8.705 2.935 ;
      RECT -8.715 2.365 -8.71 3.23 ;
      RECT -8.72 2.377 -8.715 3.23 ;
      RECT -8.725 2.387 -8.72 3.23 ;
      RECT -8.735 2.397 -8.725 3.23 ;
      RECT -8.745 2.42 -8.735 3.23 ;
      RECT -8.76 2.455 -8.745 3.23 ;
      RECT -8.8 2.517 -8.76 3.23 ;
      RECT -8.805 2.57 -8.8 3.23 ;
      RECT -8.83 2.605 -8.805 3.23 ;
      RECT -8.845 2.65 -8.83 3.23 ;
      RECT -8.85 2.672 -8.845 3.23 ;
      RECT -8.86 2.685 -8.85 3.23 ;
      RECT -8.87 2.71 -8.86 3.23 ;
      RECT -8.875 2.732 -8.87 3.23 ;
      RECT -8.9 2.77 -8.88 3.23 ;
      RECT -8.94 2.827 -8.9 3.23 ;
      RECT -8.945 2.877 -8.94 3.23 ;
      RECT -8.95 2.895 -8.945 3.23 ;
      RECT -8.955 2.907 -8.95 3.23 ;
      RECT -8.965 2.925 -8.955 3.23 ;
      RECT -8.975 2.945 -8.965 3.205 ;
      RECT -8.98 2.962 -8.975 3.205 ;
      RECT -8.99 2.975 -8.98 3.205 ;
      RECT -9.02 2.985 -8.995 3.205 ;
      RECT -9.03 2.992 -9.02 3.205 ;
      RECT -9.045 3.002 -9.03 3.2 ;
      RECT -9.415 8.575 6.435 8.88 ;
    LAYER mcon ;
      RECT 5.895 0.915 6.065 1.085 ;
      RECT 5.895 2.395 6.065 2.565 ;
      RECT 5.895 6.315 6.065 6.485 ;
      RECT 5.895 7.795 6.065 7.965 ;
      RECT 5.545 0.105 5.715 0.275 ;
      RECT 5.545 4.165 5.715 4.335 ;
      RECT 5.545 4.545 5.715 4.715 ;
      RECT 5.545 8.605 5.715 8.775 ;
      RECT 5.525 2.765 5.695 2.935 ;
      RECT 5.525 5.945 5.695 6.115 ;
      RECT 4.905 0.915 5.075 1.085 ;
      RECT 4.905 2.395 5.075 2.565 ;
      RECT 4.905 6.315 5.075 6.485 ;
      RECT 4.905 7.795 5.075 7.965 ;
      RECT 4.555 0.105 4.725 0.275 ;
      RECT 4.555 4.165 4.725 4.335 ;
      RECT 4.555 4.545 4.725 4.715 ;
      RECT 4.555 8.605 4.725 8.775 ;
      RECT 4.535 2.765 4.705 2.935 ;
      RECT 4.535 5.945 4.705 6.115 ;
      RECT 3.85 0.105 4.02 0.275 ;
      RECT 3.85 4.165 4.02 4.335 ;
      RECT 3.85 4.545 4.02 4.715 ;
      RECT 3.85 8.605 4.02 8.775 ;
      RECT 3.54 2.025 3.71 2.195 ;
      RECT 3.54 6.685 3.71 6.855 ;
      RECT 3.17 0.105 3.34 0.275 ;
      RECT 3.17 8.605 3.34 8.775 ;
      RECT 3.11 0.915 3.28 1.085 ;
      RECT 3.11 1.655 3.28 1.825 ;
      RECT 3.11 7.055 3.28 7.225 ;
      RECT 3.11 7.795 3.28 7.965 ;
      RECT 2.735 2.395 2.905 2.565 ;
      RECT 2.735 6.315 2.905 6.485 ;
      RECT 2.49 0.105 2.66 0.275 ;
      RECT 2.49 8.605 2.66 8.775 ;
      RECT 1.81 0.105 1.98 0.275 ;
      RECT 1.81 8.605 1.98 8.775 ;
      RECT 1.74 2.765 1.91 2.935 ;
      RECT 1.74 5.945 1.91 6.115 ;
      RECT 0.185 1.415 0.355 1.585 ;
      RECT 0.185 4.135 0.355 4.305 ;
      RECT -0.185 2.875 -0.015 3.045 ;
      RECT -0.275 1.415 -0.105 1.585 ;
      RECT -0.275 4.135 -0.105 4.305 ;
      RECT -0.505 2.045 -0.335 2.215 ;
      RECT -0.65 2.485 -0.48 2.655 ;
      RECT -0.735 1.415 -0.565 1.585 ;
      RECT -0.735 4.135 -0.565 4.305 ;
      RECT -1.195 1.415 -1.025 1.585 ;
      RECT -1.195 4.135 -1.025 4.305 ;
      RECT -1.26 2.525 -1.09 2.695 ;
      RECT -1.605 2.16 -1.435 2.33 ;
      RECT -1.615 3.52 -1.445 3.69 ;
      RECT -1.655 1.415 -1.485 1.585 ;
      RECT -1.655 4.135 -1.485 4.305 ;
      RECT -2.03 2.76 -1.86 2.93 ;
      RECT -2.115 1.415 -1.945 1.585 ;
      RECT -2.115 4.135 -1.945 4.305 ;
      RECT -2.38 2.235 -2.21 2.405 ;
      RECT -2.56 3.55 -2.39 3.72 ;
      RECT -2.575 1.415 -2.405 1.585 ;
      RECT -2.575 4.135 -2.405 4.305 ;
      RECT -2.84 2.865 -2.67 3.035 ;
      RECT -3.035 1.415 -2.865 1.585 ;
      RECT -3.035 4.135 -2.865 4.305 ;
      RECT -3.16 2.49 -2.99 2.66 ;
      RECT -3.495 1.415 -3.325 1.585 ;
      RECT -3.495 4.135 -3.325 4.305 ;
      RECT -3.85 1.97 -3.68 2.14 ;
      RECT -3.925 2.44 -3.755 2.61 ;
      RECT -3.955 1.415 -3.785 1.585 ;
      RECT -3.955 4.135 -3.785 4.305 ;
      RECT -4.415 1.415 -4.245 1.585 ;
      RECT -4.415 4.135 -4.245 4.305 ;
      RECT -4.775 2.165 -4.605 2.335 ;
      RECT -4.875 1.415 -4.705 1.585 ;
      RECT -4.875 4.135 -4.705 4.305 ;
      RECT -5.115 3.36 -4.945 3.53 ;
      RECT -5.15 2.695 -4.98 2.865 ;
      RECT -5.335 1.415 -5.165 1.585 ;
      RECT -5.335 4.135 -5.165 4.305 ;
      RECT -5.76 2.55 -5.59 2.72 ;
      RECT -5.795 1.415 -5.625 1.585 ;
      RECT -5.795 4.135 -5.625 4.305 ;
      RECT -5.83 3.25 -5.66 3.42 ;
      RECT -5.89 2.085 -5.72 2.255 ;
      RECT -6.255 1.415 -6.085 1.585 ;
      RECT -6.255 4.135 -6.085 4.305 ;
      RECT -6.53 3 -6.36 3.17 ;
      RECT -6.715 1.415 -6.545 1.585 ;
      RECT -6.715 4.135 -6.545 4.305 ;
      RECT -7.035 2.505 -6.865 2.675 ;
      RECT -7.175 1.415 -7.005 1.585 ;
      RECT -7.175 4.135 -7.005 4.305 ;
      RECT -7.255 3.25 -7.085 3.42 ;
      RECT -7.46 2.13 -7.29 2.3 ;
      RECT -7.635 1.415 -7.465 1.585 ;
      RECT -7.635 4.135 -7.465 4.305 ;
      RECT -7.73 3 -7.56 3.17 ;
      RECT -7.77 2.43 -7.6 2.6 ;
      RECT -8.095 1.415 -7.925 1.585 ;
      RECT -8.095 4.135 -7.925 4.305 ;
      RECT -8.315 3.475 -8.145 3.645 ;
      RECT -8.455 2.095 -8.285 2.265 ;
      RECT -8.555 1.415 -8.385 1.585 ;
      RECT -8.555 4.135 -8.385 4.305 ;
      RECT -9.015 1.415 -8.845 1.585 ;
      RECT -9.015 4.135 -8.845 4.305 ;
      RECT -9.025 3.015 -8.855 3.185 ;
    LAYER li ;
      RECT -1.03 0 -0.86 2.085 ;
      RECT -2.99 0 -2.82 2.085 ;
      RECT -5.43 0 -5.26 2.085 ;
      RECT -6.39 0 -6.22 2.085 ;
      RECT -6.91 0 -6.74 2.085 ;
      RECT -7.87 0 -7.7 2.085 ;
      RECT -8.83 0 -8.66 2.085 ;
      RECT -9.045 0 0.555 1.59 ;
      RECT -9.16 1.415 0.67 1.585 ;
      RECT -9.045 0 0.67 1.585 ;
      RECT 5.465 0 5.635 0.935 ;
      RECT 4.475 0 4.645 0.935 ;
      RECT 1.73 0 1.9 0.935 ;
      RECT -9.415 0 6.435 0.305 ;
      RECT 5.465 3.405 5.635 5.475 ;
      RECT 4.475 3.405 4.645 5.475 ;
      RECT 1.73 3.405 1.9 5.475 ;
      RECT -9.41 4.305 6.435 4.745 ;
      RECT -9.16 4.135 6.435 4.745 ;
      RECT -0.07 3.635 0.1 4.745 ;
      RECT -1.03 3.635 -0.86 4.745 ;
      RECT -3.47 3.635 -3.3 4.745 ;
      RECT -4.47 3.635 -4.3 4.745 ;
      RECT -5.43 3.635 -5.26 4.745 ;
      RECT -7.87 3.635 -7.7 4.745 ;
      RECT -9.415 8.575 6.435 8.88 ;
      RECT 5.465 7.945 5.635 8.88 ;
      RECT 4.475 7.945 4.645 8.88 ;
      RECT 1.73 7.945 1.9 8.88 ;
      RECT 5.525 1.74 5.695 2.935 ;
      RECT 5.525 1.74 5.99 1.91 ;
      RECT 5.525 6.97 5.99 7.14 ;
      RECT 5.525 5.945 5.695 7.14 ;
      RECT 4.535 1.74 4.705 2.935 ;
      RECT 4.535 1.74 5 1.91 ;
      RECT 4.535 6.97 5 7.14 ;
      RECT 4.535 5.945 4.705 7.14 ;
      RECT 2.68 2.635 2.85 3.865 ;
      RECT 2.735 0.855 2.905 2.805 ;
      RECT 2.68 0.575 2.85 1.025 ;
      RECT 2.68 7.855 2.85 8.305 ;
      RECT 2.735 6.075 2.905 8.025 ;
      RECT 2.68 5.015 2.85 6.245 ;
      RECT 2.16 0.575 2.33 3.865 ;
      RECT 2.16 2.075 2.565 2.405 ;
      RECT 2.16 1.235 2.565 1.565 ;
      RECT 2.16 5.015 2.33 8.305 ;
      RECT 2.16 7.315 2.565 7.645 ;
      RECT 2.16 6.475 2.565 6.805 ;
      RECT -0.505 1.975 0.225 2.215 ;
      RECT 0.037 1.77 0.225 2.215 ;
      RECT -0.135 1.782 0.24 2.209 ;
      RECT -0.22 1.797 0.26 2.194 ;
      RECT -0.22 1.812 0.265 2.184 ;
      RECT -0.265 1.832 0.28 2.176 ;
      RECT -0.288 1.867 0.295 2.13 ;
      RECT -0.374 1.89 0.3 2.09 ;
      RECT -0.374 1.908 0.31 2.06 ;
      RECT -0.505 1.977 0.315 2.023 ;
      RECT -0.46 1.92 0.31 2.06 ;
      RECT -0.374 1.872 0.295 2.13 ;
      RECT -0.288 1.841 0.28 2.176 ;
      RECT -0.265 1.822 0.265 2.184 ;
      RECT -0.22 1.795 0.24 2.209 ;
      RECT -0.135 1.777 0.225 2.215 ;
      RECT -0.049 1.771 0.225 2.215 ;
      RECT 0.037 1.766 0.17 2.215 ;
      RECT 0.123 1.761 0.17 2.215 ;
      RECT -0.185 2.659 -0.015 3.045 ;
      RECT -0.19 2.659 -0.015 3.04 ;
      RECT -0.215 2.659 -0.015 3.005 ;
      RECT -0.215 2.687 -0.005 2.995 ;
      RECT -0.235 2.687 -0.005 2.955 ;
      RECT -0.24 2.687 -0.005 2.928 ;
      RECT -0.24 2.705 0 2.92 ;
      RECT -0.295 2.705 0 2.855 ;
      RECT -0.295 2.722 0.01 2.838 ;
      RECT -0.305 2.722 0.01 2.778 ;
      RECT -0.305 2.739 0.015 2.775 ;
      RECT -0.31 2.575 -0.14 2.753 ;
      RECT -0.31 2.609 -0.054 2.753 ;
      RECT -0.315 3.375 -0.31 3.388 ;
      RECT -0.32 3.27 -0.315 3.393 ;
      RECT -0.345 3.13 -0.32 3.408 ;
      RECT -0.38 3.081 -0.345 3.44 ;
      RECT -0.385 3.049 -0.38 3.46 ;
      RECT -0.39 3.04 -0.385 3.46 ;
      RECT -0.47 3.005 -0.39 3.46 ;
      RECT -0.533 2.975 -0.47 3.46 ;
      RECT -0.619 2.963 -0.533 3.46 ;
      RECT -0.705 2.949 -0.619 3.46 ;
      RECT -0.785 2.936 -0.705 3.446 ;
      RECT -0.82 2.928 -0.785 3.426 ;
      RECT -0.83 2.925 -0.82 3.417 ;
      RECT -0.86 2.92 -0.83 3.404 ;
      RECT -0.91 2.895 -0.86 3.38 ;
      RECT -0.924 2.869 -0.91 3.362 ;
      RECT -1.01 2.829 -0.924 3.338 ;
      RECT -1.055 2.777 -1.01 3.307 ;
      RECT -1.065 2.752 -1.055 3.294 ;
      RECT -1.07 2.533 -1.065 2.555 ;
      RECT -1.075 2.735 -1.065 3.29 ;
      RECT -1.075 2.531 -1.07 2.645 ;
      RECT -1.085 2.527 -1.075 3.286 ;
      RECT -1.129 2.525 -1.085 3.274 ;
      RECT -1.215 2.525 -1.129 3.245 ;
      RECT -1.245 2.525 -1.215 3.218 ;
      RECT -1.26 2.525 -1.245 3.206 ;
      RECT -1.3 2.537 -1.26 3.191 ;
      RECT -1.32 2.556 -1.3 3.17 ;
      RECT -1.33 2.566 -1.32 3.154 ;
      RECT -1.34 2.572 -1.33 3.143 ;
      RECT -1.36 2.582 -1.34 3.126 ;
      RECT -1.365 2.591 -1.36 3.113 ;
      RECT -1.37 2.595 -1.365 3.063 ;
      RECT -1.38 2.601 -1.37 2.98 ;
      RECT -1.385 2.605 -1.38 2.894 ;
      RECT -1.39 2.625 -1.385 2.831 ;
      RECT -1.395 2.648 -1.39 2.778 ;
      RECT -1.4 2.666 -1.395 2.723 ;
      RECT -0.79 2.485 -0.62 2.745 ;
      RECT -0.62 2.45 -0.575 2.731 ;
      RECT -0.659 2.452 -0.57 2.714 ;
      RECT -0.77 2.469 -0.484 2.685 ;
      RECT -0.77 2.484 -0.48 2.657 ;
      RECT -0.77 2.465 -0.57 2.714 ;
      RECT -0.745 2.453 -0.62 2.745 ;
      RECT -0.659 2.451 -0.575 2.731 ;
      RECT -1.605 1.84 -1.435 2.33 ;
      RECT -1.605 1.84 -1.4 2.31 ;
      RECT -1.47 1.76 -1.36 2.27 ;
      RECT -1.489 1.764 -1.34 2.24 ;
      RECT -1.575 1.772 -1.32 2.223 ;
      RECT -1.575 1.778 -1.315 2.213 ;
      RECT -1.575 1.787 -1.295 2.201 ;
      RECT -1.6 1.812 -1.265 2.179 ;
      RECT -1.6 1.832 -1.26 2.159 ;
      RECT -1.605 1.845 -1.25 2.139 ;
      RECT -1.605 1.912 -1.245 2.12 ;
      RECT -1.605 2.045 -1.24 2.107 ;
      RECT -1.61 1.85 -1.25 1.94 ;
      RECT -1.6 1.807 -1.295 2.201 ;
      RECT -1.489 1.762 -1.36 2.27 ;
      RECT -1.615 3.515 -1.315 3.77 ;
      RECT -1.53 3.481 -1.315 3.77 ;
      RECT -1.53 3.484 -1.31 3.63 ;
      RECT -1.595 3.505 -1.31 3.63 ;
      RECT -1.56 3.495 -1.315 3.77 ;
      RECT -1.565 3.5 -1.31 3.63 ;
      RECT -1.53 3.479 -1.329 3.77 ;
      RECT -1.444 3.47 -1.329 3.77 ;
      RECT -1.444 3.464 -1.415 3.77 ;
      RECT -1.955 3.105 -1.945 3.595 ;
      RECT -2.295 3.04 -2.285 3.34 ;
      RECT -1.78 3.212 -1.775 3.431 ;
      RECT -1.79 3.192 -1.78 3.448 ;
      RECT -1.8 3.172 -1.79 3.478 ;
      RECT -1.805 3.162 -1.8 3.493 ;
      RECT -1.81 3.158 -1.805 3.498 ;
      RECT -1.825 3.15 -1.81 3.505 ;
      RECT -1.865 3.13 -1.825 3.53 ;
      RECT -1.89 3.112 -1.865 3.563 ;
      RECT -1.895 3.11 -1.89 3.576 ;
      RECT -1.915 3.107 -1.895 3.58 ;
      RECT -1.945 3.105 -1.915 3.59 ;
      RECT -2.015 3.107 -1.955 3.591 ;
      RECT -2.035 3.107 -2.015 3.585 ;
      RECT -2.06 3.105 -2.035 3.582 ;
      RECT -2.095 3.1 -2.06 3.578 ;
      RECT -2.115 3.094 -2.095 3.565 ;
      RECT -2.125 3.091 -2.115 3.553 ;
      RECT -2.145 3.088 -2.125 3.538 ;
      RECT -2.165 3.084 -2.145 3.52 ;
      RECT -2.17 3.081 -2.165 3.51 ;
      RECT -2.175 3.08 -2.17 3.508 ;
      RECT -2.185 3.077 -2.175 3.5 ;
      RECT -2.195 3.071 -2.185 3.483 ;
      RECT -2.205 3.065 -2.195 3.465 ;
      RECT -2.215 3.059 -2.205 3.453 ;
      RECT -2.225 3.053 -2.215 3.433 ;
      RECT -2.23 3.049 -2.225 3.418 ;
      RECT -2.235 3.047 -2.23 3.41 ;
      RECT -2.24 3.045 -2.235 3.403 ;
      RECT -2.245 3.043 -2.24 3.393 ;
      RECT -2.25 3.041 -2.245 3.387 ;
      RECT -2.26 3.04 -2.25 3.377 ;
      RECT -2.27 3.04 -2.26 3.368 ;
      RECT -2.285 3.04 -2.27 3.353 ;
      RECT -2.325 3.04 -2.295 3.337 ;
      RECT -2.345 3.042 -2.325 3.332 ;
      RECT -2.35 3.047 -2.345 3.33 ;
      RECT -2.38 3.055 -2.35 3.328 ;
      RECT -2.41 3.07 -2.38 3.327 ;
      RECT -2.455 3.092 -2.41 3.332 ;
      RECT -2.46 3.107 -2.455 3.336 ;
      RECT -2.475 3.112 -2.46 3.338 ;
      RECT -2.48 3.116 -2.475 3.34 ;
      RECT -2.54 3.139 -2.48 3.349 ;
      RECT -2.56 3.165 -2.54 3.362 ;
      RECT -2.57 3.172 -2.56 3.366 ;
      RECT -2.585 3.179 -2.57 3.369 ;
      RECT -2.605 3.189 -2.585 3.372 ;
      RECT -2.61 3.197 -2.605 3.375 ;
      RECT -2.655 3.202 -2.61 3.382 ;
      RECT -2.665 3.205 -2.655 3.389 ;
      RECT -2.675 3.205 -2.665 3.393 ;
      RECT -2.71 3.207 -2.675 3.405 ;
      RECT -2.73 3.21 -2.71 3.418 ;
      RECT -2.77 3.213 -2.73 3.429 ;
      RECT -2.785 3.215 -2.77 3.442 ;
      RECT -2.795 3.215 -2.785 3.447 ;
      RECT -2.82 3.216 -2.795 3.455 ;
      RECT -2.83 3.218 -2.82 3.46 ;
      RECT -2.835 3.219 -2.83 3.463 ;
      RECT -2.86 3.217 -2.835 3.466 ;
      RECT -2.875 3.215 -2.86 3.467 ;
      RECT -2.895 3.212 -2.875 3.469 ;
      RECT -2.915 3.207 -2.895 3.469 ;
      RECT -2.975 3.202 -2.915 3.466 ;
      RECT -3.01 3.177 -2.975 3.462 ;
      RECT -3.02 3.154 -3.01 3.46 ;
      RECT -3.05 3.131 -3.02 3.46 ;
      RECT -3.06 3.11 -3.05 3.46 ;
      RECT -3.085 3.092 -3.06 3.458 ;
      RECT -3.1 3.07 -3.085 3.455 ;
      RECT -3.115 3.052 -3.1 3.453 ;
      RECT -3.135 3.042 -3.115 3.451 ;
      RECT -3.15 3.037 -3.135 3.45 ;
      RECT -3.165 3.035 -3.15 3.449 ;
      RECT -3.195 3.036 -3.165 3.447 ;
      RECT -3.215 3.039 -3.195 3.445 ;
      RECT -3.272 3.043 -3.215 3.445 ;
      RECT -3.358 3.052 -3.272 3.445 ;
      RECT -3.444 3.063 -3.358 3.445 ;
      RECT -3.53 3.074 -3.444 3.445 ;
      RECT -3.55 3.081 -3.53 3.453 ;
      RECT -3.56 3.084 -3.55 3.46 ;
      RECT -3.625 3.089 -3.56 3.478 ;
      RECT -3.655 3.096 -3.625 3.503 ;
      RECT -3.665 3.099 -3.655 3.51 ;
      RECT -3.71 3.103 -3.665 3.515 ;
      RECT -3.74 3.108 -3.71 3.52 ;
      RECT -3.741 3.11 -3.74 3.52 ;
      RECT -3.827 3.116 -3.741 3.52 ;
      RECT -3.913 3.127 -3.827 3.52 ;
      RECT -3.999 3.139 -3.913 3.52 ;
      RECT -4.085 3.15 -3.999 3.52 ;
      RECT -4.1 3.157 -4.085 3.515 ;
      RECT -4.105 3.159 -4.1 3.509 ;
      RECT -4.125 3.17 -4.105 3.504 ;
      RECT -4.135 3.188 -4.125 3.498 ;
      RECT -4.14 3.2 -4.135 3.298 ;
      RECT -1.845 1.953 -1.825 2.04 ;
      RECT -1.85 1.888 -1.845 2.072 ;
      RECT -1.86 1.855 -1.85 2.077 ;
      RECT -1.865 1.835 -1.86 2.083 ;
      RECT -1.895 1.835 -1.865 2.1 ;
      RECT -1.944 1.835 -1.895 2.136 ;
      RECT -2.03 1.835 -1.944 2.194 ;
      RECT -2.059 1.845 -2.03 2.243 ;
      RECT -2.145 1.887 -2.059 2.296 ;
      RECT -2.165 1.925 -2.145 2.343 ;
      RECT -2.19 1.942 -2.165 2.363 ;
      RECT -2.2 1.956 -2.19 2.383 ;
      RECT -2.205 1.962 -2.2 2.393 ;
      RECT -2.21 1.966 -2.205 2.4 ;
      RECT -2.26 1.986 -2.21 2.405 ;
      RECT -2.325 2.03 -2.26 2.405 ;
      RECT -2.35 2.08 -2.325 2.405 ;
      RECT -2.36 2.11 -2.35 2.405 ;
      RECT -2.365 2.137 -2.36 2.405 ;
      RECT -2.37 2.155 -2.365 2.405 ;
      RECT -2.38 2.197 -2.37 2.405 ;
      RECT -2.03 2.755 -1.86 2.93 ;
      RECT -2.09 2.583 -2.03 2.918 ;
      RECT -2.1 2.576 -2.09 2.901 ;
      RECT -2.145 2.755 -1.86 2.881 ;
      RECT -2.164 2.755 -1.86 2.859 ;
      RECT -2.25 2.755 -1.86 2.824 ;
      RECT -2.27 2.575 -2.1 2.78 ;
      RECT -2.27 2.722 -1.865 2.78 ;
      RECT -2.27 2.67 -1.89 2.78 ;
      RECT -2.27 2.625 -1.925 2.78 ;
      RECT -2.27 2.607 -1.96 2.78 ;
      RECT -2.27 2.597 -1.965 2.78 ;
      RECT -2.55 3.555 -2.36 3.78 ;
      RECT -2.56 3.556 -2.355 3.775 ;
      RECT -2.56 3.558 -2.345 3.755 ;
      RECT -2.56 3.562 -2.34 3.74 ;
      RECT -2.56 3.549 -2.39 3.775 ;
      RECT -2.56 3.552 -2.365 3.775 ;
      RECT -2.55 3.548 -2.39 3.78 ;
      RECT -2.464 3.546 -2.39 3.78 ;
      RECT -2.84 2.797 -2.67 3.035 ;
      RECT -2.84 2.797 -2.584 2.949 ;
      RECT -2.84 2.797 -2.58 2.859 ;
      RECT -2.79 2.57 -2.57 2.838 ;
      RECT -2.795 2.587 -2.565 2.811 ;
      RECT -2.83 2.745 -2.565 2.811 ;
      RECT -2.81 2.595 -2.67 3.035 ;
      RECT -2.82 2.677 -2.56 2.794 ;
      RECT -2.825 2.725 -2.56 2.794 ;
      RECT -2.82 2.635 -2.565 2.811 ;
      RECT -2.795 2.572 -2.57 2.838 ;
      RECT -3.23 2.547 -3.06 2.745 ;
      RECT -3.23 2.547 -3.015 2.72 ;
      RECT -3.16 2.49 -2.99 2.678 ;
      RECT -3.185 2.505 -2.99 2.678 ;
      RECT -3.57 2.551 -3.54 2.745 ;
      RECT -3.575 2.523 -3.57 2.745 ;
      RECT -3.605 2.497 -3.575 2.747 ;
      RECT -3.63 2.455 -3.605 2.75 ;
      RECT -3.64 2.427 -3.63 2.752 ;
      RECT -3.675 2.407 -3.64 2.754 ;
      RECT -3.74 2.392 -3.675 2.76 ;
      RECT -3.79 2.39 -3.74 2.766 ;
      RECT -3.813 2.392 -3.79 2.771 ;
      RECT -3.899 2.403 -3.813 2.777 ;
      RECT -3.985 2.421 -3.899 2.787 ;
      RECT -4 2.432 -3.985 2.793 ;
      RECT -4.07 2.455 -4 2.799 ;
      RECT -4.125 2.487 -4.07 2.807 ;
      RECT -4.165 2.51 -4.125 2.813 ;
      RECT -4.179 2.523 -4.165 2.816 ;
      RECT -4.265 2.545 -4.179 2.822 ;
      RECT -4.28 2.57 -4.265 2.828 ;
      RECT -4.32 2.585 -4.28 2.832 ;
      RECT -4.37 2.6 -4.32 2.837 ;
      RECT -4.395 2.607 -4.37 2.841 ;
      RECT -4.455 2.602 -4.395 2.845 ;
      RECT -4.47 2.593 -4.455 2.849 ;
      RECT -4.54 2.583 -4.47 2.845 ;
      RECT -4.565 2.575 -4.545 2.835 ;
      RECT -4.624 2.575 -4.565 2.813 ;
      RECT -4.71 2.575 -4.624 2.77 ;
      RECT -4.545 2.575 -4.54 2.84 ;
      RECT -3.85 1.806 -3.68 2.14 ;
      RECT -3.88 1.806 -3.68 2.135 ;
      RECT -3.94 1.773 -3.88 2.123 ;
      RECT -3.94 1.829 -3.67 2.118 ;
      RECT -3.965 1.829 -3.67 2.112 ;
      RECT -3.97 1.77 -3.94 2.109 ;
      RECT -3.985 1.776 -3.85 2.107 ;
      RECT -3.99 1.784 -3.765 2.095 ;
      RECT -3.99 1.836 -3.655 2.048 ;
      RECT -4.005 1.792 -3.765 2.043 ;
      RECT -4.005 1.862 -3.645 1.984 ;
      RECT -4.035 1.812 -3.68 1.945 ;
      RECT -4.035 1.902 -3.635 1.941 ;
      RECT -3.985 1.781 -3.765 2.107 ;
      RECT -4.645 2.111 -4.59 2.375 ;
      RECT -4.645 2.111 -4.525 2.374 ;
      RECT -4.645 2.111 -4.5 2.373 ;
      RECT -4.645 2.111 -4.435 2.372 ;
      RECT -4.5 2.077 -4.42 2.371 ;
      RECT -4.685 2.121 -4.275 2.37 ;
      RECT -4.645 2.118 -4.275 2.37 ;
      RECT -4.685 2.126 -4.27 2.363 ;
      RECT -4.7 2.128 -4.27 2.362 ;
      RECT -4.7 2.135 -4.265 2.358 ;
      RECT -4.72 2.134 -4.27 2.354 ;
      RECT -4.72 2.142 -4.26 2.353 ;
      RECT -4.725 2.139 -4.265 2.349 ;
      RECT -4.725 2.152 -4.25 2.348 ;
      RECT -4.74 2.142 -4.26 2.347 ;
      RECT -4.775 2.155 -4.25 2.34 ;
      RECT -4.59 2.11 -4.28 2.37 ;
      RECT -4.59 2.095 -4.33 2.37 ;
      RECT -4.525 2.082 -4.395 2.37 ;
      RECT -4.98 3.171 -4.965 3.564 ;
      RECT -5.015 3.176 -4.965 3.563 ;
      RECT -4.98 3.175 -4.92 3.562 ;
      RECT -5.035 3.186 -4.92 3.561 ;
      RECT -5.02 3.182 -4.92 3.561 ;
      RECT -5.055 3.192 -4.845 3.558 ;
      RECT -5.055 3.211 -4.8 3.556 ;
      RECT -5.055 3.218 -4.795 3.553 ;
      RECT -5.07 3.195 -4.845 3.55 ;
      RECT -5.09 3.2 -4.845 3.543 ;
      RECT -5.095 3.204 -4.845 3.539 ;
      RECT -5.095 3.221 -4.785 3.538 ;
      RECT -5.115 3.215 -4.8 3.534 ;
      RECT -5.115 3.224 -4.78 3.528 ;
      RECT -5.12 3.23 -4.78 3.3 ;
      RECT -5.055 3.19 -4.92 3.558 ;
      RECT -5.18 2.553 -4.98 2.865 ;
      RECT -5.105 2.531 -4.98 2.865 ;
      RECT -5.165 2.55 -4.975 2.85 ;
      RECT -5.195 2.561 -4.975 2.848 ;
      RECT -5.18 2.556 -4.97 2.814 ;
      RECT -5.195 2.66 -4.965 2.781 ;
      RECT -5.165 2.532 -4.98 2.865 ;
      RECT -5.105 2.51 -5.005 2.865 ;
      RECT -5.08 2.507 -5.005 2.865 ;
      RECT -5.08 2.502 -5.06 2.865 ;
      RECT -5.675 2.57 -5.5 2.745 ;
      RECT -5.68 2.57 -5.5 2.743 ;
      RECT -5.705 2.57 -5.5 2.738 ;
      RECT -5.76 2.55 -5.59 2.728 ;
      RECT -5.76 2.557 -5.525 2.728 ;
      RECT -5.675 3.237 -5.66 3.42 ;
      RECT -5.685 3.215 -5.675 3.42 ;
      RECT -5.7 3.195 -5.685 3.42 ;
      RECT -5.71 3.17 -5.7 3.42 ;
      RECT -5.74 3.135 -5.71 3.42 ;
      RECT -5.775 3.075 -5.74 3.42 ;
      RECT -5.78 3.037 -5.775 3.42 ;
      RECT -5.83 2.988 -5.78 3.42 ;
      RECT -5.84 2.938 -5.83 3.408 ;
      RECT -5.855 2.917 -5.84 3.368 ;
      RECT -5.875 2.885 -5.855 3.318 ;
      RECT -5.9 2.841 -5.875 3.258 ;
      RECT -5.905 2.813 -5.9 3.213 ;
      RECT -5.91 2.804 -5.905 3.199 ;
      RECT -5.915 2.797 -5.91 3.186 ;
      RECT -5.92 2.792 -5.915 3.175 ;
      RECT -5.925 2.777 -5.92 3.165 ;
      RECT -5.93 2.755 -5.925 3.152 ;
      RECT -5.94 2.715 -5.93 3.127 ;
      RECT -5.965 2.645 -5.94 3.083 ;
      RECT -5.97 2.585 -5.965 3.048 ;
      RECT -5.985 2.565 -5.97 3.015 ;
      RECT -5.99 2.565 -5.985 2.99 ;
      RECT -6.02 2.565 -5.99 2.945 ;
      RECT -6.065 2.565 -6.02 2.885 ;
      RECT -6.14 2.565 -6.065 2.833 ;
      RECT -6.145 2.565 -6.14 2.798 ;
      RECT -6.15 2.565 -6.145 2.788 ;
      RECT -6.155 2.565 -6.15 2.768 ;
      RECT -5.89 1.785 -5.72 2.255 ;
      RECT -5.945 1.778 -5.75 2.239 ;
      RECT -5.945 1.792 -5.715 2.238 ;
      RECT -5.96 1.793 -5.715 2.219 ;
      RECT -5.965 1.811 -5.715 2.205 ;
      RECT -5.96 1.794 -5.71 2.203 ;
      RECT -5.975 1.825 -5.71 2.188 ;
      RECT -5.96 1.8 -5.705 2.173 ;
      RECT -5.98 1.84 -5.705 2.17 ;
      RECT -5.965 1.812 -5.7 2.155 ;
      RECT -5.965 1.824 -5.695 2.135 ;
      RECT -5.98 1.84 -5.69 2.118 ;
      RECT -5.98 1.85 -5.685 1.973 ;
      RECT -5.985 1.85 -5.685 1.93 ;
      RECT -5.985 1.865 -5.68 1.908 ;
      RECT -5.89 1.775 -5.75 2.255 ;
      RECT -5.89 1.773 -5.78 2.255 ;
      RECT -5.804 1.77 -5.78 2.255 ;
      RECT -6.145 3.437 -6.14 3.483 ;
      RECT -6.155 3.285 -6.145 3.507 ;
      RECT -6.16 3.13 -6.155 3.532 ;
      RECT -6.175 3.092 -6.16 3.543 ;
      RECT -6.18 3.075 -6.175 3.55 ;
      RECT -6.19 3.063 -6.18 3.557 ;
      RECT -6.195 3.054 -6.19 3.559 ;
      RECT -6.2 3.052 -6.195 3.563 ;
      RECT -6.245 3.043 -6.2 3.578 ;
      RECT -6.25 3.035 -6.245 3.592 ;
      RECT -6.255 3.032 -6.25 3.596 ;
      RECT -6.27 3.027 -6.255 3.604 ;
      RECT -6.325 3.017 -6.27 3.615 ;
      RECT -6.36 3.005 -6.325 3.616 ;
      RECT -6.369 3 -6.36 3.61 ;
      RECT -6.455 3 -6.369 3.6 ;
      RECT -6.485 3 -6.455 3.578 ;
      RECT -6.495 3 -6.49 3.558 ;
      RECT -6.5 3 -6.495 3.52 ;
      RECT -6.505 3 -6.5 3.478 ;
      RECT -6.51 3 -6.505 3.438 ;
      RECT -6.515 3 -6.51 3.368 ;
      RECT -6.525 3 -6.515 3.29 ;
      RECT -6.53 3 -6.525 3.19 ;
      RECT -6.49 3 -6.485 3.56 ;
      RECT -6.995 3.082 -6.905 3.56 ;
      RECT -7.01 3.085 -6.89 3.558 ;
      RECT -6.995 3.084 -6.89 3.558 ;
      RECT -7.03 3.091 -6.865 3.548 ;
      RECT -7.01 3.085 -6.865 3.548 ;
      RECT -7.045 3.097 -6.865 3.536 ;
      RECT -7.01 3.088 -6.815 3.529 ;
      RECT -7.059 3.105 -6.815 3.527 ;
      RECT -7.03 3.095 -6.805 3.515 ;
      RECT -7.059 3.116 -6.775 3.506 ;
      RECT -7.145 3.14 -6.775 3.5 ;
      RECT -7.145 3.153 -6.735 3.483 ;
      RECT -7.15 3.175 -6.735 3.476 ;
      RECT -7.18 3.19 -6.735 3.466 ;
      RECT -7.185 3.201 -6.735 3.456 ;
      RECT -7.215 3.214 -6.735 3.447 ;
      RECT -7.23 3.232 -6.735 3.436 ;
      RECT -7.255 3.245 -6.735 3.426 ;
      RECT -6.995 3.081 -6.985 3.56 ;
      RECT -6.949 2.505 -6.91 2.75 ;
      RECT -7.035 2.505 -6.9 2.748 ;
      RECT -7.15 2.53 -6.9 2.745 ;
      RECT -7.15 2.53 -6.895 2.743 ;
      RECT -7.15 2.53 -6.88 2.738 ;
      RECT -7.044 2.505 -6.865 2.718 ;
      RECT -7.13 2.513 -6.865 2.718 ;
      RECT -7.46 1.865 -7.29 2.3 ;
      RECT -7.47 1.899 -7.29 2.283 ;
      RECT -7.39 1.835 -7.22 2.27 ;
      RECT -7.485 1.91 -7.22 2.248 ;
      RECT -7.39 1.845 -7.215 2.238 ;
      RECT -7.46 1.897 -7.185 2.223 ;
      RECT -7.5 1.923 -7.185 2.208 ;
      RECT -7.5 1.965 -7.175 2.188 ;
      RECT -7.505 1.99 -7.17 2.17 ;
      RECT -7.505 2 -7.165 2.155 ;
      RECT -7.51 1.937 -7.185 2.153 ;
      RECT -7.51 2.01 -7.16 2.138 ;
      RECT -7.515 1.947 -7.185 2.135 ;
      RECT -7.52 2.031 -7.155 2.118 ;
      RECT -7.52 2.063 -7.15 2.098 ;
      RECT -7.525 1.977 -7.175 2.09 ;
      RECT -7.52 1.962 -7.185 2.118 ;
      RECT -7.505 1.932 -7.185 2.17 ;
      RECT -7.66 2.519 -7.435 2.775 ;
      RECT -7.66 2.552 -7.415 2.765 ;
      RECT -7.695 2.552 -7.415 2.763 ;
      RECT -7.695 2.565 -7.41 2.753 ;
      RECT -7.695 2.585 -7.4 2.745 ;
      RECT -7.695 2.682 -7.395 2.738 ;
      RECT -7.715 2.43 -7.585 2.728 ;
      RECT -7.76 2.585 -7.4 2.67 ;
      RECT -7.77 2.43 -7.585 2.615 ;
      RECT -7.77 2.462 -7.499 2.615 ;
      RECT -7.805 2.992 -7.785 3.17 ;
      RECT -7.84 2.945 -7.805 3.17 ;
      RECT -7.855 2.885 -7.84 3.17 ;
      RECT -7.88 2.832 -7.855 3.17 ;
      RECT -7.895 2.785 -7.88 3.17 ;
      RECT -7.915 2.762 -7.895 3.17 ;
      RECT -7.94 2.727 -7.915 3.17 ;
      RECT -7.95 2.573 -7.94 3.17 ;
      RECT -7.98 2.568 -7.95 3.161 ;
      RECT -7.985 2.565 -7.98 3.151 ;
      RECT -8 2.565 -7.985 3.125 ;
      RECT -8.005 2.565 -8 3.088 ;
      RECT -8.03 2.565 -8.005 3.04 ;
      RECT -8.05 2.565 -8.03 2.965 ;
      RECT -8.06 2.565 -8.05 2.925 ;
      RECT -8.065 2.565 -8.06 2.9 ;
      RECT -8.07 2.565 -8.065 2.883 ;
      RECT -8.075 2.565 -8.07 2.865 ;
      RECT -8.08 2.566 -8.075 2.855 ;
      RECT -8.09 2.568 -8.08 2.823 ;
      RECT -8.1 2.57 -8.09 2.79 ;
      RECT -8.11 2.573 -8.1 2.763 ;
      RECT -7.785 3 -7.56 3.17 ;
      RECT -8.455 1.812 -8.285 2.265 ;
      RECT -8.455 1.812 -8.195 2.231 ;
      RECT -8.455 1.812 -8.165 2.215 ;
      RECT -8.455 1.812 -8.135 2.188 ;
      RECT -8.199 1.79 -8.12 2.17 ;
      RECT -8.42 1.797 -8.115 2.155 ;
      RECT -8.42 1.805 -8.105 2.118 ;
      RECT -8.46 1.832 -8.105 2.09 ;
      RECT -8.475 1.845 -8.105 2.055 ;
      RECT -8.455 1.82 -8.085 2.045 ;
      RECT -8.48 1.885 -8.085 2.015 ;
      RECT -8.48 1.915 -8.08 1.998 ;
      RECT -8.485 1.945 -8.08 1.985 ;
      RECT -8.42 1.794 -8.12 2.17 ;
      RECT -8.285 1.791 -8.199 2.249 ;
      RECT -8.334 1.792 -8.12 2.17 ;
      RECT -8.19 3.452 -8.145 3.645 ;
      RECT -8.2 3.422 -8.19 3.645 ;
      RECT -8.205 3.407 -8.2 3.645 ;
      RECT -8.245 3.317 -8.205 3.645 ;
      RECT -8.25 3.23 -8.245 3.645 ;
      RECT -8.26 3.2 -8.25 3.645 ;
      RECT -8.265 3.16 -8.26 3.645 ;
      RECT -8.275 3.122 -8.265 3.645 ;
      RECT -8.28 3.087 -8.275 3.645 ;
      RECT -8.3 3.04 -8.28 3.645 ;
      RECT -8.315 2.965 -8.3 3.645 ;
      RECT -8.32 2.92 -8.315 3.64 ;
      RECT -8.325 2.9 -8.32 3.613 ;
      RECT -8.33 2.88 -8.325 3.598 ;
      RECT -8.335 2.855 -8.33 3.578 ;
      RECT -8.34 2.833 -8.335 3.563 ;
      RECT -8.345 2.811 -8.34 3.545 ;
      RECT -8.35 2.79 -8.345 3.535 ;
      RECT -8.36 2.762 -8.35 3.505 ;
      RECT -8.37 2.725 -8.36 3.473 ;
      RECT -8.38 2.685 -8.37 3.44 ;
      RECT -8.39 2.663 -8.38 3.41 ;
      RECT -8.42 2.615 -8.39 3.342 ;
      RECT -8.435 2.575 -8.42 3.269 ;
      RECT -8.445 2.575 -8.435 3.235 ;
      RECT -8.45 2.575 -8.445 3.21 ;
      RECT -8.455 2.575 -8.45 3.195 ;
      RECT -8.46 2.575 -8.455 3.173 ;
      RECT -8.465 2.575 -8.46 3.16 ;
      RECT -8.48 2.575 -8.465 3.125 ;
      RECT -8.5 2.575 -8.48 3.065 ;
      RECT -8.51 2.575 -8.5 3.015 ;
      RECT -8.53 2.575 -8.51 2.963 ;
      RECT -8.55 2.575 -8.53 2.92 ;
      RECT -8.56 2.575 -8.55 2.908 ;
      RECT -8.59 2.575 -8.56 2.895 ;
      RECT -8.62 2.596 -8.59 2.875 ;
      RECT -8.63 2.624 -8.62 2.855 ;
      RECT -8.645 2.641 -8.63 2.823 ;
      RECT -8.65 2.655 -8.645 2.79 ;
      RECT -8.655 2.663 -8.65 2.763 ;
      RECT -8.66 2.671 -8.655 2.725 ;
      RECT -8.655 3.195 -8.65 3.53 ;
      RECT -8.69 3.182 -8.655 3.529 ;
      RECT -8.76 3.122 -8.69 3.528 ;
      RECT -8.84 3.065 -8.76 3.527 ;
      RECT -8.975 3.025 -8.84 3.526 ;
      RECT -8.975 3.212 -8.64 3.515 ;
      RECT -9.015 3.212 -8.64 3.505 ;
      RECT -9.015 3.23 -8.635 3.5 ;
      RECT -9.015 3.32 -8.63 3.49 ;
      RECT -9.02 3.015 -8.855 3.47 ;
      RECT -9.025 3.015 -8.855 3.213 ;
      RECT -9.025 3.172 -8.66 3.213 ;
      RECT -9.025 3.16 -8.665 3.213 ;
      RECT 5.895 0.575 6.065 1.085 ;
      RECT 5.895 2.395 6.065 3.865 ;
      RECT 5.895 5.015 6.065 6.485 ;
      RECT 5.895 7.795 6.065 8.305 ;
      RECT 4.905 0.575 5.075 1.085 ;
      RECT 4.905 2.395 5.075 3.865 ;
      RECT 4.905 5.015 5.075 6.485 ;
      RECT 4.905 7.795 5.075 8.305 ;
      RECT 3.54 0.575 3.71 3.865 ;
      RECT 3.54 5.015 3.71 8.305 ;
      RECT 3.11 0.575 3.28 1.085 ;
      RECT 3.11 1.655 3.28 3.865 ;
      RECT 3.11 5.015 3.28 7.225 ;
      RECT 3.11 7.795 3.28 8.305 ;
      RECT 1.74 1.66 1.91 2.935 ;
      RECT 1.74 5.945 1.91 7.22 ;
  END
END sky130_osu_single_mpr2aa_8

MACRO sky130_osu_single_mpr2at_8
  CLASS CORE ;
  ORIGIN 11.495 0 ;
  FOREIGN sky130_osu_single_mpr2at_8 -11.495 0 ;
  SIZE 17.93 BY 8.88 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT -1.81 3.685 -1.255 4.015 ;
      RECT -1.81 2.02 -1.51 4.015 ;
      RECT -5.745 3.125 -5.19 3.455 ;
      RECT -5.49 2.02 -5.19 3.455 ;
      RECT -4.695 1.885 -4.545 2.535 ;
      RECT -5.49 2.02 -1.51 2.32 ;
      RECT -0.625 2.005 0.105 2.335 ;
      RECT -2.845 3.685 -2.115 4.015 ;
      RECT -4.545 3.685 -3.815 4.015 ;
      RECT -6.985 2.565 -6.255 2.895 ;
      RECT -8.425 3.125 -7.695 3.455 ;
      RECT -9.5 2.565 -8.77 2.895 ;
      RECT -10.535 2.565 -9.805 2.895 ;
      RECT -10.865 3.685 -10.135 4.015 ;
    LAYER via2 ;
      RECT -0.56 2.07 -0.36 2.27 ;
      RECT -1.52 3.75 -1.32 3.95 ;
      RECT -2.52 3.75 -2.32 3.95 ;
      RECT -4.48 3.75 -4.28 3.95 ;
      RECT -5.68 3.19 -5.48 3.39 ;
      RECT -6.92 2.63 -6.72 2.83 ;
      RECT -8.36 3.19 -8.16 3.39 ;
      RECT -9.1 2.63 -8.9 2.83 ;
      RECT -10.32 2.63 -10.12 2.83 ;
      RECT -10.8 3.75 -10.6 3.95 ;
    LAYER met2 ;
      RECT 2.705 6.28 3.025 6.605 ;
      RECT 2.735 5.695 2.905 6.605 ;
      RECT 2.735 5.695 2.91 6.045 ;
      RECT 2.735 5.695 3.71 5.87 ;
      RECT 3.535 1.965 3.71 5.87 ;
      RECT -9.13 2.59 -8.935 3.375 ;
      RECT -9.105 1.47 -8.935 3.375 ;
      RECT -9.195 3.115 -9.135 3.375 ;
      RECT -7.825 2.635 -7.565 2.895 ;
      RECT -9.14 2.59 -8.935 2.87 ;
      RECT -7.83 2.645 -7.565 2.83 ;
      RECT -8.115 2.62 -8.105 2.77 ;
      RECT 3.48 1.965 3.83 2.315 ;
      RECT 1.195 2.025 3.83 2.195 ;
      RECT 1.195 1.47 1.365 2.195 ;
      RECT -9.105 1.47 1.365 1.64 ;
      RECT -7.84 2.645 -7.83 2.829 ;
      RECT -7.85 2.644 -7.84 2.826 ;
      RECT -7.859 2.643 -7.85 2.824 ;
      RECT -7.945 2.639 -7.859 2.814 ;
      RECT -8.019 2.631 -7.945 2.796 ;
      RECT -8.105 2.624 -8.019 2.779 ;
      RECT -8.165 2.62 -8.115 2.769 ;
      RECT -8.2 2.619 -8.165 2.766 ;
      RECT -8.255 2.619 -8.2 2.768 ;
      RECT -8.29 2.619 -8.255 2.772 ;
      RECT -8.376 2.618 -8.29 2.779 ;
      RECT -8.462 2.617 -8.376 2.789 ;
      RECT -8.548 2.616 -8.462 2.8 ;
      RECT -8.634 2.616 -8.548 2.81 ;
      RECT -8.72 2.615 -8.634 2.82 ;
      RECT -8.755 2.615 -8.72 2.86 ;
      RECT -8.76 2.615 -8.755 2.903 ;
      RECT -8.785 2.615 -8.76 2.92 ;
      RECT -8.86 2.615 -8.785 2.935 ;
      RECT -8.885 2.59 -8.86 2.95 ;
      RECT -8.91 2.59 -8.885 3 ;
      RECT -8.935 2.59 -8.91 3.078 ;
      RECT -9.135 2.997 -9.13 3.375 ;
      RECT 3.505 6.655 3.83 6.98 ;
      RECT 2.39 6.745 3.83 6.915 ;
      RECT 2.39 2.395 2.55 6.915 ;
      RECT 2.705 2.365 3.025 2.685 ;
      RECT 2.39 2.395 3.025 2.565 ;
      RECT 1.65 5.84 2 6.19 ;
      RECT 1.725 2.705 1.9 6.19 ;
      RECT 1.66 2.705 2.01 3.055 ;
      RECT -4.325 4.36 1.345 4.53 ;
      RECT 1.175 3.425 1.345 4.53 ;
      RECT -4.27 3.71 -4.24 3.99 ;
      RECT -4.52 3.6 -4.5 3.99 ;
      RECT -4.565 3.6 -4.5 3.86 ;
      RECT 1.085 3.43 1.435 3.78 ;
      RECT -4.735 2.225 -4.7 2.485 ;
      RECT -4.96 2.225 -4.9 2.485 ;
      RECT -4.28 3.69 -4.27 3.99 ;
      RECT -4.285 3.65 -4.28 3.99 ;
      RECT -4.3 3.605 -4.285 3.99 ;
      RECT -4.305 3.57 -4.3 3.99 ;
      RECT -4.31 3.55 -4.305 3.99 ;
      RECT -4.325 3.508 -4.31 3.99 ;
      RECT -4.34 3.446 -4.325 4.53 ;
      RECT -4.36 3.375 -4.34 4.53 ;
      RECT -4.37 3.305 -4.36 4.53 ;
      RECT -4.415 3.245 -4.37 4.53 ;
      RECT -4.495 3.207 -4.415 4.53 ;
      RECT -4.5 3.198 -4.495 3.99 ;
      RECT -4.505 3.197 -4.5 3.57 ;
      RECT -4.515 3.196 -4.505 3.553 ;
      RECT -4.54 3.177 -4.515 3.523 ;
      RECT -4.545 3.152 -4.54 3.502 ;
      RECT -4.555 3.13 -4.545 3.493 ;
      RECT -4.56 3.101 -4.555 3.483 ;
      RECT -4.6 3.027 -4.56 3.455 ;
      RECT -4.62 2.928 -4.6 3.42 ;
      RECT -4.635 2.864 -4.62 3.403 ;
      RECT -4.665 2.788 -4.635 3.375 ;
      RECT -4.685 2.703 -4.665 3.348 ;
      RECT -4.725 2.599 -4.685 3.255 ;
      RECT -4.73 2.52 -4.725 3.163 ;
      RECT -4.735 2.503 -4.73 3.14 ;
      RECT -4.74 2.225 -4.735 3.12 ;
      RECT -4.77 2.225 -4.74 3.058 ;
      RECT -4.775 2.225 -4.77 2.99 ;
      RECT -4.785 2.225 -4.775 2.955 ;
      RECT -4.795 2.225 -4.785 2.92 ;
      RECT -4.86 2.225 -4.795 2.775 ;
      RECT -4.865 2.225 -4.86 2.645 ;
      RECT -4.895 2.225 -4.865 2.578 ;
      RECT -4.9 2.225 -4.895 2.503 ;
      RECT -0.565 2.16 -0.305 2.42 ;
      RECT -0.57 2.16 -0.305 2.368 ;
      RECT -0.575 2.16 -0.305 2.338 ;
      RECT -0.6 2.03 -0.32 2.31 ;
      RECT -1.56 3.71 -1.28 3.99 ;
      RECT -1.52 3.665 -1.255 3.925 ;
      RECT -1.53 3.7 -1.255 3.925 ;
      RECT -1.525 3.685 -1.28 3.99 ;
      RECT -1.52 3.662 -1.31 3.99 ;
      RECT -1.52 3.66 -1.325 3.99 ;
      RECT -1.48 3.65 -1.325 3.99 ;
      RECT -1.51 3.655 -1.325 3.99 ;
      RECT -1.48 3.647 -1.38 3.99 ;
      RECT -1.455 3.64 -1.38 3.99 ;
      RECT -1.475 3.642 -1.38 3.99 ;
      RECT -2.145 3.155 -1.885 3.415 ;
      RECT -2.095 3.147 -1.905 3.415 ;
      RECT -2.09 3.067 -1.905 3.415 ;
      RECT -1.97 2.455 -1.905 3.415 ;
      RECT -2.065 2.852 -1.905 3.415 ;
      RECT -1.99 2.54 -1.905 3.415 ;
      RECT -1.955 2.165 -1.819 2.893 ;
      RECT -2.01 2.662 -1.819 2.893 ;
      RECT -1.995 2.602 -1.905 3.415 ;
      RECT -1.955 2.165 -1.795 2.558 ;
      RECT -1.955 2.165 -1.785 2.455 ;
      RECT -1.965 2.165 -1.705 2.425 ;
      RECT -2.56 3.71 -2.28 3.99 ;
      RECT -2.54 3.67 -2.28 3.99 ;
      RECT -2.9 3.625 -2.795 3.885 ;
      RECT -3.045 2.115 -2.955 2.375 ;
      RECT -2.505 3.18 -2.5 3.22 ;
      RECT -2.51 3.17 -2.505 3.305 ;
      RECT -2.515 3.16 -2.51 3.398 ;
      RECT -2.525 3.14 -2.515 3.454 ;
      RECT -2.605 3.068 -2.525 3.534 ;
      RECT -2.57 3.712 -2.56 3.937 ;
      RECT -2.575 3.709 -2.57 3.932 ;
      RECT -2.59 3.706 -2.575 3.925 ;
      RECT -2.625 3.7 -2.59 3.907 ;
      RECT -2.61 3.003 -2.605 3.608 ;
      RECT -2.63 2.954 -2.61 3.623 ;
      RECT -2.64 3.687 -2.625 3.89 ;
      RECT -2.635 2.896 -2.63 3.638 ;
      RECT -2.64 2.874 -2.635 3.648 ;
      RECT -2.675 2.784 -2.64 3.885 ;
      RECT -2.69 2.662 -2.675 3.885 ;
      RECT -2.695 2.615 -2.69 3.885 ;
      RECT -2.72 2.54 -2.695 3.885 ;
      RECT -2.735 2.455 -2.72 3.885 ;
      RECT -2.74 2.402 -2.735 3.885 ;
      RECT -2.745 2.382 -2.74 3.885 ;
      RECT -2.75 2.357 -2.745 3.119 ;
      RECT -2.765 3.317 -2.745 3.885 ;
      RECT -2.755 2.335 -2.75 3.096 ;
      RECT -2.765 2.287 -2.755 3.061 ;
      RECT -2.77 2.25 -2.765 3.027 ;
      RECT -2.77 3.397 -2.765 3.885 ;
      RECT -2.785 2.227 -2.77 2.982 ;
      RECT -2.79 3.495 -2.77 3.885 ;
      RECT -2.84 2.115 -2.785 2.824 ;
      RECT -2.795 3.617 -2.79 3.885 ;
      RECT -2.855 2.115 -2.84 2.663 ;
      RECT -2.86 2.115 -2.855 2.615 ;
      RECT -2.865 2.115 -2.86 2.603 ;
      RECT -2.91 2.115 -2.865 2.54 ;
      RECT -2.935 2.115 -2.91 2.458 ;
      RECT -2.95 2.115 -2.935 2.41 ;
      RECT -2.955 2.115 -2.95 2.38 ;
      RECT -3.63 3.565 -3.585 3.825 ;
      RECT -3.725 2.1 -3.58 2.36 ;
      RECT -3.22 2.722 -3.21 2.813 ;
      RECT -3.235 2.66 -3.22 2.869 ;
      RECT -3.24 2.607 -3.235 2.915 ;
      RECT -3.29 2.554 -3.24 3.041 ;
      RECT -3.295 2.509 -3.29 3.188 ;
      RECT -3.305 2.497 -3.295 3.23 ;
      RECT -3.34 2.461 -3.305 3.335 ;
      RECT -3.345 2.429 -3.34 3.441 ;
      RECT -3.36 2.411 -3.345 3.486 ;
      RECT -3.365 2.394 -3.36 2.72 ;
      RECT -3.37 2.775 -3.36 3.543 ;
      RECT -3.375 2.38 -3.365 2.693 ;
      RECT -3.38 2.83 -3.37 3.825 ;
      RECT -3.385 2.366 -3.375 2.678 ;
      RECT -3.385 2.88 -3.38 3.825 ;
      RECT -3.4 2.343 -3.385 2.658 ;
      RECT -3.42 3.002 -3.385 3.825 ;
      RECT -3.405 2.325 -3.4 2.64 ;
      RECT -3.41 2.317 -3.405 2.63 ;
      RECT -3.44 2.285 -3.41 2.594 ;
      RECT -3.43 3.13 -3.42 3.825 ;
      RECT -3.435 3.157 -3.43 3.825 ;
      RECT -3.44 3.207 -3.435 3.825 ;
      RECT -3.45 2.251 -3.44 2.559 ;
      RECT -3.49 3.275 -3.44 3.825 ;
      RECT -3.465 2.228 -3.45 2.535 ;
      RECT -3.49 2.1 -3.465 2.498 ;
      RECT -3.495 2.1 -3.49 2.47 ;
      RECT -3.525 3.375 -3.49 3.825 ;
      RECT -3.5 2.1 -3.495 2.463 ;
      RECT -3.505 2.1 -3.5 2.453 ;
      RECT -3.52 2.1 -3.505 2.438 ;
      RECT -3.535 2.1 -3.52 2.41 ;
      RECT -3.57 3.48 -3.525 3.825 ;
      RECT -3.55 2.1 -3.535 2.383 ;
      RECT -3.58 2.1 -3.55 2.368 ;
      RECT -3.585 3.552 -3.57 3.825 ;
      RECT -3.66 2.635 -3.62 2.895 ;
      RECT -3.885 2.582 -3.88 2.84 ;
      RECT -7.93 2.06 -7.67 2.32 ;
      RECT -7.93 2.085 -7.655 2.3 ;
      RECT -5.54 1.91 -5.535 2.055 ;
      RECT -3.67 2.63 -3.66 2.895 ;
      RECT -3.69 2.622 -3.67 2.895 ;
      RECT -3.708 2.618 -3.69 2.895 ;
      RECT -3.794 2.607 -3.708 2.895 ;
      RECT -3.88 2.59 -3.794 2.895 ;
      RECT -3.935 2.577 -3.885 2.825 ;
      RECT -3.969 2.569 -3.935 2.8 ;
      RECT -4.055 2.558 -3.969 2.765 ;
      RECT -4.09 2.535 -4.055 2.73 ;
      RECT -4.1 2.497 -4.09 2.716 ;
      RECT -4.105 2.47 -4.1 2.712 ;
      RECT -4.11 2.457 -4.105 2.709 ;
      RECT -4.12 2.437 -4.11 2.705 ;
      RECT -4.125 2.412 -4.12 2.701 ;
      RECT -4.15 2.367 -4.125 2.695 ;
      RECT -4.16 2.308 -4.15 2.687 ;
      RECT -4.17 2.276 -4.16 2.678 ;
      RECT -4.19 2.228 -4.17 2.658 ;
      RECT -4.195 2.188 -4.19 2.628 ;
      RECT -4.21 2.162 -4.195 2.602 ;
      RECT -4.215 2.14 -4.21 2.578 ;
      RECT -4.23 2.112 -4.215 2.554 ;
      RECT -4.245 2.085 -4.23 2.518 ;
      RECT -4.26 2.062 -4.245 2.48 ;
      RECT -4.265 2.052 -4.26 2.455 ;
      RECT -4.275 2.045 -4.265 2.438 ;
      RECT -4.29 2.032 -4.275 2.408 ;
      RECT -4.295 2.022 -4.29 2.383 ;
      RECT -4.3 2.017 -4.295 2.37 ;
      RECT -4.31 2.01 -4.3 2.35 ;
      RECT -4.315 2.003 -4.31 2.335 ;
      RECT -4.34 1.996 -4.315 2.293 ;
      RECT -4.355 1.986 -4.34 2.243 ;
      RECT -4.365 1.981 -4.355 2.213 ;
      RECT -4.375 1.977 -4.365 2.188 ;
      RECT -4.39 1.974 -4.375 2.178 ;
      RECT -4.44 1.971 -4.39 2.163 ;
      RECT -4.46 1.969 -4.44 2.148 ;
      RECT -4.509 1.967 -4.46 2.143 ;
      RECT -4.595 1.963 -4.509 2.138 ;
      RECT -4.634 1.96 -4.595 2.134 ;
      RECT -4.72 1.956 -4.634 2.129 ;
      RECT -4.77 1.953 -4.72 2.123 ;
      RECT -4.819 1.95 -4.77 2.118 ;
      RECT -4.905 1.947 -4.819 2.113 ;
      RECT -4.909 1.945 -4.905 2.11 ;
      RECT -4.995 1.942 -4.909 2.105 ;
      RECT -5.044 1.938 -4.995 2.098 ;
      RECT -5.13 1.935 -5.044 2.093 ;
      RECT -5.154 1.932 -5.13 2.089 ;
      RECT -5.24 1.93 -5.154 2.084 ;
      RECT -5.305 1.926 -5.24 2.077 ;
      RECT -5.308 1.925 -5.305 2.074 ;
      RECT -5.394 1.922 -5.308 2.071 ;
      RECT -5.48 1.916 -5.394 2.064 ;
      RECT -5.51 1.912 -5.48 2.06 ;
      RECT -5.535 1.91 -5.51 2.058 ;
      RECT -5.59 1.907 -5.54 2.055 ;
      RECT -5.67 1.906 -5.59 2.055 ;
      RECT -5.725 1.908 -5.67 2.058 ;
      RECT -5.74 1.909 -5.725 2.062 ;
      RECT -5.795 1.917 -5.74 2.072 ;
      RECT -5.825 1.925 -5.795 2.085 ;
      RECT -5.844 1.926 -5.825 2.091 ;
      RECT -5.93 1.929 -5.844 2.096 ;
      RECT -6 1.934 -5.93 2.105 ;
      RECT -6.019 1.937 -6 2.111 ;
      RECT -6.105 1.941 -6.019 2.116 ;
      RECT -6.145 1.945 -6.105 2.123 ;
      RECT -6.154 1.947 -6.145 2.126 ;
      RECT -6.24 1.951 -6.154 2.131 ;
      RECT -6.243 1.954 -6.24 2.135 ;
      RECT -6.329 1.957 -6.243 2.139 ;
      RECT -6.415 1.963 -6.329 2.147 ;
      RECT -6.439 1.967 -6.415 2.151 ;
      RECT -6.525 1.971 -6.439 2.156 ;
      RECT -6.57 1.976 -6.525 2.163 ;
      RECT -6.65 1.981 -6.57 2.17 ;
      RECT -6.73 1.987 -6.65 2.185 ;
      RECT -6.755 1.991 -6.73 2.198 ;
      RECT -6.82 1.994 -6.755 2.21 ;
      RECT -6.875 1.999 -6.82 2.225 ;
      RECT -6.905 2.002 -6.875 2.243 ;
      RECT -6.915 2.004 -6.905 2.256 ;
      RECT -6.975 2.019 -6.915 2.266 ;
      RECT -6.99 2.036 -6.975 2.275 ;
      RECT -6.995 2.045 -6.99 2.275 ;
      RECT -7.005 2.055 -6.995 2.275 ;
      RECT -7.015 2.072 -7.005 2.275 ;
      RECT -7.035 2.082 -7.015 2.276 ;
      RECT -7.08 2.092 -7.035 2.277 ;
      RECT -7.115 2.101 -7.08 2.279 ;
      RECT -7.18 2.106 -7.115 2.281 ;
      RECT -7.26 2.107 -7.18 2.284 ;
      RECT -7.264 2.105 -7.26 2.285 ;
      RECT -7.35 2.102 -7.264 2.287 ;
      RECT -7.397 2.099 -7.35 2.289 ;
      RECT -7.483 2.095 -7.397 2.292 ;
      RECT -7.569 2.091 -7.483 2.295 ;
      RECT -7.655 2.087 -7.569 2.299 ;
      RECT -5.72 3.15 -5.44 3.43 ;
      RECT -5.68 3.13 -5.42 3.39 ;
      RECT -5.69 3.14 -5.42 3.39 ;
      RECT -5.68 3.067 -5.465 3.43 ;
      RECT -5.625 2.99 -5.47 3.43 ;
      RECT -5.62 2.775 -5.47 3.43 ;
      RECT -5.63 2.577 -5.48 2.828 ;
      RECT -5.64 2.577 -5.48 2.695 ;
      RECT -5.645 2.455 -5.485 2.598 ;
      RECT -5.66 2.455 -5.485 2.503 ;
      RECT -5.665 2.165 -5.49 2.48 ;
      RECT -5.68 2.165 -5.49 2.45 ;
      RECT -5.72 2.165 -5.46 2.425 ;
      RECT -5.81 3.635 -5.73 3.895 ;
      RECT -6.405 2.355 -6.4 2.62 ;
      RECT -6.525 2.355 -6.4 2.615 ;
      RECT -5.85 3.6 -5.81 3.895 ;
      RECT -5.895 3.522 -5.85 3.895 ;
      RECT -5.915 3.45 -5.895 3.895 ;
      RECT -5.925 3.402 -5.915 3.895 ;
      RECT -5.96 3.335 -5.925 3.895 ;
      RECT -5.99 3.235 -5.96 3.895 ;
      RECT -6.01 3.16 -5.99 3.695 ;
      RECT -6.02 3.11 -6.01 3.65 ;
      RECT -6.025 3.087 -6.02 3.623 ;
      RECT -6.03 3.072 -6.025 3.61 ;
      RECT -6.035 3.057 -6.03 3.588 ;
      RECT -6.04 3.042 -6.035 3.57 ;
      RECT -6.065 2.997 -6.04 3.525 ;
      RECT -6.075 2.945 -6.065 3.468 ;
      RECT -6.085 2.915 -6.075 3.435 ;
      RECT -6.095 2.88 -6.085 3.403 ;
      RECT -6.13 2.812 -6.095 3.335 ;
      RECT -6.135 2.751 -6.13 3.27 ;
      RECT -6.145 2.739 -6.135 3.25 ;
      RECT -6.15 2.727 -6.145 3.23 ;
      RECT -6.155 2.719 -6.15 3.218 ;
      RECT -6.16 2.711 -6.155 3.198 ;
      RECT -6.17 2.699 -6.16 3.17 ;
      RECT -6.18 2.683 -6.17 3.14 ;
      RECT -6.205 2.655 -6.18 3.078 ;
      RECT -6.215 2.626 -6.205 3.023 ;
      RECT -6.23 2.605 -6.215 2.983 ;
      RECT -6.235 2.589 -6.23 2.955 ;
      RECT -6.24 2.577 -6.235 2.945 ;
      RECT -6.245 2.572 -6.24 2.918 ;
      RECT -6.25 2.565 -6.245 2.905 ;
      RECT -6.265 2.548 -6.25 2.878 ;
      RECT -6.275 2.355 -6.265 2.838 ;
      RECT -6.285 2.355 -6.275 2.805 ;
      RECT -6.295 2.355 -6.285 2.78 ;
      RECT -6.365 2.355 -6.295 2.715 ;
      RECT -6.375 2.355 -6.365 2.663 ;
      RECT -6.39 2.355 -6.375 2.645 ;
      RECT -6.4 2.355 -6.39 2.63 ;
      RECT -6.57 3.225 -6.31 3.485 ;
      RECT -8.035 3.26 -8.03 3.467 ;
      RECT -8.4 3.15 -8.325 3.465 ;
      RECT -8.585 3.205 -8.43 3.465 ;
      RECT -8.4 3.15 -8.295 3.43 ;
      RECT -6.585 3.322 -6.57 3.483 ;
      RECT -6.61 3.33 -6.585 3.488 ;
      RECT -6.635 3.337 -6.61 3.493 ;
      RECT -6.698 3.348 -6.635 3.502 ;
      RECT -6.784 3.367 -6.698 3.519 ;
      RECT -6.87 3.389 -6.784 3.538 ;
      RECT -6.885 3.402 -6.87 3.549 ;
      RECT -6.925 3.41 -6.885 3.556 ;
      RECT -6.945 3.415 -6.925 3.563 ;
      RECT -6.983 3.416 -6.945 3.566 ;
      RECT -7.069 3.419 -6.983 3.567 ;
      RECT -7.155 3.423 -7.069 3.568 ;
      RECT -7.204 3.425 -7.155 3.57 ;
      RECT -7.29 3.425 -7.204 3.572 ;
      RECT -7.33 3.42 -7.29 3.574 ;
      RECT -7.34 3.414 -7.33 3.575 ;
      RECT -7.38 3.409 -7.34 3.572 ;
      RECT -7.39 3.402 -7.38 3.568 ;
      RECT -7.405 3.398 -7.39 3.566 ;
      RECT -7.422 3.394 -7.405 3.564 ;
      RECT -7.508 3.384 -7.422 3.556 ;
      RECT -7.594 3.366 -7.508 3.542 ;
      RECT -7.68 3.349 -7.594 3.528 ;
      RECT -7.705 3.337 -7.68 3.519 ;
      RECT -7.775 3.327 -7.705 3.512 ;
      RECT -7.82 3.315 -7.775 3.503 ;
      RECT -7.88 3.302 -7.82 3.495 ;
      RECT -7.885 3.294 -7.88 3.49 ;
      RECT -7.92 3.289 -7.885 3.488 ;
      RECT -7.975 3.28 -7.92 3.481 ;
      RECT -8.015 3.269 -7.975 3.473 ;
      RECT -8.03 3.262 -8.015 3.469 ;
      RECT -8.05 3.255 -8.035 3.466 ;
      RECT -8.065 3.245 -8.05 3.464 ;
      RECT -8.08 3.232 -8.065 3.461 ;
      RECT -8.105 3.215 -8.08 3.457 ;
      RECT -8.12 3.197 -8.105 3.454 ;
      RECT -8.145 3.15 -8.12 3.452 ;
      RECT -8.169 3.15 -8.145 3.449 ;
      RECT -8.255 3.15 -8.169 3.441 ;
      RECT -8.295 3.15 -8.255 3.433 ;
      RECT -8.43 3.197 -8.4 3.465 ;
      RECT -6.75 2.78 -6.49 3.04 ;
      RECT -6.79 2.78 -6.49 2.918 ;
      RECT -6.825 2.78 -6.49 2.903 ;
      RECT -6.88 2.78 -6.49 2.883 ;
      RECT -6.96 2.59 -6.68 2.87 ;
      RECT -6.96 2.772 -6.61 2.87 ;
      RECT -6.96 2.715 -6.625 2.87 ;
      RECT -6.96 2.662 -6.675 2.87 ;
      RECT -9.8 2.949 -9.785 3.405 ;
      RECT -9.805 3.021 -9.699 3.403 ;
      RECT -9.785 2.115 -9.65 3.401 ;
      RECT -9.8 2.965 -9.645 3.4 ;
      RECT -9.8 3.015 -9.64 3.398 ;
      RECT -9.815 3.08 -9.64 3.397 ;
      RECT -9.805 3.072 -9.635 3.394 ;
      RECT -9.825 3.12 -9.635 3.389 ;
      RECT -9.825 3.12 -9.62 3.386 ;
      RECT -9.83 3.12 -9.62 3.383 ;
      RECT -9.855 3.12 -9.595 3.38 ;
      RECT -9.785 2.115 -9.625 2.768 ;
      RECT -9.79 2.115 -9.625 2.74 ;
      RECT -9.795 2.115 -9.625 2.568 ;
      RECT -9.795 2.115 -9.605 2.508 ;
      RECT -9.84 2.115 -9.58 2.375 ;
      RECT -10.36 2.59 -10.08 2.87 ;
      RECT -10.37 2.605 -10.08 2.865 ;
      RECT -10.415 2.667 -10.08 2.863 ;
      RECT -10.34 2.582 -10.175 2.87 ;
      RECT -10.34 2.567 -10.219 2.87 ;
      RECT -10.305 2.56 -10.219 2.87 ;
      RECT -10.84 3.71 -10.56 3.99 ;
      RECT -10.88 3.672 -10.585 3.783 ;
      RECT -10.895 3.622 -10.605 3.678 ;
      RECT -10.95 3.385 -10.69 3.645 ;
      RECT -10.95 3.587 -10.61 3.645 ;
      RECT -10.95 3.527 -10.615 3.645 ;
      RECT -10.95 3.477 -10.635 3.645 ;
      RECT -10.95 3.457 -10.64 3.645 ;
      RECT -10.95 3.435 -10.645 3.645 ;
      RECT -10.95 3.42 -10.675 3.645 ;
    LAYER via1 ;
      RECT 3.595 6.74 3.745 6.89 ;
      RECT 3.58 2.065 3.73 2.215 ;
      RECT 2.79 2.45 2.94 2.6 ;
      RECT 2.79 6.37 2.94 6.52 ;
      RECT 1.76 2.805 1.91 2.955 ;
      RECT 1.75 5.94 1.9 6.09 ;
      RECT 1.185 3.53 1.335 3.68 ;
      RECT -0.51 2.215 -0.36 2.365 ;
      RECT -1.46 3.72 -1.31 3.87 ;
      RECT -1.91 2.22 -1.76 2.37 ;
      RECT -2.09 3.21 -1.94 3.36 ;
      RECT -2.485 3.725 -2.335 3.875 ;
      RECT -2.845 3.68 -2.695 3.83 ;
      RECT -2.99 2.17 -2.84 2.32 ;
      RECT -3.575 3.62 -3.425 3.77 ;
      RECT -3.67 2.155 -3.52 2.305 ;
      RECT -3.825 2.69 -3.675 2.84 ;
      RECT -4.51 3.655 -4.36 3.805 ;
      RECT -4.905 2.28 -4.755 2.43 ;
      RECT -5.625 3.185 -5.475 3.335 ;
      RECT -5.665 2.22 -5.515 2.37 ;
      RECT -5.935 3.69 -5.785 3.84 ;
      RECT -6.47 2.41 -6.32 2.56 ;
      RECT -6.515 3.28 -6.365 3.43 ;
      RECT -6.695 2.835 -6.545 2.985 ;
      RECT -7.77 2.69 -7.62 2.84 ;
      RECT -7.875 2.115 -7.725 2.265 ;
      RECT -8.53 3.26 -8.38 3.41 ;
      RECT -9.14 3.17 -8.99 3.32 ;
      RECT -9.785 2.17 -9.635 2.32 ;
      RECT -9.8 3.175 -9.65 3.325 ;
      RECT -10.315 2.66 -10.165 2.81 ;
      RECT -10.895 3.44 -10.745 3.59 ;
    LAYER met1 ;
      RECT -11.115 0 0.845 1.89 ;
      RECT -11.12 0 0.845 1.68 ;
      RECT -11.49 0 6.435 0.305 ;
      RECT -11.49 4.285 6.435 4.745 ;
      RECT -11.115 4.135 6.435 4.745 ;
      RECT -11.115 4.13 0.845 4.745 ;
      RECT 5.835 2.365 6.125 2.595 ;
      RECT 5.895 0.885 6.065 2.595 ;
      RECT 5.835 0.885 6.125 1.115 ;
      RECT 5.835 7.765 6.125 7.995 ;
      RECT 5.895 6.285 6.065 7.995 ;
      RECT 5.835 6.285 6.125 6.515 ;
      RECT 5.425 2.735 5.755 2.965 ;
      RECT 5.425 2.765 5.925 2.935 ;
      RECT 5.425 2.395 5.615 2.965 ;
      RECT 4.845 2.365 5.135 2.595 ;
      RECT 4.845 2.395 5.615 2.565 ;
      RECT 4.905 0.885 5.075 2.595 ;
      RECT 4.845 0.885 5.135 1.115 ;
      RECT 4.845 7.765 5.135 7.995 ;
      RECT 4.905 6.285 5.075 7.995 ;
      RECT 4.845 6.285 5.135 6.515 ;
      RECT 4.845 6.325 5.695 6.485 ;
      RECT 5.525 5.915 5.695 6.485 ;
      RECT 4.845 6.32 5.235 6.485 ;
      RECT 5.465 5.915 5.755 6.145 ;
      RECT 5.465 5.945 5.925 6.115 ;
      RECT 4.475 2.735 4.765 2.965 ;
      RECT 4.475 2.765 4.935 2.935 ;
      RECT 4.535 1.655 4.7 2.965 ;
      RECT 3.05 1.625 3.34 1.855 ;
      RECT 3.05 1.655 4.7 1.825 ;
      RECT 3.11 0.885 3.28 1.855 ;
      RECT 3.05 0.885 3.34 1.115 ;
      RECT 3.05 7.765 3.34 7.995 ;
      RECT 3.11 7.025 3.28 7.995 ;
      RECT 3.11 7.12 4.7 7.29 ;
      RECT 4.53 5.915 4.7 7.29 ;
      RECT 3.05 7.025 3.34 7.255 ;
      RECT 4.475 5.915 4.765 6.145 ;
      RECT 4.475 5.945 4.935 6.115 ;
      RECT 3.48 1.965 3.83 2.315 ;
      RECT 3.31 2.025 3.83 2.195 ;
      RECT 3.505 6.655 3.83 6.98 ;
      RECT 3.48 6.655 3.83 6.885 ;
      RECT 3.31 6.685 3.83 6.855 ;
      RECT 1.085 3.43 1.435 3.78 ;
      RECT 1.175 2.395 1.345 3.78 ;
      RECT 2.705 2.365 3.025 2.685 ;
      RECT 2.675 2.365 3.025 2.595 ;
      RECT 1.175 2.395 3.025 2.565 ;
      RECT 2.705 6.28 3.025 6.605 ;
      RECT 2.675 6.285 3.025 6.515 ;
      RECT 2.505 6.315 3.025 6.485 ;
      RECT 1.66 2.705 2.01 3.055 ;
      RECT 1.66 2.765 2.14 2.935 ;
      RECT 1.65 5.84 2 6.19 ;
      RECT 1.65 5.945 2.14 6.115 ;
      RECT -1.515 3.665 -1.475 3.925 ;
      RECT -1.475 3.645 -1.47 3.655 ;
      RECT -0.135 2.735 0.02 3.055 ;
      RECT -0.215 2.735 -0.135 3.22 ;
      RECT -0.225 2.735 -0.215 3.363 ;
      RECT -0.25 2.735 -0.225 3.41 ;
      RECT -0.275 2.735 -0.25 3.488 ;
      RECT -0.295 2.735 -0.275 3.558 ;
      RECT -0.3 2.735 -0.295 3.588 ;
      RECT -0.32 2.885 -0.3 3.6 ;
      RECT -0.33 2.885 -0.32 3.618 ;
      RECT -0.34 2.887 -0.33 3.626 ;
      RECT -0.345 2.892 -0.34 3.083 ;
      RECT -0.345 3.092 -0.34 3.627 ;
      RECT -0.35 3.137 -0.345 3.628 ;
      RECT -0.36 3.202 -0.35 3.629 ;
      RECT -0.37 3.297 -0.36 3.631 ;
      RECT -0.375 3.35 -0.37 3.633 ;
      RECT -0.38 3.37 -0.375 3.634 ;
      RECT -0.435 3.395 -0.38 3.64 ;
      RECT -0.475 3.43 -0.435 3.649 ;
      RECT -0.485 3.447 -0.475 3.654 ;
      RECT -0.494 3.453 -0.485 3.656 ;
      RECT -0.58 3.491 -0.494 3.667 ;
      RECT -0.585 3.53 -0.58 3.677 ;
      RECT -0.66 3.537 -0.585 3.687 ;
      RECT -0.68 3.547 -0.66 3.698 ;
      RECT -0.71 3.554 -0.68 3.706 ;
      RECT -0.735 3.561 -0.71 3.713 ;
      RECT -0.759 3.567 -0.735 3.718 ;
      RECT -0.845 3.58 -0.759 3.73 ;
      RECT -0.923 3.587 -0.845 3.748 ;
      RECT -1.009 3.582 -0.923 3.766 ;
      RECT -1.095 3.577 -1.009 3.786 ;
      RECT -1.175 3.571 -1.095 3.803 ;
      RECT -1.24 3.567 -1.175 3.832 ;
      RECT -1.245 3.281 -1.24 3.305 ;
      RECT -1.255 3.557 -1.24 3.86 ;
      RECT -1.25 3.275 -1.245 3.345 ;
      RECT -1.255 3.269 -1.25 3.415 ;
      RECT -1.26 3.263 -1.255 3.493 ;
      RECT -1.26 3.54 -1.255 3.925 ;
      RECT -1.268 3.26 -1.26 3.925 ;
      RECT -1.354 3.258 -1.268 3.925 ;
      RECT -1.44 3.256 -1.354 3.925 ;
      RECT -1.45 3.257 -1.44 3.925 ;
      RECT -1.455 3.262 -1.45 3.925 ;
      RECT -1.465 3.275 -1.455 3.925 ;
      RECT -1.47 3.297 -1.465 3.925 ;
      RECT -1.475 3.657 -1.47 3.925 ;
      RECT -0.845 3.125 -0.84 3.345 ;
      RECT -0.34 2.16 -0.305 2.42 ;
      RECT -0.355 2.16 -0.34 2.428 ;
      RECT -0.384 2.16 -0.355 2.45 ;
      RECT -0.47 2.16 -0.384 2.51 ;
      RECT -0.49 2.16 -0.47 2.575 ;
      RECT -0.55 2.16 -0.49 2.74 ;
      RECT -0.555 2.16 -0.55 2.888 ;
      RECT -0.56 2.16 -0.555 2.9 ;
      RECT -0.565 2.16 -0.56 2.926 ;
      RECT -0.595 2.346 -0.565 3.006 ;
      RECT -0.6 2.394 -0.595 3.095 ;
      RECT -0.605 2.408 -0.6 3.11 ;
      RECT -0.61 2.427 -0.605 3.14 ;
      RECT -0.615 2.442 -0.61 3.156 ;
      RECT -0.62 2.457 -0.615 3.178 ;
      RECT -0.625 2.477 -0.62 3.2 ;
      RECT -0.635 2.497 -0.625 3.233 ;
      RECT -0.65 2.539 -0.635 3.295 ;
      RECT -0.655 2.57 -0.65 3.335 ;
      RECT -0.66 2.582 -0.655 3.34 ;
      RECT -0.665 2.594 -0.66 3.345 ;
      RECT -0.67 2.607 -0.665 3.345 ;
      RECT -0.675 2.625 -0.67 3.345 ;
      RECT -0.68 2.645 -0.675 3.345 ;
      RECT -0.685 2.657 -0.68 3.345 ;
      RECT -0.69 2.67 -0.685 3.345 ;
      RECT -0.71 2.705 -0.69 3.345 ;
      RECT -0.76 2.807 -0.71 3.345 ;
      RECT -0.765 2.892 -0.76 3.345 ;
      RECT -0.77 2.9 -0.765 3.345 ;
      RECT -0.775 2.917 -0.77 3.345 ;
      RECT -0.78 2.932 -0.775 3.345 ;
      RECT -0.815 2.997 -0.78 3.345 ;
      RECT -0.83 3.062 -0.815 3.345 ;
      RECT -0.835 3.092 -0.83 3.345 ;
      RECT -0.84 3.117 -0.835 3.345 ;
      RECT -0.855 3.127 -0.845 3.345 ;
      RECT -0.87 3.14 -0.855 3.338 ;
      RECT -1.125 2.73 -1.055 2.94 ;
      RECT -1.335 2.707 -1.33 2.9 ;
      RECT -3.88 2.635 -3.62 2.895 ;
      RECT -1.045 2.917 -1.04 2.92 ;
      RECT -1.055 2.735 -1.045 2.935 ;
      RECT -1.154 2.728 -1.125 2.94 ;
      RECT -1.24 2.72 -1.154 2.94 ;
      RECT -1.255 2.714 -1.24 2.938 ;
      RECT -1.275 2.713 -1.255 2.925 ;
      RECT -1.28 2.712 -1.275 2.908 ;
      RECT -1.33 2.709 -1.28 2.903 ;
      RECT -1.36 2.706 -1.335 2.898 ;
      RECT -1.38 2.704 -1.36 2.893 ;
      RECT -1.395 2.702 -1.38 2.89 ;
      RECT -1.425 2.7 -1.395 2.888 ;
      RECT -1.49 2.696 -1.425 2.88 ;
      RECT -1.52 2.691 -1.49 2.875 ;
      RECT -1.54 2.689 -1.52 2.873 ;
      RECT -1.57 2.686 -1.54 2.868 ;
      RECT -1.63 2.682 -1.57 2.86 ;
      RECT -1.635 2.679 -1.63 2.855 ;
      RECT -1.705 2.677 -1.635 2.85 ;
      RECT -1.734 2.673 -1.705 2.843 ;
      RECT -1.82 2.668 -1.734 2.835 ;
      RECT -1.854 2.663 -1.82 2.827 ;
      RECT -1.94 2.655 -1.854 2.819 ;
      RECT -1.979 2.648 -1.94 2.811 ;
      RECT -2.065 2.643 -1.979 2.803 ;
      RECT -2.13 2.637 -2.065 2.793 ;
      RECT -2.15 2.632 -2.13 2.788 ;
      RECT -2.159 2.629 -2.15 2.787 ;
      RECT -2.245 2.625 -2.159 2.781 ;
      RECT -2.285 2.621 -2.245 2.773 ;
      RECT -2.305 2.617 -2.285 2.771 ;
      RECT -2.365 2.617 -2.305 2.768 ;
      RECT -2.385 2.62 -2.365 2.766 ;
      RECT -2.406 2.62 -2.385 2.766 ;
      RECT -2.492 2.622 -2.406 2.77 ;
      RECT -2.578 2.624 -2.492 2.776 ;
      RECT -2.664 2.626 -2.578 2.783 ;
      RECT -2.75 2.629 -2.664 2.789 ;
      RECT -2.784 2.63 -2.75 2.794 ;
      RECT -2.87 2.633 -2.784 2.799 ;
      RECT -2.899 2.64 -2.87 2.804 ;
      RECT -2.985 2.64 -2.899 2.809 ;
      RECT -3.018 2.64 -2.985 2.814 ;
      RECT -3.104 2.642 -3.018 2.819 ;
      RECT -3.19 2.644 -3.104 2.826 ;
      RECT -3.254 2.646 -3.19 2.832 ;
      RECT -3.34 2.648 -3.254 2.838 ;
      RECT -3.343 2.65 -3.34 2.841 ;
      RECT -3.429 2.651 -3.343 2.845 ;
      RECT -3.515 2.654 -3.429 2.852 ;
      RECT -3.534 2.656 -3.515 2.856 ;
      RECT -3.62 2.658 -3.534 2.861 ;
      RECT -3.89 2.67 -3.88 2.865 ;
      RECT -1.655 2.25 -1.47 2.46 ;
      RECT -1.66 2.251 -1.465 2.458 ;
      RECT -1.665 2.256 -1.455 2.453 ;
      RECT -1.67 2.232 -1.665 2.45 ;
      RECT -1.7 2.229 -1.67 2.443 ;
      RECT -1.705 2.225 -1.7 2.434 ;
      RECT -1.74 2.256 -1.455 2.429 ;
      RECT -1.965 2.165 -1.705 2.425 ;
      RECT -1.665 2.234 -1.66 2.453 ;
      RECT -1.66 2.235 -1.655 2.458 ;
      RECT -1.965 2.247 -1.585 2.425 ;
      RECT -1.965 2.245 -1.6 2.425 ;
      RECT -1.965 2.24 -1.61 2.425 ;
      RECT -2.01 3.155 -1.96 3.44 ;
      RECT -2.065 3.125 -2.06 3.44 ;
      RECT -2.095 3.105 -2.09 3.44 ;
      RECT -1.945 3.155 -1.885 3.415 ;
      RECT -1.95 3.155 -1.945 3.423 ;
      RECT -1.96 3.155 -1.95 3.435 ;
      RECT -2.045 3.145 -2.01 3.44 ;
      RECT -2.05 3.132 -2.045 3.44 ;
      RECT -2.06 3.127 -2.05 3.44 ;
      RECT -2.08 3.117 -2.065 3.44 ;
      RECT -2.09 3.11 -2.08 3.44 ;
      RECT -2.1 3.102 -2.095 3.44 ;
      RECT -2.13 3.092 -2.1 3.44 ;
      RECT -2.145 3.08 -2.13 3.44 ;
      RECT -2.16 3.07 -2.145 3.435 ;
      RECT -2.18 3.06 -2.16 3.41 ;
      RECT -2.19 3.052 -2.18 3.387 ;
      RECT -2.22 3.035 -2.19 3.377 ;
      RECT -2.225 3.012 -2.22 3.368 ;
      RECT -2.23 2.999 -2.225 3.366 ;
      RECT -2.245 2.975 -2.23 3.36 ;
      RECT -2.25 2.951 -2.245 3.354 ;
      RECT -2.26 2.94 -2.25 3.349 ;
      RECT -2.265 2.93 -2.26 3.345 ;
      RECT -2.27 2.922 -2.265 3.342 ;
      RECT -2.28 2.917 -2.27 3.338 ;
      RECT -2.285 2.912 -2.28 3.334 ;
      RECT -2.37 2.91 -2.285 3.309 ;
      RECT -2.4 2.91 -2.37 3.275 ;
      RECT -2.415 2.91 -2.4 3.258 ;
      RECT -2.47 2.91 -2.415 3.203 ;
      RECT -2.475 2.915 -2.47 3.152 ;
      RECT -2.485 2.92 -2.475 3.142 ;
      RECT -2.49 2.93 -2.485 3.128 ;
      RECT -2.54 3.67 -2.28 3.93 ;
      RECT -2.62 3.685 -2.28 3.906 ;
      RECT -2.64 3.685 -2.28 3.901 ;
      RECT -2.664 3.685 -2.28 3.899 ;
      RECT -2.75 3.685 -2.28 3.894 ;
      RECT -2.9 3.625 -2.64 3.89 ;
      RECT -2.945 3.685 -2.28 3.885 ;
      RECT -2.95 3.692 -2.28 3.88 ;
      RECT -2.935 3.68 -2.62 3.89 ;
      RECT -3.045 2.115 -2.785 2.375 ;
      RECT -3.045 2.172 -2.78 2.368 ;
      RECT -3.045 2.202 -2.775 2.3 ;
      RECT -2.985 2.633 -2.87 2.635 ;
      RECT -2.899 2.63 -2.87 2.635 ;
      RECT -3.875 3.634 -3.85 3.874 ;
      RECT -3.89 3.637 -3.8 3.868 ;
      RECT -3.895 3.642 -3.714 3.863 ;
      RECT -3.9 3.65 -3.65 3.861 ;
      RECT -3.9 3.65 -3.64 3.86 ;
      RECT -3.905 3.657 -3.63 3.853 ;
      RECT -3.905 3.657 -3.544 3.842 ;
      RECT -3.91 3.692 -3.544 3.838 ;
      RECT -3.91 3.692 -3.535 3.827 ;
      RECT -3.63 3.565 -3.37 3.825 ;
      RECT -3.92 3.742 -3.37 3.823 ;
      RECT -3.65 3.61 -3.63 3.858 ;
      RECT -3.714 3.613 -3.65 3.862 ;
      RECT -3.8 3.618 -3.714 3.867 ;
      RECT -3.87 3.629 -3.37 3.825 ;
      RECT -3.85 3.623 -3.8 3.872 ;
      RECT -3.725 2.1 -3.715 2.362 ;
      RECT -3.735 2.157 -3.725 2.365 ;
      RECT -3.76 2.162 -3.735 2.371 ;
      RECT -3.785 2.166 -3.76 2.383 ;
      RECT -3.795 2.169 -3.785 2.393 ;
      RECT -3.8 2.17 -3.795 2.398 ;
      RECT -3.805 2.171 -3.8 2.403 ;
      RECT -3.81 2.172 -3.805 2.405 ;
      RECT -3.835 2.175 -3.81 2.408 ;
      RECT -3.865 2.181 -3.835 2.411 ;
      RECT -3.93 2.192 -3.865 2.414 ;
      RECT -3.975 2.2 -3.93 2.418 ;
      RECT -3.99 2.2 -3.975 2.426 ;
      RECT -3.995 2.201 -3.99 2.433 ;
      RECT -4 2.203 -3.995 2.436 ;
      RECT -4.005 2.207 -4 2.439 ;
      RECT -4.015 2.215 -4.005 2.443 ;
      RECT -4.02 2.228 -4.015 2.448 ;
      RECT -4.025 2.236 -4.02 2.45 ;
      RECT -4.03 2.242 -4.025 2.45 ;
      RECT -4.035 2.246 -4.03 2.453 ;
      RECT -4.04 2.248 -4.035 2.456 ;
      RECT -4.045 2.251 -4.04 2.459 ;
      RECT -4.055 2.256 -4.045 2.463 ;
      RECT -4.06 2.262 -4.055 2.468 ;
      RECT -4.07 2.268 -4.06 2.472 ;
      RECT -4.085 2.275 -4.07 2.478 ;
      RECT -4.114 2.289 -4.085 2.488 ;
      RECT -4.2 2.324 -4.114 2.52 ;
      RECT -4.22 2.357 -4.2 2.549 ;
      RECT -4.24 2.37 -4.22 2.56 ;
      RECT -4.26 2.382 -4.24 2.571 ;
      RECT -4.31 2.404 -4.26 2.591 ;
      RECT -4.325 2.422 -4.31 2.608 ;
      RECT -4.33 2.428 -4.325 2.611 ;
      RECT -4.335 2.432 -4.33 2.614 ;
      RECT -4.34 2.436 -4.335 2.618 ;
      RECT -4.345 2.438 -4.34 2.621 ;
      RECT -4.355 2.445 -4.345 2.624 ;
      RECT -4.36 2.45 -4.355 2.628 ;
      RECT -4.365 2.452 -4.36 2.631 ;
      RECT -4.37 2.456 -4.365 2.634 ;
      RECT -4.375 2.458 -4.37 2.638 ;
      RECT -4.39 2.463 -4.375 2.643 ;
      RECT -4.395 2.468 -4.39 2.646 ;
      RECT -4.4 2.476 -4.395 2.649 ;
      RECT -4.405 2.478 -4.4 2.652 ;
      RECT -4.41 2.48 -4.405 2.655 ;
      RECT -4.42 2.482 -4.41 2.661 ;
      RECT -4.455 2.496 -4.42 2.673 ;
      RECT -4.465 2.511 -4.455 2.683 ;
      RECT -4.54 2.54 -4.465 2.707 ;
      RECT -4.545 2.565 -4.54 2.73 ;
      RECT -4.56 2.569 -4.545 2.736 ;
      RECT -4.57 2.577 -4.56 2.741 ;
      RECT -4.6 2.59 -4.57 2.745 ;
      RECT -4.61 2.605 -4.6 2.75 ;
      RECT -4.62 2.61 -4.61 2.753 ;
      RECT -4.625 2.612 -4.62 2.755 ;
      RECT -4.64 2.615 -4.625 2.758 ;
      RECT -4.645 2.617 -4.64 2.761 ;
      RECT -4.665 2.622 -4.645 2.765 ;
      RECT -4.695 2.627 -4.665 2.773 ;
      RECT -4.72 2.634 -4.695 2.781 ;
      RECT -4.725 2.639 -4.72 2.786 ;
      RECT -4.755 2.642 -4.725 2.79 ;
      RECT -4.795 2.645 -4.755 2.8 ;
      RECT -4.83 2.642 -4.795 2.812 ;
      RECT -4.84 2.638 -4.83 2.819 ;
      RECT -4.865 2.634 -4.84 2.825 ;
      RECT -4.87 2.63 -4.865 2.83 ;
      RECT -4.91 2.627 -4.87 2.83 ;
      RECT -4.925 2.612 -4.91 2.831 ;
      RECT -4.948 2.6 -4.925 2.831 ;
      RECT -5.034 2.6 -4.948 2.832 ;
      RECT -5.12 2.6 -5.034 2.834 ;
      RECT -5.14 2.6 -5.12 2.831 ;
      RECT -5.145 2.605 -5.14 2.826 ;
      RECT -5.15 2.61 -5.145 2.824 ;
      RECT -5.16 2.62 -5.15 2.822 ;
      RECT -5.165 2.626 -5.16 2.815 ;
      RECT -5.17 2.628 -5.165 2.8 ;
      RECT -5.175 2.632 -5.17 2.79 ;
      RECT -3.715 2.1 -3.465 2.36 ;
      RECT -5.99 3.635 -5.73 3.895 ;
      RECT -3.695 3.125 -3.69 3.335 ;
      RECT -3.69 3.13 -3.68 3.33 ;
      RECT -3.74 3.125 -3.695 3.35 ;
      RECT -3.75 3.125 -3.74 3.37 ;
      RECT -3.769 3.125 -3.75 3.375 ;
      RECT -3.855 3.125 -3.769 3.372 ;
      RECT -3.885 3.127 -3.855 3.37 ;
      RECT -3.94 3.137 -3.885 3.368 ;
      RECT -4.005 3.151 -3.94 3.366 ;
      RECT -4.01 3.159 -4.005 3.365 ;
      RECT -4.025 3.162 -4.01 3.363 ;
      RECT -4.09 3.172 -4.025 3.359 ;
      RECT -4.138 3.186 -4.09 3.36 ;
      RECT -4.224 3.203 -4.138 3.374 ;
      RECT -4.31 3.224 -4.224 3.391 ;
      RECT -4.33 3.237 -4.31 3.401 ;
      RECT -4.375 3.245 -4.33 3.408 ;
      RECT -4.41 3.253 -4.375 3.416 ;
      RECT -4.444 3.261 -4.41 3.424 ;
      RECT -4.53 3.275 -4.444 3.436 ;
      RECT -4.565 3.292 -4.53 3.448 ;
      RECT -4.574 3.301 -4.565 3.452 ;
      RECT -4.66 3.319 -4.574 3.469 ;
      RECT -4.719 3.346 -4.66 3.496 ;
      RECT -4.805 3.373 -4.719 3.524 ;
      RECT -4.825 3.395 -4.805 3.544 ;
      RECT -4.885 3.41 -4.825 3.56 ;
      RECT -4.895 3.422 -4.885 3.573 ;
      RECT -4.9 3.427 -4.895 3.576 ;
      RECT -4.91 3.43 -4.9 3.579 ;
      RECT -4.915 3.432 -4.91 3.582 ;
      RECT -4.945 3.44 -4.915 3.589 ;
      RECT -4.96 3.447 -4.945 3.597 ;
      RECT -4.97 3.452 -4.96 3.601 ;
      RECT -4.975 3.455 -4.97 3.604 ;
      RECT -4.985 3.457 -4.975 3.607 ;
      RECT -5.02 3.467 -4.985 3.616 ;
      RECT -5.095 3.49 -5.02 3.638 ;
      RECT -5.115 3.508 -5.095 3.656 ;
      RECT -5.145 3.515 -5.115 3.666 ;
      RECT -5.165 3.523 -5.145 3.676 ;
      RECT -5.175 3.529 -5.165 3.683 ;
      RECT -5.194 3.534 -5.175 3.689 ;
      RECT -5.28 3.554 -5.194 3.709 ;
      RECT -5.295 3.574 -5.28 3.728 ;
      RECT -5.34 3.586 -5.295 3.739 ;
      RECT -5.405 3.607 -5.34 3.762 ;
      RECT -5.445 3.627 -5.405 3.783 ;
      RECT -5.455 3.637 -5.445 3.793 ;
      RECT -5.505 3.649 -5.455 3.804 ;
      RECT -5.525 3.665 -5.505 3.816 ;
      RECT -5.555 3.675 -5.525 3.822 ;
      RECT -5.565 3.68 -5.555 3.824 ;
      RECT -5.634 3.681 -5.565 3.83 ;
      RECT -5.72 3.683 -5.634 3.84 ;
      RECT -5.73 3.684 -5.72 3.845 ;
      RECT -4.46 3.71 -4.27 3.92 ;
      RECT -4.47 3.715 -4.26 3.913 ;
      RECT -4.485 3.715 -4.26 3.878 ;
      RECT -4.565 3.6 -4.305 3.86 ;
      RECT -5.65 3.13 -5.465 3.425 ;
      RECT -5.66 3.13 -5.465 3.423 ;
      RECT -5.675 3.13 -5.46 3.418 ;
      RECT -5.675 3.13 -5.455 3.415 ;
      RECT -5.68 3.13 -5.455 3.413 ;
      RECT -5.685 3.385 -5.455 3.403 ;
      RECT -5.68 3.13 -5.42 3.39 ;
      RECT -5.72 2.165 -5.46 2.425 ;
      RECT -5.91 2.09 -5.824 2.423 ;
      RECT -5.935 2.094 -5.78 2.419 ;
      RECT -5.824 2.086 -5.78 2.419 ;
      RECT -5.824 2.087 -5.775 2.418 ;
      RECT -5.91 2.092 -5.76 2.417 ;
      RECT -5.935 2.1 -5.72 2.416 ;
      RECT -5.94 2.095 -5.76 2.411 ;
      RECT -5.95 2.11 -5.72 2.318 ;
      RECT -5.95 2.162 -5.52 2.318 ;
      RECT -5.95 2.155 -5.54 2.318 ;
      RECT -5.95 2.142 -5.57 2.318 ;
      RECT -5.95 2.13 -5.63 2.318 ;
      RECT -5.95 2.115 -5.655 2.318 ;
      RECT -6.75 2.745 -6.615 3.04 ;
      RECT -6.49 2.768 -6.485 2.955 ;
      RECT -5.77 2.665 -5.625 2.9 ;
      RECT -5.61 2.665 -5.605 2.89 ;
      RECT -5.575 2.676 -5.57 2.87 ;
      RECT -5.58 2.668 -5.575 2.875 ;
      RECT -5.6 2.665 -5.58 2.88 ;
      RECT -5.605 2.665 -5.6 2.888 ;
      RECT -5.615 2.665 -5.61 2.893 ;
      RECT -5.625 2.665 -5.615 2.898 ;
      RECT -5.795 2.667 -5.77 2.9 ;
      RECT -5.845 2.674 -5.795 2.9 ;
      RECT -5.85 2.679 -5.845 2.9 ;
      RECT -5.889 2.684 -5.85 2.901 ;
      RECT -5.975 2.696 -5.889 2.902 ;
      RECT -5.984 2.706 -5.975 2.902 ;
      RECT -6.07 2.715 -5.984 2.904 ;
      RECT -6.094 2.725 -6.07 2.906 ;
      RECT -6.18 2.736 -6.094 2.907 ;
      RECT -6.21 2.747 -6.18 2.909 ;
      RECT -6.24 2.752 -6.21 2.911 ;
      RECT -6.265 2.758 -6.24 2.914 ;
      RECT -6.28 2.763 -6.265 2.915 ;
      RECT -6.325 2.769 -6.28 2.915 ;
      RECT -6.33 2.774 -6.325 2.916 ;
      RECT -6.35 2.774 -6.33 2.918 ;
      RECT -6.37 2.772 -6.35 2.923 ;
      RECT -6.405 2.771 -6.37 2.93 ;
      RECT -6.435 2.77 -6.405 2.94 ;
      RECT -6.485 2.769 -6.435 2.95 ;
      RECT -6.575 2.766 -6.49 3.04 ;
      RECT -6.6 2.76 -6.575 3.04 ;
      RECT -6.615 2.75 -6.6 3.04 ;
      RECT -6.8 2.745 -6.75 2.96 ;
      RECT -6.81 2.75 -6.8 2.95 ;
      RECT -6.57 3.225 -6.31 3.485 ;
      RECT -6.57 3.225 -6.28 3.378 ;
      RECT -6.57 3.225 -6.245 3.363 ;
      RECT -6.315 3.145 -6.125 3.355 ;
      RECT -6.325 3.15 -6.115 3.348 ;
      RECT -6.36 3.22 -6.115 3.348 ;
      RECT -6.33 3.162 -6.31 3.485 ;
      RECT -6.345 3.21 -6.115 3.348 ;
      RECT -6.34 3.182 -6.31 3.485 ;
      RECT -7.26 2.25 -7.19 3.355 ;
      RECT -6.525 2.355 -6.265 2.615 ;
      RECT -6.945 2.401 -6.93 2.61 ;
      RECT -6.609 2.414 -6.525 2.565 ;
      RECT -6.695 2.411 -6.609 2.565 ;
      RECT -6.734 2.409 -6.695 2.565 ;
      RECT -6.82 2.407 -6.734 2.565 ;
      RECT -6.88 2.405 -6.82 2.576 ;
      RECT -6.915 2.403 -6.88 2.594 ;
      RECT -6.93 2.401 -6.915 2.605 ;
      RECT -6.96 2.401 -6.945 2.618 ;
      RECT -6.97 2.401 -6.96 2.623 ;
      RECT -6.995 2.4 -6.97 2.628 ;
      RECT -7.01 2.395 -6.995 2.634 ;
      RECT -7.015 2.388 -7.01 2.639 ;
      RECT -7.04 2.379 -7.015 2.645 ;
      RECT -7.085 2.358 -7.04 2.658 ;
      RECT -7.095 2.342 -7.085 2.668 ;
      RECT -7.11 2.335 -7.095 2.678 ;
      RECT -7.12 2.328 -7.11 2.695 ;
      RECT -7.125 2.325 -7.12 2.725 ;
      RECT -7.13 2.323 -7.125 2.755 ;
      RECT -7.135 2.321 -7.13 2.792 ;
      RECT -7.15 2.317 -7.135 2.859 ;
      RECT -7.15 3.15 -7.14 3.35 ;
      RECT -7.155 2.313 -7.15 2.985 ;
      RECT -7.155 3.137 -7.15 3.355 ;
      RECT -7.16 2.311 -7.155 3.07 ;
      RECT -7.16 3.127 -7.155 3.355 ;
      RECT -7.175 2.282 -7.16 3.355 ;
      RECT -7.19 2.255 -7.175 3.355 ;
      RECT -7.265 2.25 -7.26 2.605 ;
      RECT -7.265 2.66 -7.26 3.355 ;
      RECT -7.28 2.25 -7.265 2.583 ;
      RECT -7.27 2.682 -7.265 3.355 ;
      RECT -7.28 2.722 -7.27 3.355 ;
      RECT -7.315 2.25 -7.28 2.525 ;
      RECT -7.285 2.757 -7.28 3.355 ;
      RECT -7.3 2.812 -7.285 3.355 ;
      RECT -7.305 2.877 -7.3 3.355 ;
      RECT -7.32 2.925 -7.305 3.355 ;
      RECT -7.345 2.25 -7.315 2.48 ;
      RECT -7.325 2.98 -7.32 3.355 ;
      RECT -7.34 3.04 -7.325 3.355 ;
      RECT -7.345 3.088 -7.34 3.353 ;
      RECT -7.35 2.25 -7.345 2.473 ;
      RECT -7.35 3.12 -7.345 3.348 ;
      RECT -7.375 2.25 -7.35 2.465 ;
      RECT -7.385 2.255 -7.375 2.455 ;
      RECT -7.17 3.53 -7.15 3.77 ;
      RECT -7.94 3.46 -7.935 3.67 ;
      RECT -6.66 3.533 -6.65 3.728 ;
      RECT -6.665 3.523 -6.66 3.731 ;
      RECT -6.745 3.52 -6.665 3.754 ;
      RECT -6.749 3.52 -6.745 3.776 ;
      RECT -6.835 3.52 -6.749 3.786 ;
      RECT -6.85 3.52 -6.835 3.794 ;
      RECT -6.879 3.521 -6.85 3.792 ;
      RECT -6.965 3.526 -6.879 3.788 ;
      RECT -6.978 3.53 -6.965 3.784 ;
      RECT -7.064 3.53 -6.978 3.78 ;
      RECT -7.15 3.53 -7.064 3.774 ;
      RECT -7.234 3.53 -7.17 3.768 ;
      RECT -7.32 3.53 -7.234 3.763 ;
      RECT -7.34 3.53 -7.32 3.759 ;
      RECT -7.4 3.525 -7.34 3.756 ;
      RECT -7.428 3.519 -7.4 3.753 ;
      RECT -7.514 3.514 -7.428 3.749 ;
      RECT -7.6 3.508 -7.514 3.743 ;
      RECT -7.675 3.49 -7.6 3.738 ;
      RECT -7.71 3.467 -7.675 3.734 ;
      RECT -7.72 3.457 -7.71 3.733 ;
      RECT -7.775 3.455 -7.72 3.732 ;
      RECT -7.85 3.455 -7.775 3.728 ;
      RECT -7.86 3.455 -7.85 3.723 ;
      RECT -7.875 3.455 -7.86 3.715 ;
      RECT -7.925 3.457 -7.875 3.693 ;
      RECT -7.935 3.46 -7.925 3.673 ;
      RECT -7.945 3.465 -7.94 3.668 ;
      RECT -7.95 3.47 -7.945 3.663 ;
      RECT -7.825 2.635 -7.565 2.895 ;
      RECT -7.825 2.65 -7.545 2.86 ;
      RECT -7.825 2.655 -7.535 2.855 ;
      RECT -9.84 2.115 -9.58 2.375 ;
      RECT -9.85 2.145 -9.58 2.355 ;
      RECT -7.93 2.06 -7.67 2.32 ;
      RECT -7.935 2.135 -7.93 2.321 ;
      RECT -7.96 2.14 -7.935 2.323 ;
      RECT -7.975 2.147 -7.96 2.326 ;
      RECT -8.035 2.165 -7.975 2.331 ;
      RECT -8.065 2.185 -8.035 2.338 ;
      RECT -8.09 2.193 -8.065 2.343 ;
      RECT -8.115 2.201 -8.09 2.345 ;
      RECT -8.133 2.205 -8.115 2.344 ;
      RECT -8.219 2.203 -8.133 2.344 ;
      RECT -8.305 2.201 -8.219 2.344 ;
      RECT -8.391 2.199 -8.305 2.343 ;
      RECT -8.477 2.197 -8.391 2.343 ;
      RECT -8.563 2.195 -8.477 2.343 ;
      RECT -8.649 2.193 -8.563 2.343 ;
      RECT -8.735 2.191 -8.649 2.342 ;
      RECT -8.753 2.19 -8.735 2.342 ;
      RECT -8.839 2.189 -8.753 2.342 ;
      RECT -8.925 2.187 -8.839 2.342 ;
      RECT -9.011 2.186 -8.925 2.341 ;
      RECT -9.097 2.185 -9.011 2.341 ;
      RECT -9.183 2.183 -9.097 2.341 ;
      RECT -9.269 2.182 -9.183 2.341 ;
      RECT -9.355 2.18 -9.269 2.34 ;
      RECT -9.379 2.178 -9.355 2.34 ;
      RECT -9.465 2.171 -9.379 2.34 ;
      RECT -9.494 2.163 -9.465 2.34 ;
      RECT -9.58 2.155 -9.494 2.34 ;
      RECT -9.86 2.152 -9.85 2.35 ;
      RECT -8.355 3.115 -8.35 3.465 ;
      RECT -8.585 3.205 -8.445 3.465 ;
      RECT -8.11 2.89 -8.065 3.1 ;
      RECT -8.055 2.901 -8.045 3.095 ;
      RECT -8.065 2.893 -8.055 3.1 ;
      RECT -8.13 2.89 -8.11 3.105 ;
      RECT -8.16 2.89 -8.13 3.128 ;
      RECT -8.17 2.89 -8.16 3.153 ;
      RECT -8.175 2.89 -8.17 3.163 ;
      RECT -8.23 2.89 -8.175 3.203 ;
      RECT -8.235 2.89 -8.23 3.243 ;
      RECT -8.24 2.892 -8.235 3.248 ;
      RECT -8.255 2.902 -8.24 3.259 ;
      RECT -8.3 2.96 -8.255 3.295 ;
      RECT -8.31 3.015 -8.3 3.329 ;
      RECT -8.325 3.042 -8.31 3.345 ;
      RECT -8.335 3.069 -8.325 3.465 ;
      RECT -8.35 3.092 -8.335 3.465 ;
      RECT -8.36 3.132 -8.355 3.465 ;
      RECT -8.365 3.142 -8.36 3.465 ;
      RECT -8.37 3.157 -8.365 3.465 ;
      RECT -8.38 3.162 -8.37 3.465 ;
      RECT -8.445 3.185 -8.38 3.465 ;
      RECT -8.945 2.68 -8.755 2.89 ;
      RECT -10.37 2.605 -10.11 2.865 ;
      RECT -10.02 2.6 -9.925 2.81 ;
      RECT -10.045 2.615 -10.035 2.81 ;
      RECT -8.755 2.687 -8.745 2.885 ;
      RECT -8.955 2.687 -8.945 2.885 ;
      RECT -8.97 2.702 -8.955 2.875 ;
      RECT -8.975 2.71 -8.97 2.868 ;
      RECT -8.985 2.713 -8.975 2.865 ;
      RECT -9.02 2.712 -8.985 2.863 ;
      RECT -9.049 2.708 -9.02 2.86 ;
      RECT -9.135 2.703 -9.049 2.857 ;
      RECT -9.195 2.697 -9.135 2.853 ;
      RECT -9.224 2.693 -9.195 2.85 ;
      RECT -9.31 2.685 -9.224 2.847 ;
      RECT -9.319 2.679 -9.31 2.845 ;
      RECT -9.405 2.674 -9.319 2.843 ;
      RECT -9.428 2.669 -9.405 2.84 ;
      RECT -9.514 2.663 -9.428 2.837 ;
      RECT -9.6 2.654 -9.514 2.832 ;
      RECT -9.61 2.649 -9.6 2.83 ;
      RECT -9.629 2.648 -9.61 2.829 ;
      RECT -9.715 2.643 -9.629 2.825 ;
      RECT -9.735 2.638 -9.715 2.821 ;
      RECT -9.795 2.633 -9.735 2.818 ;
      RECT -9.82 2.623 -9.795 2.816 ;
      RECT -9.825 2.616 -9.82 2.815 ;
      RECT -9.835 2.607 -9.825 2.814 ;
      RECT -9.839 2.6 -9.835 2.814 ;
      RECT -9.925 2.6 -9.839 2.812 ;
      RECT -10.035 2.607 -10.02 2.81 ;
      RECT -10.05 2.617 -10.045 2.81 ;
      RECT -10.07 2.62 -10.05 2.807 ;
      RECT -10.1 2.62 -10.07 2.803 ;
      RECT -10.11 2.62 -10.1 2.803 ;
      RECT -9.195 3.115 -8.935 3.375 ;
      RECT -9.265 3.125 -8.935 3.335 ;
      RECT -9.275 3.132 -8.935 3.33 ;
      RECT -9.855 3.12 -9.595 3.38 ;
      RECT -9.855 3.16 -9.49 3.37 ;
      RECT -9.855 3.162 -9.485 3.369 ;
      RECT -9.855 3.17 -9.48 3.366 ;
      RECT -10.93 2.245 -10.83 3.77 ;
      RECT -10.74 3.385 -10.69 3.645 ;
      RECT -10.745 2.258 -10.74 2.445 ;
      RECT -10.75 3.366 -10.74 3.645 ;
      RECT -10.75 2.255 -10.745 2.453 ;
      RECT -10.765 2.249 -10.75 2.46 ;
      RECT -10.755 3.354 -10.75 3.728 ;
      RECT -10.765 3.342 -10.755 3.765 ;
      RECT -10.775 2.245 -10.765 2.467 ;
      RECT -10.775 3.327 -10.765 3.77 ;
      RECT -10.78 2.245 -10.775 2.475 ;
      RECT -10.8 3.297 -10.775 3.77 ;
      RECT -10.82 2.245 -10.78 2.523 ;
      RECT -10.81 3.257 -10.8 3.77 ;
      RECT -10.82 3.212 -10.81 3.77 ;
      RECT -10.825 2.245 -10.82 2.593 ;
      RECT -10.825 3.17 -10.82 3.77 ;
      RECT -10.83 2.245 -10.825 3.07 ;
      RECT -10.83 3.152 -10.825 3.77 ;
      RECT -10.94 2.248 -10.93 3.77 ;
      RECT -10.955 2.255 -10.94 3.766 ;
      RECT -10.96 2.265 -10.955 3.761 ;
      RECT -10.965 2.465 -10.96 3.653 ;
      RECT -10.97 2.55 -10.965 3.205 ;
      RECT -11.485 8.575 6.435 8.88 ;
      RECT -4.96 2.225 -4.7 2.485 ;
    LAYER mcon ;
      RECT 5.895 0.915 6.065 1.085 ;
      RECT 5.895 2.395 6.065 2.565 ;
      RECT 5.895 6.315 6.065 6.485 ;
      RECT 5.895 7.795 6.065 7.965 ;
      RECT 5.545 0.105 5.715 0.275 ;
      RECT 5.545 4.165 5.715 4.335 ;
      RECT 5.545 4.545 5.715 4.715 ;
      RECT 5.545 8.605 5.715 8.775 ;
      RECT 5.525 2.765 5.695 2.935 ;
      RECT 5.525 5.945 5.695 6.115 ;
      RECT 4.905 0.915 5.075 1.085 ;
      RECT 4.905 2.395 5.075 2.565 ;
      RECT 4.905 6.315 5.075 6.485 ;
      RECT 4.905 7.795 5.075 7.965 ;
      RECT 4.555 0.105 4.725 0.275 ;
      RECT 4.555 4.165 4.725 4.335 ;
      RECT 4.555 4.545 4.725 4.715 ;
      RECT 4.555 8.605 4.725 8.775 ;
      RECT 4.535 2.765 4.705 2.935 ;
      RECT 4.535 5.945 4.705 6.115 ;
      RECT 3.85 0.105 4.02 0.275 ;
      RECT 3.85 4.165 4.02 4.335 ;
      RECT 3.85 4.545 4.02 4.715 ;
      RECT 3.85 8.605 4.02 8.775 ;
      RECT 3.54 2.025 3.71 2.195 ;
      RECT 3.54 6.685 3.71 6.855 ;
      RECT 3.17 0.105 3.34 0.275 ;
      RECT 3.17 8.605 3.34 8.775 ;
      RECT 3.11 0.915 3.28 1.085 ;
      RECT 3.11 1.655 3.28 1.825 ;
      RECT 3.11 7.055 3.28 7.225 ;
      RECT 3.11 7.795 3.28 7.965 ;
      RECT 2.735 2.395 2.905 2.565 ;
      RECT 2.735 6.315 2.905 6.485 ;
      RECT 2.49 0.105 2.66 0.275 ;
      RECT 2.49 8.605 2.66 8.775 ;
      RECT 1.81 0.105 1.98 0.275 ;
      RECT 1.81 8.605 1.98 8.775 ;
      RECT 1.74 2.765 1.91 2.935 ;
      RECT 1.74 5.945 1.91 6.115 ;
      RECT 0.53 1.565 0.7 1.735 ;
      RECT 0.53 4.285 0.7 4.455 ;
      RECT 0.07 1.565 0.24 1.735 ;
      RECT 0.07 4.285 0.24 4.455 ;
      RECT -0.325 2.905 -0.155 3.075 ;
      RECT -0.39 1.565 -0.22 1.735 ;
      RECT -0.39 4.285 -0.22 4.455 ;
      RECT -0.535 2.245 -0.365 2.415 ;
      RECT -0.85 1.565 -0.68 1.735 ;
      RECT -0.85 3.155 -0.68 3.325 ;
      RECT -0.85 4.285 -0.68 4.455 ;
      RECT -1.235 2.75 -1.065 2.92 ;
      RECT -1.31 1.565 -1.14 1.735 ;
      RECT -1.31 4.285 -1.14 4.455 ;
      RECT -1.45 3.315 -1.28 3.485 ;
      RECT -1.47 3.715 -1.3 3.885 ;
      RECT -1.645 2.27 -1.475 2.44 ;
      RECT -1.77 1.565 -1.6 1.735 ;
      RECT -1.77 4.285 -1.6 4.455 ;
      RECT -2.14 3.25 -1.97 3.42 ;
      RECT -2.23 1.565 -2.06 1.735 ;
      RECT -2.23 4.285 -2.06 4.455 ;
      RECT -2.465 2.935 -2.295 3.105 ;
      RECT -2.53 3.715 -2.36 3.885 ;
      RECT -2.69 1.565 -2.52 1.735 ;
      RECT -2.69 4.285 -2.52 4.455 ;
      RECT -2.93 3.7 -2.76 3.87 ;
      RECT -2.97 2.185 -2.8 2.355 ;
      RECT -3.15 1.565 -2.98 1.735 ;
      RECT -3.15 4.285 -2.98 4.455 ;
      RECT -3.61 1.565 -3.44 1.735 ;
      RECT -3.61 4.285 -3.44 4.455 ;
      RECT -3.87 2.685 -3.7 2.855 ;
      RECT -3.87 3.145 -3.7 3.315 ;
      RECT -3.87 3.66 -3.7 3.83 ;
      RECT -3.985 2.22 -3.815 2.39 ;
      RECT -4.07 1.565 -3.9 1.735 ;
      RECT -4.07 4.285 -3.9 4.455 ;
      RECT -4.45 3.73 -4.28 3.9 ;
      RECT -4.53 1.565 -4.36 1.735 ;
      RECT -4.53 4.285 -4.36 4.455 ;
      RECT -4.93 2.26 -4.76 2.43 ;
      RECT -4.99 1.565 -4.82 1.735 ;
      RECT -4.99 4.285 -4.82 4.455 ;
      RECT -5.145 2.635 -4.975 2.805 ;
      RECT -5.45 1.565 -5.28 1.735 ;
      RECT -5.45 4.285 -5.28 4.455 ;
      RECT -5.645 3.235 -5.475 3.405 ;
      RECT -5.76 2.685 -5.59 2.855 ;
      RECT -5.91 1.565 -5.74 1.735 ;
      RECT -5.91 4.285 -5.74 4.455 ;
      RECT -5.93 2.135 -5.76 2.305 ;
      RECT -6.305 3.165 -6.135 3.335 ;
      RECT -6.37 1.565 -6.2 1.735 ;
      RECT -6.37 4.285 -6.2 4.455 ;
      RECT -6.79 2.765 -6.62 2.935 ;
      RECT -6.83 1.565 -6.66 1.735 ;
      RECT -6.83 4.285 -6.66 4.455 ;
      RECT -6.84 3.54 -6.67 3.71 ;
      RECT -7.29 1.565 -7.12 1.735 ;
      RECT -7.29 4.285 -7.12 4.455 ;
      RECT -7.33 3.165 -7.16 3.335 ;
      RECT -7.365 2.27 -7.195 2.44 ;
      RECT -7.725 2.67 -7.555 2.84 ;
      RECT -7.75 1.565 -7.58 1.735 ;
      RECT -7.75 4.285 -7.58 4.455 ;
      RECT -7.93 3.48 -7.76 3.65 ;
      RECT -8.21 1.565 -8.04 1.735 ;
      RECT -8.21 4.285 -8.04 4.455 ;
      RECT -8.235 2.91 -8.065 3.08 ;
      RECT -8.67 1.565 -8.5 1.735 ;
      RECT -8.67 4.285 -8.5 4.455 ;
      RECT -8.935 2.7 -8.765 2.87 ;
      RECT -9.13 1.565 -8.96 1.735 ;
      RECT -9.13 4.285 -8.96 4.455 ;
      RECT -9.255 3.145 -9.085 3.315 ;
      RECT -9.59 1.565 -9.42 1.735 ;
      RECT -9.59 4.285 -9.42 4.455 ;
      RECT -9.67 3.18 -9.5 3.35 ;
      RECT -9.84 2.165 -9.67 2.335 ;
      RECT -10.015 2.62 -9.845 2.79 ;
      RECT -10.05 1.565 -9.88 1.735 ;
      RECT -10.05 4.285 -9.88 4.455 ;
      RECT -10.51 1.565 -10.34 1.735 ;
      RECT -10.51 4.285 -10.34 4.455 ;
      RECT -10.935 2.27 -10.765 2.44 ;
      RECT -10.94 3.585 -10.77 3.755 ;
      RECT -10.97 1.565 -10.8 1.735 ;
      RECT -10.97 4.285 -10.8 4.455 ;
    LAYER li ;
      RECT -0.065 0 0.105 2.235 ;
      RECT -1.025 0 -0.855 2.235 ;
      RECT -1.985 0 -1.815 2.235 ;
      RECT -2.505 0 -2.335 2.235 ;
      RECT -3.465 0 -3.295 2.235 ;
      RECT -4.465 0 -4.295 2.235 ;
      RECT -5.425 0 -5.255 2.235 ;
      RECT -6.905 0 -6.735 2.235 ;
      RECT -8.825 0 -8.655 2.235 ;
      RECT -10.305 0 -10.135 2.235 ;
      RECT -11.115 0 0.845 1.735 ;
      RECT -11.12 0 0.845 1.68 ;
      RECT 5.465 0 5.635 0.935 ;
      RECT 4.475 0 4.645 0.935 ;
      RECT 1.73 0 1.9 0.935 ;
      RECT -11.49 0 6.435 0.305 ;
      RECT 5.465 3.405 5.635 5.475 ;
      RECT 4.475 3.405 4.645 5.475 ;
      RECT 1.73 3.405 1.9 5.475 ;
      RECT -11.49 4.285 6.435 4.745 ;
      RECT 0.475 4.135 6.435 4.745 ;
      RECT -1.025 3.785 -0.855 4.745 ;
      RECT -3.465 3.785 -3.295 4.745 ;
      RECT -5.425 3.785 -5.255 4.745 ;
      RECT -6.385 3.785 -6.215 4.745 ;
      RECT -8.345 3.785 -8.175 4.745 ;
      RECT -9.345 3.785 -9.175 4.745 ;
      RECT -10.305 3.785 -10.135 4.745 ;
      RECT -11.485 8.575 6.435 8.88 ;
      RECT 5.465 7.945 5.635 8.88 ;
      RECT 4.475 7.945 4.645 8.88 ;
      RECT 1.73 7.945 1.9 8.88 ;
      RECT 5.525 1.74 5.695 2.935 ;
      RECT 5.525 1.74 5.99 1.91 ;
      RECT 5.525 6.97 5.99 7.14 ;
      RECT 5.525 5.945 5.695 7.14 ;
      RECT 4.535 1.74 4.705 2.935 ;
      RECT 4.535 1.74 5 1.91 ;
      RECT 4.535 6.97 5 7.14 ;
      RECT 4.535 5.945 4.705 7.14 ;
      RECT 2.68 2.635 2.85 3.865 ;
      RECT 2.735 0.855 2.905 2.805 ;
      RECT 2.68 0.575 2.85 1.025 ;
      RECT 2.68 7.855 2.85 8.305 ;
      RECT 2.735 6.075 2.905 8.025 ;
      RECT 2.68 5.015 2.85 6.245 ;
      RECT 2.16 0.575 2.33 3.865 ;
      RECT 2.16 2.075 2.565 2.405 ;
      RECT 2.16 1.235 2.565 1.565 ;
      RECT 2.16 5.015 2.33 8.305 ;
      RECT 2.16 7.315 2.565 7.645 ;
      RECT 2.16 6.475 2.565 6.805 ;
      RECT 0.26 3.392 0.275 3.443 ;
      RECT 0.255 3.372 0.26 3.49 ;
      RECT 0.24 3.362 0.255 3.558 ;
      RECT 0.215 3.342 0.24 3.613 ;
      RECT 0.175 3.327 0.215 3.633 ;
      RECT 0.13 3.321 0.175 3.661 ;
      RECT 0.06 3.311 0.13 3.678 ;
      RECT 0.04 3.303 0.06 3.678 ;
      RECT -0.02 3.297 0.04 3.67 ;
      RECT -0.079 3.288 -0.02 3.658 ;
      RECT -0.165 3.277 -0.079 3.641 ;
      RECT -0.187 3.268 -0.165 3.629 ;
      RECT -0.273 3.261 -0.187 3.616 ;
      RECT -0.359 3.248 -0.273 3.597 ;
      RECT -0.445 3.236 -0.359 3.577 ;
      RECT -0.475 3.225 -0.445 3.564 ;
      RECT -0.525 3.211 -0.475 3.556 ;
      RECT -0.545 3.2 -0.525 3.548 ;
      RECT -0.594 3.189 -0.545 3.54 ;
      RECT -0.68 3.168 -0.594 3.525 ;
      RECT -0.725 3.155 -0.68 3.51 ;
      RECT -0.77 3.155 -0.725 3.49 ;
      RECT -0.825 3.155 -0.77 3.425 ;
      RECT -0.85 3.155 -0.825 3.348 ;
      RECT -0.325 2.892 -0.155 3.075 ;
      RECT -0.325 2.892 -0.14 3.033 ;
      RECT -0.325 2.892 -0.135 2.975 ;
      RECT -0.265 2.66 -0.13 2.951 ;
      RECT -0.265 2.664 -0.125 2.934 ;
      RECT -0.32 2.827 -0.125 2.934 ;
      RECT -0.295 2.672 -0.155 3.075 ;
      RECT -0.295 2.676 -0.115 2.875 ;
      RECT -0.31 2.762 -0.115 2.875 ;
      RECT -0.3 2.692 -0.155 3.075 ;
      RECT -0.3 2.695 -0.105 2.788 ;
      RECT -0.305 2.712 -0.105 2.788 ;
      RECT -0.535 1.932 -0.365 2.415 ;
      RECT -0.54 1.927 -0.39 2.405 ;
      RECT -0.54 1.934 -0.36 2.399 ;
      RECT -0.55 1.928 -0.39 2.378 ;
      RECT -0.55 1.944 -0.345 2.337 ;
      RECT -0.58 1.929 -0.39 2.3 ;
      RECT -0.58 1.959 -0.335 2.24 ;
      RECT -0.585 1.931 -0.39 2.238 ;
      RECT -0.605 1.94 -0.36 2.195 ;
      RECT -0.63 1.956 -0.345 2.107 ;
      RECT -0.63 1.975 -0.32 2.098 ;
      RECT -0.635 2.012 -0.32 2.05 ;
      RECT -0.63 1.992 -0.315 2.018 ;
      RECT -0.535 1.926 -0.425 2.415 ;
      RECT -0.449 1.925 -0.425 2.415 ;
      RECT -1.215 2.71 -1.21 2.921 ;
      RECT -0.615 2.71 -0.61 2.895 ;
      RECT -0.55 2.75 -0.545 2.863 ;
      RECT -0.555 2.742 -0.55 2.869 ;
      RECT -0.56 2.732 -0.555 2.877 ;
      RECT -0.565 2.722 -0.56 2.886 ;
      RECT -0.57 2.712 -0.565 2.89 ;
      RECT -0.61 2.71 -0.57 2.893 ;
      RECT -0.638 2.709 -0.615 2.897 ;
      RECT -0.724 2.706 -0.638 2.904 ;
      RECT -0.81 2.702 -0.724 2.915 ;
      RECT -0.83 2.7 -0.81 2.921 ;
      RECT -0.848 2.699 -0.83 2.924 ;
      RECT -0.934 2.697 -0.848 2.931 ;
      RECT -1.02 2.692 -0.934 2.944 ;
      RECT -1.039 2.689 -1.02 2.949 ;
      RECT -1.125 2.687 -1.039 2.94 ;
      RECT -1.135 2.687 -1.125 2.933 ;
      RECT -1.21 2.7 -1.135 2.927 ;
      RECT -1.225 2.711 -1.215 2.921 ;
      RECT -1.235 2.713 -1.225 2.92 ;
      RECT -1.245 2.717 -1.235 2.916 ;
      RECT -1.25 2.72 -1.245 2.91 ;
      RECT -1.26 2.722 -1.25 2.904 ;
      RECT -1.265 2.725 -1.26 2.898 ;
      RECT -1.285 3.311 -1.28 3.515 ;
      RECT -1.3 3.298 -1.285 3.608 ;
      RECT -1.315 3.279 -1.3 3.885 ;
      RECT -1.35 3.245 -1.315 3.885 ;
      RECT -1.354 3.215 -1.35 3.885 ;
      RECT -1.44 3.097 -1.354 3.885 ;
      RECT -1.45 2.972 -1.44 3.885 ;
      RECT -1.465 2.94 -1.45 3.885 ;
      RECT -1.47 2.915 -1.465 3.885 ;
      RECT -1.475 2.905 -1.47 3.841 ;
      RECT -1.49 2.877 -1.475 3.746 ;
      RECT -1.505 2.843 -1.49 3.645 ;
      RECT -1.51 2.821 -1.505 3.598 ;
      RECT -1.515 2.81 -1.51 3.568 ;
      RECT -1.52 2.8 -1.515 3.534 ;
      RECT -1.53 2.787 -1.52 3.502 ;
      RECT -1.555 2.763 -1.53 3.428 ;
      RECT -1.56 2.743 -1.555 3.353 ;
      RECT -1.565 2.737 -1.56 3.328 ;
      RECT -1.57 2.732 -1.565 3.293 ;
      RECT -1.575 2.727 -1.57 3.268 ;
      RECT -1.58 2.725 -1.575 3.248 ;
      RECT -1.585 2.725 -1.58 3.233 ;
      RECT -1.59 2.725 -1.585 3.193 ;
      RECT -1.6 2.725 -1.59 3.165 ;
      RECT -1.61 2.725 -1.6 3.11 ;
      RECT -1.625 2.725 -1.61 3.048 ;
      RECT -1.63 2.724 -1.625 2.993 ;
      RECT -1.645 2.723 -1.63 2.973 ;
      RECT -1.705 2.721 -1.645 2.947 ;
      RECT -1.74 2.722 -1.705 2.927 ;
      RECT -1.745 2.724 -1.74 2.917 ;
      RECT -1.755 2.743 -1.745 2.907 ;
      RECT -1.76 2.77 -1.755 2.838 ;
      RECT -1.645 2.195 -1.475 2.44 ;
      RECT -1.61 1.966 -1.475 2.44 ;
      RECT -1.61 1.968 -1.465 2.435 ;
      RECT -1.61 1.97 -1.44 2.423 ;
      RECT -1.61 1.973 -1.415 2.405 ;
      RECT -1.61 1.978 -1.365 2.378 ;
      RECT -1.61 1.983 -1.345 2.343 ;
      RECT -1.63 1.985 -1.335 2.318 ;
      RECT -1.64 2.08 -1.335 2.318 ;
      RECT -1.61 1.965 -1.5 2.44 ;
      RECT -1.6 1.962 -1.505 2.44 ;
      RECT -2.08 3.227 -1.89 3.585 ;
      RECT -2.08 3.239 -1.855 3.584 ;
      RECT -2.08 3.267 -1.835 3.582 ;
      RECT -2.08 3.292 -1.83 3.581 ;
      RECT -2.08 3.35 -1.815 3.58 ;
      RECT -2.095 3.223 -1.935 3.565 ;
      RECT -2.115 3.232 -1.89 3.518 ;
      RECT -2.14 3.243 -1.855 3.455 ;
      RECT -2.14 3.327 -1.82 3.455 ;
      RECT -2.14 3.302 -1.825 3.455 ;
      RECT -2.08 3.218 -1.935 3.585 ;
      RECT -1.994 3.217 -1.935 3.585 ;
      RECT -1.994 3.216 -1.95 3.585 ;
      RECT -2.295 2.732 -2.29 3.11 ;
      RECT -2.3 2.7 -2.295 3.11 ;
      RECT -2.305 2.672 -2.3 3.11 ;
      RECT -2.31 2.652 -2.305 3.11 ;
      RECT -2.365 2.635 -2.31 3.11 ;
      RECT -2.405 2.62 -2.365 3.11 ;
      RECT -2.46 2.607 -2.405 3.11 ;
      RECT -2.495 2.598 -2.46 3.11 ;
      RECT -2.499 2.596 -2.495 3.109 ;
      RECT -2.585 2.592 -2.499 3.092 ;
      RECT -2.67 2.584 -2.585 3.055 ;
      RECT -2.68 2.58 -2.67 3.028 ;
      RECT -2.69 2.58 -2.68 3.01 ;
      RECT -2.7 2.582 -2.69 2.993 ;
      RECT -2.705 2.587 -2.7 2.979 ;
      RECT -2.71 2.591 -2.705 2.966 ;
      RECT -2.72 2.596 -2.71 2.95 ;
      RECT -2.735 2.61 -2.72 2.925 ;
      RECT -2.74 2.616 -2.735 2.905 ;
      RECT -2.745 2.618 -2.74 2.898 ;
      RECT -2.75 2.622 -2.745 2.773 ;
      RECT -2.57 3.422 -2.325 3.885 ;
      RECT -2.65 3.395 -2.33 3.881 ;
      RECT -2.72 3.43 -2.325 3.874 ;
      RECT -2.93 3.685 -2.325 3.87 ;
      RECT -2.75 3.453 -2.325 3.87 ;
      RECT -2.91 3.645 -2.325 3.87 ;
      RECT -2.76 3.465 -2.325 3.87 ;
      RECT -2.875 3.582 -2.325 3.87 ;
      RECT -2.82 3.507 -2.325 3.87 ;
      RECT -2.57 3.372 -2.33 3.885 ;
      RECT -2.54 3.365 -2.33 3.885 ;
      RECT -2.55 3.367 -2.33 3.885 ;
      RECT -2.54 3.362 -2.41 3.885 ;
      RECT -2.985 1.925 -2.899 2.364 ;
      RECT -2.99 1.925 -2.899 2.362 ;
      RECT -2.99 1.925 -2.83 2.361 ;
      RECT -2.99 1.925 -2.8 2.358 ;
      RECT -3.005 1.932 -2.8 2.349 ;
      RECT -3.005 1.932 -2.795 2.345 ;
      RECT -3.01 1.942 -2.795 2.338 ;
      RECT -3.015 1.947 -2.795 2.313 ;
      RECT -3.015 1.947 -2.78 2.295 ;
      RECT -2.99 1.925 -2.76 2.21 ;
      RECT -3.02 1.952 -2.76 2.208 ;
      RECT -3.01 1.945 -2.755 2.146 ;
      RECT -3.02 2.067 -2.75 2.129 ;
      RECT -3.035 1.962 -2.755 2.08 ;
      RECT -3.04 1.972 -2.755 1.98 ;
      RECT -2.96 2.743 -2.955 2.82 ;
      RECT -2.97 2.737 -2.96 3.01 ;
      RECT -2.98 2.729 -2.97 3.031 ;
      RECT -2.99 2.72 -2.98 3.053 ;
      RECT -2.995 2.715 -2.99 3.07 ;
      RECT -3.035 2.715 -2.995 3.11 ;
      RECT -3.055 2.715 -3.035 3.165 ;
      RECT -3.06 2.715 -3.055 3.193 ;
      RECT -3.07 2.715 -3.06 3.208 ;
      RECT -3.105 2.715 -3.07 3.25 ;
      RECT -3.11 2.715 -3.105 3.293 ;
      RECT -3.12 2.715 -3.11 3.308 ;
      RECT -3.135 2.715 -3.12 3.328 ;
      RECT -3.15 2.715 -3.135 3.355 ;
      RECT -3.155 2.716 -3.15 3.373 ;
      RECT -3.175 2.717 -3.155 3.38 ;
      RECT -3.23 2.718 -3.175 3.4 ;
      RECT -3.24 2.719 -3.23 3.414 ;
      RECT -3.245 2.722 -3.24 3.413 ;
      RECT -3.285 2.795 -3.245 3.411 ;
      RECT -3.3 2.875 -3.285 3.409 ;
      RECT -3.325 2.93 -3.3 3.407 ;
      RECT -3.34 2.995 -3.325 3.406 ;
      RECT -3.385 3.027 -3.34 3.403 ;
      RECT -3.47 3.05 -3.385 3.398 ;
      RECT -3.495 3.07 -3.47 3.393 ;
      RECT -3.565 3.075 -3.495 3.389 ;
      RECT -3.585 3.077 -3.565 3.386 ;
      RECT -3.67 3.088 -3.585 3.38 ;
      RECT -3.675 3.099 -3.67 3.375 ;
      RECT -3.685 3.101 -3.675 3.375 ;
      RECT -3.72 3.105 -3.685 3.373 ;
      RECT -3.77 3.115 -3.72 3.36 ;
      RECT -3.79 3.123 -3.77 3.345 ;
      RECT -3.87 3.135 -3.79 3.328 ;
      RECT -3.705 2.685 -3.535 2.895 ;
      RECT -3.589 2.681 -3.535 2.895 ;
      RECT -3.784 2.685 -3.535 2.886 ;
      RECT -3.784 2.685 -3.53 2.875 ;
      RECT -3.87 2.685 -3.53 2.866 ;
      RECT -3.87 2.693 -3.52 2.81 ;
      RECT -3.87 2.705 -3.515 2.723 ;
      RECT -3.87 2.712 -3.51 2.715 ;
      RECT -3.675 2.683 -3.535 2.895 ;
      RECT -3.92 3.628 -3.675 3.96 ;
      RECT -3.925 3.62 -3.92 3.957 ;
      RECT -3.955 3.64 -3.675 3.938 ;
      RECT -3.975 3.672 -3.675 3.911 ;
      RECT -3.925 3.625 -3.748 3.957 ;
      RECT -3.925 3.622 -3.834 3.957 ;
      RECT -3.985 1.97 -3.815 2.39 ;
      RECT -3.99 1.97 -3.815 2.388 ;
      RECT -3.99 1.97 -3.79 2.378 ;
      RECT -3.99 1.97 -3.77 2.353 ;
      RECT -3.995 1.97 -3.77 2.348 ;
      RECT -3.995 1.97 -3.76 2.338 ;
      RECT -3.995 1.97 -3.755 2.333 ;
      RECT -3.995 1.975 -3.75 2.328 ;
      RECT -3.995 2.007 -3.735 2.318 ;
      RECT -3.995 2.077 -3.71 2.301 ;
      RECT -4.015 2.077 -3.71 2.293 ;
      RECT -4.015 2.137 -3.7 2.27 ;
      RECT -4.015 2.177 -3.69 2.215 ;
      RECT -4.03 1.97 -3.755 2.195 ;
      RECT -4.04 1.985 -3.75 2.093 ;
      RECT -4.45 3.375 -4.28 3.9 ;
      RECT -4.455 3.375 -4.28 3.893 ;
      RECT -4.465 3.375 -4.275 3.858 ;
      RECT -4.47 3.385 -4.275 3.83 ;
      RECT -4.475 3.405 -4.275 3.813 ;
      RECT -4.465 3.38 -4.27 3.803 ;
      RECT -4.48 3.425 -4.27 3.795 ;
      RECT -4.485 3.445 -4.27 3.78 ;
      RECT -4.49 3.475 -4.27 3.77 ;
      RECT -4.5 3.52 -4.27 3.745 ;
      RECT -4.47 3.39 -4.265 3.728 ;
      RECT -4.505 3.572 -4.265 3.723 ;
      RECT -4.47 3.4 -4.26 3.693 ;
      RECT -4.51 3.605 -4.26 3.69 ;
      RECT -4.515 3.63 -4.26 3.67 ;
      RECT -4.475 3.417 -4.25 3.61 ;
      RECT -4.48 3.439 -4.24 3.503 ;
      RECT -4.53 2.686 -4.515 2.955 ;
      RECT -4.575 2.67 -4.53 3 ;
      RECT -4.58 2.658 -4.575 3.05 ;
      RECT -4.59 2.654 -4.58 3.083 ;
      RECT -4.595 2.651 -4.59 3.111 ;
      RECT -4.61 2.653 -4.595 3.153 ;
      RECT -4.615 2.657 -4.61 3.193 ;
      RECT -4.635 2.662 -4.615 3.245 ;
      RECT -4.639 2.667 -4.635 3.302 ;
      RECT -4.725 2.686 -4.639 3.339 ;
      RECT -4.735 2.707 -4.725 3.375 ;
      RECT -4.74 2.715 -4.735 3.376 ;
      RECT -4.745 2.757 -4.74 3.377 ;
      RECT -4.76 2.845 -4.745 3.378 ;
      RECT -4.77 2.995 -4.76 3.38 ;
      RECT -4.775 3.04 -4.77 3.382 ;
      RECT -4.81 3.082 -4.775 3.385 ;
      RECT -4.815 3.1 -4.81 3.388 ;
      RECT -4.892 3.106 -4.815 3.394 ;
      RECT -4.978 3.12 -4.892 3.407 ;
      RECT -5.064 3.134 -4.978 3.421 ;
      RECT -5.15 3.148 -5.064 3.434 ;
      RECT -5.21 3.16 -5.15 3.446 ;
      RECT -5.235 3.167 -5.21 3.453 ;
      RECT -5.249 3.17 -5.235 3.458 ;
      RECT -5.335 3.178 -5.249 3.474 ;
      RECT -5.34 3.185 -5.335 3.489 ;
      RECT -5.364 3.185 -5.34 3.496 ;
      RECT -5.45 3.188 -5.364 3.524 ;
      RECT -5.535 3.192 -5.45 3.568 ;
      RECT -5.6 3.196 -5.535 3.605 ;
      RECT -5.625 3.199 -5.6 3.621 ;
      RECT -5.7 3.212 -5.625 3.625 ;
      RECT -5.725 3.23 -5.7 3.629 ;
      RECT -5.735 3.237 -5.725 3.631 ;
      RECT -5.75 3.24 -5.735 3.632 ;
      RECT -5.81 3.252 -5.75 3.636 ;
      RECT -5.82 3.266 -5.81 3.64 ;
      RECT -5.875 3.276 -5.82 3.628 ;
      RECT -5.9 3.297 -5.875 3.611 ;
      RECT -5.92 3.317 -5.9 3.602 ;
      RECT -5.925 3.33 -5.92 3.597 ;
      RECT -5.94 3.342 -5.925 3.593 ;
      RECT -4.705 1.997 -4.7 2.02 ;
      RECT -4.71 1.988 -4.705 2.06 ;
      RECT -4.715 1.986 -4.71 2.103 ;
      RECT -4.72 1.977 -4.715 2.138 ;
      RECT -4.725 1.967 -4.72 2.21 ;
      RECT -4.73 1.957 -4.725 2.275 ;
      RECT -4.735 1.954 -4.73 2.315 ;
      RECT -4.76 1.948 -4.735 2.405 ;
      RECT -4.795 1.936 -4.76 2.43 ;
      RECT -4.805 1.927 -4.795 2.43 ;
      RECT -4.94 1.925 -4.93 2.413 ;
      RECT -4.95 1.925 -4.94 2.38 ;
      RECT -4.955 1.925 -4.95 2.355 ;
      RECT -4.96 1.925 -4.955 2.343 ;
      RECT -4.965 1.925 -4.96 2.325 ;
      RECT -4.975 1.925 -4.965 2.29 ;
      RECT -4.98 1.927 -4.975 2.268 ;
      RECT -4.985 1.933 -4.98 2.253 ;
      RECT -4.99 1.939 -4.985 2.238 ;
      RECT -5.005 1.951 -4.99 2.211 ;
      RECT -5.01 1.962 -5.005 2.179 ;
      RECT -5.015 1.972 -5.01 2.163 ;
      RECT -5.025 1.98 -5.015 2.132 ;
      RECT -5.03 1.99 -5.025 2.106 ;
      RECT -5.035 2.047 -5.03 2.089 ;
      RECT -4.93 1.925 -4.805 2.43 ;
      RECT -5.215 2.612 -4.955 2.91 ;
      RECT -5.22 2.619 -4.955 2.908 ;
      RECT -5.215 2.614 -4.94 2.903 ;
      RECT -5.225 2.627 -4.94 2.9 ;
      RECT -5.225 2.632 -4.935 2.893 ;
      RECT -5.23 2.64 -4.935 2.89 ;
      RECT -5.23 2.657 -4.93 2.688 ;
      RECT -5.215 2.609 -4.984 2.91 ;
      RECT -5.16 2.608 -4.984 2.91 ;
      RECT -5.16 2.605 -5.07 2.91 ;
      RECT -5.16 2.602 -5.074 2.91 ;
      RECT -5.47 2.875 -5.465 2.888 ;
      RECT -5.475 2.842 -5.47 2.893 ;
      RECT -5.48 2.797 -5.475 2.9 ;
      RECT -5.485 2.752 -5.48 2.908 ;
      RECT -5.49 2.72 -5.485 2.916 ;
      RECT -5.495 2.68 -5.49 2.917 ;
      RECT -5.51 2.66 -5.495 2.919 ;
      RECT -5.585 2.642 -5.51 2.931 ;
      RECT -5.595 2.635 -5.585 2.942 ;
      RECT -5.6 2.635 -5.595 2.944 ;
      RECT -5.63 2.641 -5.6 2.948 ;
      RECT -5.67 2.654 -5.63 2.948 ;
      RECT -5.695 2.665 -5.67 2.934 ;
      RECT -5.71 2.671 -5.695 2.917 ;
      RECT -5.72 2.673 -5.71 2.908 ;
      RECT -5.725 2.674 -5.72 2.903 ;
      RECT -5.73 2.675 -5.725 2.898 ;
      RECT -5.735 2.676 -5.73 2.895 ;
      RECT -5.76 2.681 -5.735 2.885 ;
      RECT -5.77 2.697 -5.76 2.872 ;
      RECT -5.775 2.717 -5.77 2.867 ;
      RECT -5.765 2.11 -5.76 2.306 ;
      RECT -5.78 2.074 -5.765 2.308 ;
      RECT -5.79 2.056 -5.78 2.313 ;
      RECT -5.8 2.042 -5.79 2.317 ;
      RECT -5.845 2.026 -5.8 2.327 ;
      RECT -5.85 2.016 -5.845 2.336 ;
      RECT -5.895 2.005 -5.85 2.342 ;
      RECT -5.9 1.993 -5.895 2.349 ;
      RECT -5.915 1.988 -5.9 2.353 ;
      RECT -5.93 1.98 -5.915 2.358 ;
      RECT -5.94 1.973 -5.93 2.363 ;
      RECT -5.95 1.97 -5.94 2.368 ;
      RECT -5.96 1.97 -5.95 2.369 ;
      RECT -5.965 1.967 -5.96 2.368 ;
      RECT -6 1.962 -5.975 2.367 ;
      RECT -6.024 1.958 -6 2.366 ;
      RECT -6.11 1.949 -6.024 2.363 ;
      RECT -6.125 1.941 -6.11 2.36 ;
      RECT -6.147 1.94 -6.125 2.359 ;
      RECT -6.233 1.94 -6.147 2.357 ;
      RECT -6.319 1.94 -6.233 2.355 ;
      RECT -6.405 1.94 -6.319 2.352 ;
      RECT -6.415 1.94 -6.405 2.343 ;
      RECT -6.445 1.94 -6.415 2.303 ;
      RECT -6.455 1.95 -6.445 2.258 ;
      RECT -6.46 1.99 -6.455 2.243 ;
      RECT -6.465 2.005 -6.46 2.23 ;
      RECT -6.495 2.085 -6.465 2.192 ;
      RECT -5.975 1.965 -5.965 2.368 ;
      RECT -6.15 2.73 -6.135 3.335 ;
      RECT -6.145 2.725 -6.135 3.335 ;
      RECT -5.98 2.725 -5.975 2.908 ;
      RECT -5.99 2.725 -5.98 2.938 ;
      RECT -6.005 2.725 -5.99 2.998 ;
      RECT -6.01 2.725 -6.005 3.043 ;
      RECT -6.015 2.725 -6.01 3.073 ;
      RECT -6.02 2.725 -6.015 3.093 ;
      RECT -6.03 2.725 -6.02 3.128 ;
      RECT -6.045 2.725 -6.03 3.16 ;
      RECT -6.09 2.725 -6.045 3.188 ;
      RECT -6.095 2.725 -6.09 3.218 ;
      RECT -6.1 2.725 -6.095 3.23 ;
      RECT -6.105 2.725 -6.1 3.238 ;
      RECT -6.115 2.725 -6.105 3.253 ;
      RECT -6.12 2.725 -6.115 3.275 ;
      RECT -6.13 2.725 -6.12 3.298 ;
      RECT -6.135 2.725 -6.13 3.318 ;
      RECT -6.17 2.74 -6.15 3.335 ;
      RECT -6.195 2.757 -6.17 3.335 ;
      RECT -6.2 2.767 -6.195 3.335 ;
      RECT -6.23 2.782 -6.2 3.335 ;
      RECT -6.305 2.824 -6.23 3.335 ;
      RECT -6.31 2.855 -6.305 3.318 ;
      RECT -6.315 2.859 -6.31 3.3 ;
      RECT -6.32 2.863 -6.315 3.263 ;
      RECT -6.325 3.047 -6.32 3.23 ;
      RECT -6.84 3.236 -6.754 3.801 ;
      RECT -6.885 3.238 -6.72 3.795 ;
      RECT -6.754 3.235 -6.72 3.795 ;
      RECT -6.84 3.237 -6.635 3.789 ;
      RECT -6.885 3.247 -6.625 3.785 ;
      RECT -6.91 3.239 -6.635 3.781 ;
      RECT -6.915 3.242 -6.635 3.776 ;
      RECT -6.94 3.257 -6.625 3.77 ;
      RECT -6.94 3.282 -6.585 3.765 ;
      RECT -6.98 3.29 -6.585 3.74 ;
      RECT -6.98 3.317 -6.57 3.738 ;
      RECT -6.98 3.347 -6.56 3.725 ;
      RECT -6.985 3.492 -6.56 3.713 ;
      RECT -6.98 3.421 -6.54 3.71 ;
      RECT -6.98 3.478 -6.535 3.518 ;
      RECT -6.79 2.757 -6.62 2.935 ;
      RECT -6.84 2.696 -6.79 2.92 ;
      RECT -7.105 2.676 -6.84 2.905 ;
      RECT -7.145 2.74 -6.67 2.905 ;
      RECT -7.145 2.73 -6.715 2.905 ;
      RECT -7.145 2.727 -6.725 2.905 ;
      RECT -7.145 2.715 -6.735 2.905 ;
      RECT -7.145 2.7 -6.79 2.905 ;
      RECT -7.105 2.672 -6.904 2.905 ;
      RECT -7.095 2.65 -6.904 2.905 ;
      RECT -7.07 2.635 -6.99 2.905 ;
      RECT -7.315 3.165 -7.195 3.61 ;
      RECT -7.33 3.165 -7.195 3.609 ;
      RECT -7.375 3.187 -7.195 3.604 ;
      RECT -7.415 3.236 -7.195 3.598 ;
      RECT -7.415 3.236 -7.19 3.573 ;
      RECT -7.415 3.236 -7.17 3.463 ;
      RECT -7.42 3.266 -7.17 3.46 ;
      RECT -7.33 3.165 -7.16 3.355 ;
      RECT -7.67 1.95 -7.665 2.395 ;
      RECT -7.86 1.95 -7.84 2.36 ;
      RECT -7.89 1.95 -7.885 2.335 ;
      RECT -7.21 2.257 -7.195 2.445 ;
      RECT -7.215 2.242 -7.21 2.451 ;
      RECT -7.235 2.215 -7.215 2.454 ;
      RECT -7.285 2.182 -7.235 2.463 ;
      RECT -7.315 2.162 -7.285 2.467 ;
      RECT -7.334 2.15 -7.315 2.463 ;
      RECT -7.42 2.122 -7.334 2.453 ;
      RECT -7.43 2.097 -7.42 2.443 ;
      RECT -7.5 2.065 -7.43 2.435 ;
      RECT -7.525 2.025 -7.5 2.427 ;
      RECT -7.545 2.007 -7.525 2.421 ;
      RECT -7.555 1.997 -7.545 2.418 ;
      RECT -7.565 1.99 -7.555 2.416 ;
      RECT -7.585 1.977 -7.565 2.413 ;
      RECT -7.595 1.967 -7.585 2.41 ;
      RECT -7.605 1.96 -7.595 2.408 ;
      RECT -7.655 1.952 -7.605 2.402 ;
      RECT -7.665 1.95 -7.655 2.396 ;
      RECT -7.695 1.95 -7.67 2.393 ;
      RECT -7.724 1.95 -7.695 2.388 ;
      RECT -7.81 1.95 -7.724 2.378 ;
      RECT -7.84 1.95 -7.81 2.365 ;
      RECT -7.885 1.95 -7.86 2.348 ;
      RECT -7.9 1.95 -7.89 2.33 ;
      RECT -7.92 1.957 -7.9 2.315 ;
      RECT -7.925 1.972 -7.92 2.303 ;
      RECT -7.93 1.977 -7.925 2.243 ;
      RECT -7.935 1.982 -7.93 2.085 ;
      RECT -7.94 1.985 -7.935 2.003 ;
      RECT -7.675 2.67 -7.589 2.991 ;
      RECT -7.675 2.67 -7.555 2.984 ;
      RECT -7.725 2.67 -7.555 2.98 ;
      RECT -7.725 2.672 -7.469 2.978 ;
      RECT -7.725 2.674 -7.445 2.972 ;
      RECT -7.725 2.681 -7.435 2.971 ;
      RECT -7.725 2.69 -7.43 2.968 ;
      RECT -7.725 2.696 -7.425 2.963 ;
      RECT -7.725 2.74 -7.42 2.96 ;
      RECT -7.725 2.832 -7.415 2.957 ;
      RECT -8.2 3.275 -8.165 3.595 ;
      RECT -7.615 3.46 -7.61 3.642 ;
      RECT -7.66 3.342 -7.615 3.661 ;
      RECT -7.675 3.319 -7.66 3.684 ;
      RECT -7.685 3.309 -7.675 3.694 ;
      RECT -7.705 3.304 -7.685 3.707 ;
      RECT -7.73 3.302 -7.705 3.728 ;
      RECT -7.749 3.301 -7.73 3.74 ;
      RECT -7.835 3.298 -7.749 3.74 ;
      RECT -7.905 3.293 -7.835 3.728 ;
      RECT -7.98 3.289 -7.905 3.703 ;
      RECT -8.045 3.285 -7.98 3.67 ;
      RECT -8.115 3.282 -8.045 3.63 ;
      RECT -8.145 3.278 -8.115 3.605 ;
      RECT -8.165 3.276 -8.145 3.598 ;
      RECT -8.249 3.274 -8.2 3.596 ;
      RECT -8.335 3.271 -8.249 3.597 ;
      RECT -8.41 3.27 -8.335 3.599 ;
      RECT -8.495 3.27 -8.41 3.625 ;
      RECT -8.572 3.271 -8.495 3.65 ;
      RECT -8.658 3.272 -8.572 3.65 ;
      RECT -8.744 3.272 -8.658 3.65 ;
      RECT -8.83 3.273 -8.744 3.65 ;
      RECT -8.85 3.274 -8.83 3.642 ;
      RECT -8.865 3.28 -8.85 3.627 ;
      RECT -8.9 3.3 -8.865 3.607 ;
      RECT -8.91 3.32 -8.9 3.589 ;
      RECT -7.94 2.625 -7.935 2.895 ;
      RECT -7.945 2.616 -7.94 2.9 ;
      RECT -7.955 2.606 -7.945 2.912 ;
      RECT -7.96 2.595 -7.955 2.923 ;
      RECT -7.98 2.589 -7.96 2.941 ;
      RECT -8.025 2.586 -7.98 2.99 ;
      RECT -8.04 2.585 -8.025 3.035 ;
      RECT -8.045 2.585 -8.04 3.048 ;
      RECT -8.055 2.585 -8.045 3.06 ;
      RECT -8.06 2.586 -8.055 3.075 ;
      RECT -8.08 2.594 -8.06 3.08 ;
      RECT -8.11 2.61 -8.08 3.08 ;
      RECT -8.12 2.622 -8.115 3.08 ;
      RECT -8.155 2.637 -8.12 3.08 ;
      RECT -8.185 2.657 -8.155 3.08 ;
      RECT -8.195 2.682 -8.185 3.08 ;
      RECT -8.2 2.71 -8.195 3.08 ;
      RECT -8.205 2.74 -8.2 3.08 ;
      RECT -8.21 2.757 -8.205 3.08 ;
      RECT -8.22 2.785 -8.21 3.08 ;
      RECT -8.23 2.82 -8.22 3.08 ;
      RECT -8.235 2.855 -8.23 3.08 ;
      RECT -8.115 2.62 -8.11 3.08 ;
      RECT -8.6 2.722 -8.415 2.895 ;
      RECT -8.64 2.64 -8.455 2.893 ;
      RECT -8.679 2.645 -8.455 2.889 ;
      RECT -8.765 2.654 -8.455 2.884 ;
      RECT -8.849 2.67 -8.45 2.879 ;
      RECT -8.935 2.69 -8.425 2.873 ;
      RECT -8.935 2.71 -8.42 2.873 ;
      RECT -8.849 2.68 -8.425 2.879 ;
      RECT -8.765 2.655 -8.45 2.884 ;
      RECT -8.6 2.637 -8.455 2.895 ;
      RECT -8.6 2.632 -8.5 2.895 ;
      RECT -8.514 2.626 -8.5 2.895 ;
      RECT -9.125 1.95 -9.12 2.349 ;
      RECT -9.38 1.95 -9.345 2.347 ;
      RECT -9.785 1.985 -9.78 2.341 ;
      RECT -9.04 1.988 -9.035 2.243 ;
      RECT -9.045 1.986 -9.04 2.249 ;
      RECT -9.05 1.985 -9.045 2.256 ;
      RECT -9.075 1.978 -9.05 2.28 ;
      RECT -9.08 1.971 -9.075 2.304 ;
      RECT -9.085 1.967 -9.08 2.313 ;
      RECT -9.095 1.962 -9.085 2.326 ;
      RECT -9.1 1.959 -9.095 2.335 ;
      RECT -9.105 1.957 -9.1 2.34 ;
      RECT -9.12 1.953 -9.105 2.35 ;
      RECT -9.135 1.947 -9.125 2.349 ;
      RECT -9.173 1.945 -9.135 2.349 ;
      RECT -9.259 1.947 -9.173 2.349 ;
      RECT -9.345 1.949 -9.259 2.348 ;
      RECT -9.416 1.95 -9.38 2.347 ;
      RECT -9.502 1.952 -9.416 2.347 ;
      RECT -9.588 1.954 -9.502 2.346 ;
      RECT -9.674 1.956 -9.588 2.346 ;
      RECT -9.76 1.959 -9.674 2.345 ;
      RECT -9.77 1.965 -9.76 2.344 ;
      RECT -9.78 1.977 -9.77 2.342 ;
      RECT -9.84 2.012 -9.785 2.338 ;
      RECT -9.845 2.042 -9.84 2.1 ;
      RECT -9.1 3.122 -9.085 3.315 ;
      RECT -9.105 3.09 -9.1 3.315 ;
      RECT -9.115 3.065 -9.105 3.315 ;
      RECT -9.12 3.037 -9.115 3.315 ;
      RECT -9.15 2.96 -9.12 3.315 ;
      RECT -9.175 2.842 -9.15 3.315 ;
      RECT -9.18 2.78 -9.175 3.315 ;
      RECT -9.19 2.767 -9.18 3.315 ;
      RECT -9.21 2.757 -9.19 3.315 ;
      RECT -9.225 2.74 -9.21 3.315 ;
      RECT -9.255 2.728 -9.225 3.315 ;
      RECT -9.26 2.727 -9.255 3.26 ;
      RECT -9.265 2.727 -9.26 3.218 ;
      RECT -9.28 2.726 -9.265 3.17 ;
      RECT -9.295 2.726 -9.28 3.108 ;
      RECT -9.315 2.726 -9.295 3.068 ;
      RECT -9.32 2.726 -9.315 3.053 ;
      RECT -9.345 2.725 -9.32 3.048 ;
      RECT -9.415 2.724 -9.345 3.035 ;
      RECT -9.43 2.723 -9.415 3.02 ;
      RECT -9.46 2.722 -9.43 3.003 ;
      RECT -9.465 2.722 -9.46 2.988 ;
      RECT -9.515 2.721 -9.465 2.968 ;
      RECT -9.58 2.72 -9.515 2.923 ;
      RECT -9.585 2.72 -9.58 2.895 ;
      RECT -9.5 3.257 -9.495 3.514 ;
      RECT -9.52 3.176 -9.5 3.531 ;
      RECT -9.54 3.17 -9.52 3.56 ;
      RECT -9.6 3.157 -9.54 3.58 ;
      RECT -9.645 3.141 -9.6 3.581 ;
      RECT -9.729 3.129 -9.645 3.569 ;
      RECT -9.815 3.116 -9.729 3.553 ;
      RECT -9.825 3.109 -9.815 3.545 ;
      RECT -9.87 3.106 -9.825 3.485 ;
      RECT -9.89 3.102 -9.87 3.4 ;
      RECT -9.905 3.1 -9.89 3.353 ;
      RECT -9.935 3.097 -9.905 3.323 ;
      RECT -9.97 3.093 -9.935 3.3 ;
      RECT -10.013 3.088 -9.97 3.288 ;
      RECT -10.099 3.079 -10.013 3.297 ;
      RECT -10.185 3.068 -10.099 3.309 ;
      RECT -10.25 3.059 -10.185 3.318 ;
      RECT -10.27 3.05 -10.25 3.323 ;
      RECT -10.275 3.043 -10.27 3.325 ;
      RECT -10.315 3.028 -10.275 3.322 ;
      RECT -10.335 3.007 -10.315 3.317 ;
      RECT -10.35 2.995 -10.335 3.31 ;
      RECT -10.355 2.987 -10.35 3.303 ;
      RECT -10.37 2.967 -10.355 3.296 ;
      RECT -10.375 2.83 -10.37 3.29 ;
      RECT -10.455 2.719 -10.375 3.262 ;
      RECT -10.464 2.712 -10.455 3.228 ;
      RECT -10.55 2.706 -10.464 3.153 ;
      RECT -10.575 2.697 -10.55 3.065 ;
      RECT -10.605 2.692 -10.575 3.04 ;
      RECT -10.67 2.701 -10.605 3.025 ;
      RECT -10.69 2.717 -10.67 3 ;
      RECT -10.7 2.723 -10.69 2.948 ;
      RECT -10.72 2.745 -10.7 2.83 ;
      RECT -10.065 2.71 -9.895 2.895 ;
      RECT -10.065 2.71 -9.86 2.893 ;
      RECT -10.015 2.62 -9.845 2.884 ;
      RECT -10.065 2.777 -9.84 2.877 ;
      RECT -10.05 2.655 -9.845 2.884 ;
      RECT -10.85 3.388 -10.785 3.831 ;
      RECT -10.91 3.413 -10.785 3.829 ;
      RECT -10.91 3.413 -10.73 3.823 ;
      RECT -10.925 3.438 -10.73 3.822 ;
      RECT -10.785 3.375 -10.71 3.819 ;
      RECT -10.85 3.4 -10.63 3.813 ;
      RECT -10.925 3.439 -10.585 3.807 ;
      RECT -10.94 3.466 -10.585 3.798 ;
      RECT -10.925 3.459 -10.565 3.79 ;
      RECT -10.94 3.468 -10.56 3.773 ;
      RECT -10.945 3.485 -10.56 3.6 ;
      RECT -10.94 2.207 -10.905 2.445 ;
      RECT -10.94 2.207 -10.875 2.444 ;
      RECT -10.94 2.207 -10.76 2.44 ;
      RECT -10.94 2.207 -10.705 2.418 ;
      RECT -10.93 2.15 -10.65 2.318 ;
      RECT -10.825 1.99 -10.795 2.441 ;
      RECT -10.795 1.985 -10.615 2.198 ;
      RECT -10.925 2.126 -10.615 2.198 ;
      RECT -10.875 2.022 -10.825 2.442 ;
      RECT -10.905 2.078 -10.615 2.198 ;
      RECT 5.895 0.575 6.065 1.085 ;
      RECT 5.895 2.395 6.065 3.865 ;
      RECT 5.895 5.015 6.065 6.485 ;
      RECT 5.895 7.795 6.065 8.305 ;
      RECT 4.905 0.575 5.075 1.085 ;
      RECT 4.905 2.395 5.075 3.865 ;
      RECT 4.905 5.015 5.075 6.485 ;
      RECT 4.905 7.795 5.075 8.305 ;
      RECT 3.54 0.575 3.71 3.865 ;
      RECT 3.54 5.015 3.71 8.305 ;
      RECT 3.11 0.575 3.28 1.085 ;
      RECT 3.11 1.655 3.28 3.865 ;
      RECT 3.11 5.015 3.28 7.225 ;
      RECT 3.11 7.795 3.28 8.305 ;
      RECT 1.74 1.66 1.91 2.935 ;
      RECT 1.74 5.945 1.91 7.22 ;
  END
END sky130_osu_single_mpr2at_8

MACRO sky130_osu_single_mpr2ca_8
  CLASS CORE ;
  ORIGIN 8.04 0 ;
  FOREIGN sky130_osu_single_mpr2ca_8 -8.04 0 ;
  SIZE 14.475 BY 8.88 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT -1.66 2.735 -1.33 3.065 ;
      RECT -1.66 2.75 -0.86 3.05 ;
      RECT -1.66 3.755 -1.33 4.085 ;
      RECT -1.66 3.77 -0.86 4.07 ;
      RECT -1.655 3.705 -1.355 4.085 ;
      RECT -2.34 5.795 -2.01 6.125 ;
      RECT -2.34 5.81 -1.54 6.11 ;
      RECT -2.335 5.79 -2.035 6.125 ;
      RECT -2.36 3.075 -2.03 3.405 ;
      RECT -2.83 3.09 -2.03 3.39 ;
      RECT -2.335 3.06 -2.035 3.405 ;
      RECT -3.02 4.775 -2.69 5.105 ;
      RECT -3.02 4.79 -2.22 5.09 ;
      RECT -3.385 5.795 -3.055 6.125 ;
      RECT -3.855 5.81 -3.055 6.11 ;
      RECT -3.7 2.39 -3.37 2.72 ;
      RECT -4.17 2.41 -3.81 2.71 ;
      RECT -3.81 2.405 -3.37 2.705 ;
      RECT -4.09 6.49 -3.79 6.905 ;
      RECT -4.06 6.475 -3.73 6.805 ;
      RECT -4.53 6.49 -3.73 6.79 ;
    LAYER via2 ;
      RECT -1.595 2.8 -1.395 3 ;
      RECT -1.595 3.82 -1.395 4.02 ;
      RECT -2.275 5.86 -2.075 6.06 ;
      RECT -2.295 3.14 -2.095 3.34 ;
      RECT -2.955 4.84 -2.755 5.04 ;
      RECT -3.32 5.86 -3.12 6.06 ;
      RECT -3.635 2.455 -3.435 2.655 ;
      RECT -3.995 6.54 -3.795 6.74 ;
    LAYER met2 ;
      RECT 2.705 6.28 3.025 6.605 ;
      RECT 2.735 5.695 2.905 6.605 ;
      RECT 2.735 5.695 2.91 6.045 ;
      RECT 2.735 5.695 3.71 5.87 ;
      RECT 3.535 1.965 3.71 5.87 ;
      RECT 1.035 1.995 1.36 2.32 ;
      RECT 3.48 1.965 3.83 2.315 ;
      RECT 1.035 2.025 3.83 2.195 ;
      RECT 3.505 6.655 3.83 6.98 ;
      RECT 2.39 6.745 3.83 6.915 ;
      RECT 2.39 2.395 2.55 6.915 ;
      RECT 0.45 3.185 0.775 3.51 ;
      RECT 0.45 3.225 2.55 3.4 ;
      RECT 0.495 1.605 0.695 3.51 ;
      RECT -3.675 2.37 -3.395 2.74 ;
      RECT 2.705 2.365 3.025 2.685 ;
      RECT 2.39 2.395 3.025 2.565 ;
      RECT -3.655 1.605 -3.455 2.74 ;
      RECT -3.655 1.605 0.695 1.805 ;
      RECT 1.665 5.865 1.99 6.19 ;
      RECT 1.73 3.635 1.905 6.19 ;
      RECT 1.66 3.635 1.985 3.96 ;
      RECT -4.035 6.455 -3.755 6.825 ;
      RECT -4.035 6.625 1.24 6.79 ;
      RECT 1.075 3.655 1.24 6.79 ;
      RECT 0.95 3.655 1.275 3.98 ;
      RECT 0.065 4.78 0.325 5.1 ;
      RECT 0.125 2.74 0.265 5.1 ;
      RECT 0.065 2.74 0.325 3.06 ;
      RECT -0.955 5.8 -0.695 6.12 ;
      RECT -1.575 5.89 -0.695 6.03 ;
      RECT -1.575 3.735 -1.435 6.03 ;
      RECT -1.635 3.735 -1.355 4.105 ;
      RECT -2.315 5.775 -2.035 6.145 ;
      RECT -2.255 3.85 -2.115 6.145 ;
      RECT -2.255 3.85 -1.775 3.99 ;
      RECT -1.915 2.06 -1.775 3.99 ;
      RECT -1.975 2.06 -1.715 2.38 ;
      RECT -2.995 4.755 -2.715 5.125 ;
      RECT -2.935 2.4 -2.795 5.125 ;
      RECT -2.995 2.4 -2.735 2.72 ;
      RECT -3.36 5.775 -3.08 6.145 ;
      RECT -3.36 5.8 -3.075 6.12 ;
      RECT -1.635 2.715 -1.355 3.085 ;
      RECT -2.335 3.055 -2.055 3.425 ;
    LAYER via1 ;
      RECT 3.595 6.74 3.745 6.89 ;
      RECT 3.58 2.065 3.73 2.215 ;
      RECT 2.79 2.45 2.94 2.6 ;
      RECT 2.79 6.37 2.94 6.52 ;
      RECT 1.755 5.95 1.905 6.1 ;
      RECT 1.75 3.72 1.9 3.87 ;
      RECT 1.125 2.08 1.275 2.23 ;
      RECT 1.04 3.74 1.19 3.89 ;
      RECT 0.54 3.27 0.69 3.42 ;
      RECT 0.12 2.825 0.27 2.975 ;
      RECT 0.12 4.865 0.27 5.015 ;
      RECT -0.9 5.885 -0.75 6.035 ;
      RECT -1.58 2.825 -1.43 2.975 ;
      RECT -1.58 3.845 -1.43 3.995 ;
      RECT -1.92 2.145 -1.77 2.295 ;
      RECT -2.26 3.165 -2.11 3.315 ;
      RECT -2.26 5.885 -2.11 6.035 ;
      RECT -2.94 2.485 -2.79 2.635 ;
      RECT -2.94 4.865 -2.79 5.015 ;
      RECT -3.28 5.885 -3.13 6.035 ;
      RECT -3.62 2.48 -3.47 2.63 ;
      RECT -3.96 6.565 -3.81 6.715 ;
    LAYER met1 ;
      RECT -6.435 0 0.465 1.95 ;
      RECT -6.435 0 0.655 1.795 ;
      RECT -6.69 0 0.655 1.655 ;
      RECT -8.035 0 6.435 0.305 ;
      RECT 0.495 4.15 6.435 4.745 ;
      RECT 0.955 4.135 6.435 4.745 ;
      RECT -8.035 4.13 -6.575 4.74 ;
      RECT -8.035 4.19 6.435 4.67 ;
      RECT 0.365 4.15 6.435 4.67 ;
      RECT -8.035 8.575 6.435 8.88 ;
      RECT -6.73 7.18 0.47 8.88 ;
      RECT -6.435 6.91 0.465 8.88 ;
      RECT 5.835 2.365 6.125 2.595 ;
      RECT 5.895 0.885 6.065 2.595 ;
      RECT 5.835 0.885 6.125 1.115 ;
      RECT 5.835 7.765 6.125 7.995 ;
      RECT 5.895 6.285 6.065 7.995 ;
      RECT 5.835 6.285 6.125 6.515 ;
      RECT 5.425 2.735 5.755 2.965 ;
      RECT 5.425 2.765 5.925 2.935 ;
      RECT 5.425 2.395 5.615 2.965 ;
      RECT 4.845 2.365 5.135 2.595 ;
      RECT 4.845 2.395 5.615 2.565 ;
      RECT 4.905 0.885 5.075 2.595 ;
      RECT 4.845 0.885 5.135 1.115 ;
      RECT 4.845 7.765 5.135 7.995 ;
      RECT 4.905 6.285 5.075 7.995 ;
      RECT 4.845 6.285 5.135 6.515 ;
      RECT 4.845 6.325 5.695 6.485 ;
      RECT 5.525 5.915 5.695 6.485 ;
      RECT 4.845 6.32 5.235 6.485 ;
      RECT 5.465 5.915 5.755 6.145 ;
      RECT 5.465 5.945 5.925 6.115 ;
      RECT 4.475 2.735 4.765 2.965 ;
      RECT 4.475 2.765 4.935 2.935 ;
      RECT 4.535 1.655 4.7 2.965 ;
      RECT 3.05 1.625 3.34 1.855 ;
      RECT 3.05 1.655 4.7 1.825 ;
      RECT 3.11 0.885 3.28 1.855 ;
      RECT 3.05 0.885 3.34 1.115 ;
      RECT 3.05 7.765 3.34 7.995 ;
      RECT 3.11 7.025 3.28 7.995 ;
      RECT 3.11 7.12 4.7 7.29 ;
      RECT 4.53 5.915 4.7 7.29 ;
      RECT 3.05 7.025 3.34 7.255 ;
      RECT 4.475 5.915 4.765 6.145 ;
      RECT 4.475 5.945 4.935 6.115 ;
      RECT 3.48 1.965 3.83 2.315 ;
      RECT 3.31 2.025 3.83 2.195 ;
      RECT 3.505 6.655 3.83 6.98 ;
      RECT 3.48 6.655 3.83 6.885 ;
      RECT 3.31 6.685 3.83 6.855 ;
      RECT 2.705 2.365 3.025 2.685 ;
      RECT 2.675 2.365 3.025 2.595 ;
      RECT 2.39 2.395 3.025 2.565 ;
      RECT 2.705 6.28 3.025 6.605 ;
      RECT 2.675 6.285 3.025 6.515 ;
      RECT 2.505 6.315 3.025 6.485 ;
      RECT 1.66 3.635 1.985 3.96 ;
      RECT 1.735 2.735 1.915 3.96 ;
      RECT 1.68 2.735 1.97 2.965 ;
      RECT 1.68 2.765 2.14 2.935 ;
      RECT 1.665 5.865 1.99 6.19 ;
      RECT 1.665 5.945 2.14 6.115 ;
      RECT 0.955 3.655 1.275 3.995 ;
      RECT 0.95 3.655 1.275 3.67 ;
      RECT 1.075 1.995 1.24 3.995 ;
      RECT 1.035 1.995 1.36 2.32 ;
      RECT 0.035 2.77 0.355 3.03 ;
      RECT -0.24 2.83 0.355 2.97 ;
      RECT -2.345 3.11 -2.025 3.37 ;
      RECT -0.37 3.125 -0.08 3.355 ;
      RECT -2.345 3.17 -0.08 3.31 ;
      RECT -0.985 5.83 -0.665 6.09 ;
      RECT -0.985 5.89 -0.39 6.03 ;
      RECT -1.665 2.77 -1.345 3.03 ;
      RECT -6.405 2.785 -6.115 3.015 ;
      RECT -6.405 2.83 -1.345 2.97 ;
      RECT -1.575 2.49 -1.435 3.03 ;
      RECT -1.575 2.49 -1.095 2.63 ;
      RECT -1.235 2.105 -1.095 2.63 ;
      RECT -1.31 2.105 -1.02 2.335 ;
      RECT -1.665 3.79 -1.345 4.05 ;
      RECT -2.33 3.805 -2.04 4.035 ;
      RECT -4.54 3.805 -4.25 4.035 ;
      RECT -4.54 3.85 -1.345 3.99 ;
      RECT -3.365 5.83 -3.045 6.09 ;
      RECT -1.65 5.845 -1.36 6.075 ;
      RECT -4.03 5.845 -3.74 6.075 ;
      RECT -4.03 5.89 -3.045 6.03 ;
      RECT -1.575 5.55 -1.435 6.075 ;
      RECT -3.275 5.55 -3.135 6.09 ;
      RECT -3.275 5.55 -1.435 5.69 ;
      RECT -4.37 2.445 -4.08 2.675 ;
      RECT -4.295 2.15 -4.155 2.675 ;
      RECT -2.005 2.09 -1.685 2.35 ;
      RECT -2.105 2.105 -1.685 2.335 ;
      RECT -4.295 2.15 -1.685 2.29 ;
      RECT -3.025 2.43 -2.705 2.69 ;
      RECT -3.025 2.49 -2.43 2.63 ;
      RECT -4.045 6.51 -3.725 6.77 ;
      RECT -4.975 6.57 -2.625 6.71 ;
      RECT -2.765 5.845 -2.625 6.71 ;
      RECT -4.975 5.845 -4.835 6.71 ;
      RECT -2.84 5.845 -2.55 6.075 ;
      RECT -5.05 5.845 -4.76 6.075 ;
      RECT -3.025 4.81 -2.705 5.07 ;
      RECT -5.73 4.825 -5.44 5.055 ;
      RECT -5.73 4.87 -2.705 5.01 ;
      RECT -3.7 2.39 -3.37 2.72 ;
      RECT -3.705 2.425 -3.37 2.685 ;
      RECT -3.355 2.445 -3.24 2.675 ;
      RECT -3.705 2.44 -3.355 2.67 ;
      RECT -3.705 2.49 -3.225 2.63 ;
      RECT -3.82 2.49 -3.81 2.63 ;
      RECT -3.81 2.485 -3.24 2.625 ;
      RECT 0.45 3.185 0.775 3.51 ;
      RECT -0.29 4.81 0.355 5.07 ;
      RECT -2.345 5.83 -2.025 6.09 ;
    LAYER mcon ;
      RECT 5.895 0.915 6.065 1.085 ;
      RECT 5.895 2.395 6.065 2.565 ;
      RECT 5.895 6.315 6.065 6.485 ;
      RECT 5.895 7.795 6.065 7.965 ;
      RECT 5.545 0.105 5.715 0.275 ;
      RECT 5.545 4.165 5.715 4.335 ;
      RECT 5.545 4.545 5.715 4.715 ;
      RECT 5.545 8.605 5.715 8.775 ;
      RECT 5.525 2.765 5.695 2.935 ;
      RECT 5.525 5.945 5.695 6.115 ;
      RECT 4.905 0.915 5.075 1.085 ;
      RECT 4.905 2.395 5.075 2.565 ;
      RECT 4.905 6.315 5.075 6.485 ;
      RECT 4.905 7.795 5.075 7.965 ;
      RECT 4.555 0.105 4.725 0.275 ;
      RECT 4.555 4.165 4.725 4.335 ;
      RECT 4.555 4.545 4.725 4.715 ;
      RECT 4.555 8.605 4.725 8.775 ;
      RECT 4.535 2.765 4.705 2.935 ;
      RECT 4.535 5.945 4.705 6.115 ;
      RECT 3.85 0.105 4.02 0.275 ;
      RECT 3.85 4.165 4.02 4.335 ;
      RECT 3.85 4.545 4.02 4.715 ;
      RECT 3.85 8.605 4.02 8.775 ;
      RECT 3.54 2.025 3.71 2.195 ;
      RECT 3.54 6.685 3.71 6.855 ;
      RECT 3.17 0.105 3.34 0.275 ;
      RECT 3.17 8.605 3.34 8.775 ;
      RECT 3.11 0.915 3.28 1.085 ;
      RECT 3.11 1.655 3.28 1.825 ;
      RECT 3.11 7.055 3.28 7.225 ;
      RECT 3.11 7.795 3.28 7.965 ;
      RECT 2.735 2.395 2.905 2.565 ;
      RECT 2.735 6.315 2.905 6.485 ;
      RECT 2.49 0.105 2.66 0.275 ;
      RECT 2.49 8.605 2.66 8.775 ;
      RECT 1.81 0.105 1.98 0.275 ;
      RECT 1.81 8.605 1.98 8.775 ;
      RECT 1.74 2.765 1.91 2.935 ;
      RECT 1.74 5.945 1.91 6.115 ;
      RECT 0.15 1.625 0.32 1.795 ;
      RECT 0.15 4.345 0.32 4.515 ;
      RECT 0.15 7.065 0.32 7.235 ;
      RECT 0.11 2.815 0.28 2.985 ;
      RECT -0.23 4.855 -0.06 5.025 ;
      RECT -0.31 1.625 -0.14 1.795 ;
      RECT -0.31 3.155 -0.14 3.325 ;
      RECT -0.31 4.345 -0.14 4.515 ;
      RECT -0.31 7.065 -0.14 7.235 ;
      RECT -0.77 1.625 -0.6 1.795 ;
      RECT -0.77 4.345 -0.6 4.515 ;
      RECT -0.77 7.065 -0.6 7.235 ;
      RECT -0.91 5.875 -0.74 6.045 ;
      RECT -1.23 1.625 -1.06 1.795 ;
      RECT -1.23 4.345 -1.06 4.515 ;
      RECT -1.23 7.065 -1.06 7.235 ;
      RECT -1.25 2.135 -1.08 2.305 ;
      RECT -1.59 5.875 -1.42 6.045 ;
      RECT -1.69 1.625 -1.52 1.795 ;
      RECT -1.69 4.345 -1.52 4.515 ;
      RECT -1.69 7.065 -1.52 7.235 ;
      RECT -2.045 2.135 -1.875 2.305 ;
      RECT -2.15 1.625 -1.98 1.795 ;
      RECT -2.15 4.345 -1.98 4.515 ;
      RECT -2.15 7.065 -1.98 7.235 ;
      RECT -2.27 3.835 -2.1 4.005 ;
      RECT -2.27 5.875 -2.1 6.045 ;
      RECT -2.61 1.625 -2.44 1.795 ;
      RECT -2.61 4.345 -2.44 4.515 ;
      RECT -2.61 7.065 -2.44 7.235 ;
      RECT -2.78 5.875 -2.61 6.045 ;
      RECT -2.95 2.475 -2.78 2.645 ;
      RECT -3.07 1.625 -2.9 1.795 ;
      RECT -3.07 4.345 -2.9 4.515 ;
      RECT -3.07 7.065 -2.9 7.235 ;
      RECT -3.53 1.625 -3.36 1.795 ;
      RECT -3.53 4.345 -3.36 4.515 ;
      RECT -3.53 7.065 -3.36 7.235 ;
      RECT -3.97 5.875 -3.8 6.045 ;
      RECT -3.99 1.625 -3.82 1.795 ;
      RECT -3.99 4.345 -3.82 4.515 ;
      RECT -3.99 7.065 -3.82 7.235 ;
      RECT -4.31 2.475 -4.14 2.645 ;
      RECT -4.45 1.625 -4.28 1.795 ;
      RECT -4.45 4.345 -4.28 4.515 ;
      RECT -4.45 7.065 -4.28 7.235 ;
      RECT -4.48 3.835 -4.31 4.005 ;
      RECT -4.91 1.625 -4.74 1.795 ;
      RECT -4.91 4.345 -4.74 4.515 ;
      RECT -4.91 7.065 -4.74 7.235 ;
      RECT -4.99 5.875 -4.82 6.045 ;
      RECT -5.37 1.625 -5.2 1.795 ;
      RECT -5.37 4.345 -5.2 4.515 ;
      RECT -5.37 7.065 -5.2 7.235 ;
      RECT -5.67 4.855 -5.5 5.025 ;
      RECT -5.83 1.625 -5.66 1.795 ;
      RECT -5.83 4.345 -5.66 4.515 ;
      RECT -5.83 7.065 -5.66 7.235 ;
      RECT -6.29 1.625 -6.12 1.795 ;
      RECT -6.29 4.345 -6.12 4.515 ;
      RECT -6.29 7.065 -6.12 7.235 ;
      RECT -6.345 2.815 -6.175 2.985 ;
    LAYER li ;
      RECT -6.35 0 -6.09 2.615 ;
      RECT 0.1 0 0.37 2.605 ;
      RECT -0.81 0 -0.57 2.605 ;
      RECT -1.68 0 -1.43 2.335 ;
      RECT -4.06 0 -3.73 2.255 ;
      RECT -6.435 0 0.655 1.795 ;
      RECT -6.69 0 0.655 1.655 ;
      RECT 5.465 0 5.635 0.935 ;
      RECT 4.475 0 4.645 0.935 ;
      RECT 1.73 0 1.9 0.935 ;
      RECT -8.035 0 6.435 0.305 ;
      RECT 5.465 3.405 5.635 5.475 ;
      RECT 4.475 3.405 4.645 5.475 ;
      RECT 1.73 3.405 1.9 5.475 ;
      RECT -3.08 3.69 -2.815 5.295 ;
      RECT -5.24 3.84 -4.91 5.235 ;
      RECT -4.24 4.345 -3.96 5.185 ;
      RECT -2.265 4.345 -1.89 4.895 ;
      RECT 0.495 4.135 6.435 4.745 ;
      RECT -8.035 4.13 -6.575 4.74 ;
      RECT 0.365 4.135 6.435 4.67 ;
      RECT -8.035 4.345 6.435 4.515 ;
      RECT 0.04 3.205 0.37 4.515 ;
      RECT -1.7 3.8 -1.445 4.515 ;
      RECT -3.13 3.69 -2.525 4.515 ;
      RECT -4 3.8 -3.785 4.515 ;
      RECT -5.43 3.84 -4.815 4.515 ;
      RECT -5.01 3.475 -4.815 4.515 ;
      RECT -6.35 3.835 -6.09 4.515 ;
      RECT -2.7 3.42 -2.515 3.79 ;
      RECT -2.7 3.42 -2.37 3.665 ;
      RECT -5.01 3.475 -4.68 3.665 ;
      RECT -8.035 8.575 6.435 8.88 ;
      RECT 5.465 7.945 5.635 8.88 ;
      RECT 4.475 7.945 4.645 8.88 ;
      RECT 1.73 7.945 1.9 8.88 ;
      RECT -6.73 7.18 0.47 8.88 ;
      RECT -6.435 7.065 0.465 8.88 ;
      RECT -1 6.555 -0.55 8.88 ;
      RECT -3.09 6.665 -2.76 8.88 ;
      RECT -5.16 6.605 -4.91 8.88 ;
      RECT 5.525 1.74 5.695 2.935 ;
      RECT 5.525 1.74 5.99 1.91 ;
      RECT 5.525 6.97 5.99 7.14 ;
      RECT 5.525 5.945 5.695 7.14 ;
      RECT 4.535 1.74 4.705 2.935 ;
      RECT 4.535 1.74 5 1.91 ;
      RECT 4.535 6.97 5 7.14 ;
      RECT 4.535 5.945 4.705 7.14 ;
      RECT 2.68 2.635 2.85 3.865 ;
      RECT 2.735 0.855 2.905 2.805 ;
      RECT 2.68 0.575 2.85 1.025 ;
      RECT 2.68 7.855 2.85 8.305 ;
      RECT 2.735 6.075 2.905 8.025 ;
      RECT 2.68 5.015 2.85 6.245 ;
      RECT 2.16 0.575 2.33 3.865 ;
      RECT 2.16 2.075 2.565 2.405 ;
      RECT 2.16 1.235 2.565 1.565 ;
      RECT 2.16 5.015 2.33 8.305 ;
      RECT 2.16 7.315 2.565 7.645 ;
      RECT 2.16 6.475 2.565 6.805 ;
      RECT -2.58 6.645 -1.275 6.895 ;
      RECT -2.58 6.325 -2.4 6.895 ;
      RECT -3.13 6.325 -2.4 6.495 ;
      RECT -3.13 5.485 -2.96 6.495 ;
      RECT -2.295 5.525 -0.55 5.705 ;
      RECT -0.88 4.685 -0.55 5.705 ;
      RECT -3.13 5.485 -2.07 5.655 ;
      RECT -0.88 4.855 -0.06 5.025 ;
      RECT -1.72 4.685 -1.39 4.895 ;
      RECT -1.72 4.685 -0.55 4.855 ;
      RECT -0.82 3.205 -0.49 4.16 ;
      RECT -0.82 3.205 -0.14 3.375 ;
      RECT -0.31 1.965 -0.14 3.375 ;
      RECT -0.4 1.965 -0.07 2.605 ;
      RECT -1.275 3.475 -1 4.175 ;
      RECT -1.17 1.965 -1 4.175 ;
      RECT -0.83 2.785 -0.48 3.035 ;
      RECT -1.17 2.815 -0.48 2.985 ;
      RECT -1.26 1.965 -1 2.445 ;
      RECT -1.93 5.115 -1.05 5.355 ;
      RECT -1.28 5.025 -1.05 5.355 ;
      RECT -2.58 5.115 -1.05 5.315 ;
      RECT -1.665 5.065 -1.05 5.355 ;
      RECT -2.58 4.985 -2.41 5.315 ;
      RECT -1.695 5.875 -1.445 6.475 ;
      RECT -1.695 5.875 -1.22 6.075 ;
      RECT -2.2 3.095 -1.445 3.595 ;
      RECT -3.13 2.9 -2.87 3.52 ;
      RECT -2.215 3.04 -2.2 3.345 ;
      RECT -2.23 3.025 -2.21 3.31 ;
      RECT -1.57 2.7 -1.34 3.3 ;
      RECT -2.255 2.97 -2.235 3.285 ;
      RECT -2.275 3.095 -1.34 3.27 ;
      RECT -2.3 3.095 -1.34 3.26 ;
      RECT -2.37 3.095 -1.34 3.25 ;
      RECT -2.39 3.095 -1.34 3.22 ;
      RECT -2.41 2.005 -2.24 3.19 ;
      RECT -2.44 3.095 -1.34 3.16 ;
      RECT -2.475 3.095 -1.34 3.135 ;
      RECT -2.505 3.09 -2.115 3.1 ;
      RECT -2.505 3.08 -2.14 3.1 ;
      RECT -2.505 3.075 -2.155 3.1 ;
      RECT -2.505 3.065 -2.17 3.1 ;
      RECT -3.13 2.9 -2.24 3.07 ;
      RECT -3.13 3.055 -2.18 3.07 ;
      RECT -3.13 3.05 -2.19 3.07 ;
      RECT -2.235 2.995 -2.225 3.3 ;
      RECT -3.13 3.03 -2.205 3.07 ;
      RECT -3.13 3.01 -2.22 3.07 ;
      RECT -3.13 2.005 -2.24 2.175 ;
      RECT -2.07 2.5 -1.74 2.925 ;
      RECT -2.07 2.015 -1.85 2.925 ;
      RECT -2.155 5.875 -1.945 6.475 ;
      RECT -2.295 5.875 -1.945 6.075 ;
      RECT -3.575 3.475 -3.3 4.175 ;
      RECT -3.355 1.965 -3.3 4.175 ;
      RECT -3.47 2.77 -3.3 4.175 ;
      RECT -3.47 1.965 -3.3 2.765 ;
      RECT -3.56 1.965 -3.3 2.44 ;
      RECT -5.43 3.135 -5.18 3.67 ;
      RECT -4.46 3.135 -3.745 3.6 ;
      RECT -5.43 3.135 -3.64 3.305 ;
      RECT -3.87 2.77 -3.64 3.305 ;
      RECT -4.875 2.015 -4.62 3.305 ;
      RECT -3.87 2.705 -3.81 3.6 ;
      RECT -3.81 2.7 -3.64 2.765 ;
      RECT -5.41 2.015 -4.62 2.28 ;
      RECT -4.45 5.825 -3.775 6.075 ;
      RECT -4.04 5.465 -3.775 6.075 ;
      RECT -4.29 6.245 -3.96 6.795 ;
      RECT -5.35 6.245 -3.96 6.435 ;
      RECT -5.35 5.405 -5.18 6.435 ;
      RECT -5.47 5.825 -5.18 6.155 ;
      RECT -5.35 5.405 -4.41 5.575 ;
      RECT -4.71 4.855 -4.41 5.575 ;
      RECT -4.45 2.435 -4.04 2.955 ;
      RECT -4.45 2.015 -4.25 2.955 ;
      RECT -5.84 2.195 -5.67 4.175 ;
      RECT -5.84 2.705 -5.045 2.955 ;
      RECT -5.84 2.195 -5.59 2.955 ;
      RECT -5.92 2.195 -5.59 2.615 ;
      RECT -5.89 6.605 -5.33 6.895 ;
      RECT -5.89 4.685 -5.64 6.895 ;
      RECT -5.89 4.685 -5.43 5.235 ;
      RECT 5.895 0.575 6.065 1.085 ;
      RECT 5.895 2.395 6.065 3.865 ;
      RECT 5.895 5.015 6.065 6.485 ;
      RECT 5.895 7.795 6.065 8.305 ;
      RECT 4.905 0.575 5.075 1.085 ;
      RECT 4.905 2.395 5.075 3.865 ;
      RECT 4.905 5.015 5.075 6.485 ;
      RECT 4.905 7.795 5.075 8.305 ;
      RECT 3.54 0.575 3.71 3.865 ;
      RECT 3.54 5.015 3.71 8.305 ;
      RECT 3.11 0.575 3.28 1.085 ;
      RECT 3.11 1.655 3.28 3.865 ;
      RECT 3.11 5.015 3.28 7.225 ;
      RECT 3.11 7.795 3.28 8.305 ;
      RECT 1.74 1.66 1.91 2.935 ;
      RECT 1.74 5.945 1.91 7.22 ;
      RECT 0.03 2.785 0.38 3.035 ;
      RECT -1.03 5.875 -0.58 6.385 ;
      RECT -2.35 3.835 -1.87 4.175 ;
      RECT -2.79 5.825 -2.465 6.155 ;
      RECT -3.13 2.345 -2.58 2.73 ;
      RECT -4.645 3.835 -4.17 4.175 ;
      RECT -5.01 5.825 -4.67 6.075 ;
      RECT -6.35 2.785 -6.01 3.665 ;
  END
END sky130_osu_single_mpr2ca_8

MACRO sky130_osu_single_mpr2ct_8
  CLASS CORE ;
  ORIGIN 8.04 0 ;
  FOREIGN sky130_osu_single_mpr2ct_8 -8.04 0 ;
  SIZE 14.475 BY 8.88 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT -1.885 5.79 -1.555 6.12 ;
      RECT -1.885 5.805 -1.085 6.105 ;
      RECT -1.83 5.765 -1.53 6.105 ;
      RECT -2.235 3.755 -1.905 4.085 ;
      RECT -2.235 3.77 -1.435 4.07 ;
      RECT -2.22 3.725 -1.92 4.085 ;
      RECT -2.575 3.075 -2.245 3.405 ;
      RECT -2.575 3.09 -1.775 3.39 ;
      RECT -2.49 3.065 -2.19 3.39 ;
      RECT -2.925 5.79 -2.595 6.12 ;
      RECT -3.395 5.805 -2.595 6.105 ;
      RECT -2.9 5.745 -2.6 6.12 ;
      RECT -3.255 4.155 -2.925 4.485 ;
      RECT -5.295 4.155 -4.965 4.485 ;
      RECT -5.295 4.17 -2.925 4.47 ;
      RECT -3.605 3.415 -3.275 3.745 ;
      RECT -4.065 3.43 -3.265 3.73 ;
      RECT -3.935 2.225 -3.605 2.555 ;
      RECT -4.405 2.24 -3.605 2.54 ;
      RECT -3.945 2.235 -3.605 2.54 ;
      RECT -3.935 6.48 -3.605 6.81 ;
      RECT -4.405 6.495 -3.605 6.795 ;
      RECT -4.025 6.455 -3.725 6.795 ;
      RECT -4.615 5.79 -4.285 6.12 ;
      RECT -5.085 5.805 -4.285 6.105 ;
    LAYER via2 ;
      RECT -1.82 5.855 -1.62 6.055 ;
      RECT -2.17 3.82 -1.97 4.02 ;
      RECT -2.51 3.14 -2.31 3.34 ;
      RECT -2.86 5.855 -2.66 6.055 ;
      RECT -3.19 4.22 -2.99 4.42 ;
      RECT -3.54 3.48 -3.34 3.68 ;
      RECT -3.87 2.29 -3.67 2.49 ;
      RECT -3.87 6.545 -3.67 6.745 ;
      RECT -4.55 5.855 -4.35 6.055 ;
      RECT -5.23 4.22 -5.03 4.42 ;
    LAYER met2 ;
      RECT 2.705 6.28 3.025 6.605 ;
      RECT 2.735 5.695 2.905 6.605 ;
      RECT 2.735 5.695 2.91 6.045 ;
      RECT 2.735 5.695 3.71 5.87 ;
      RECT 3.535 1.965 3.71 5.87 ;
      RECT 1.035 1.995 1.36 2.32 ;
      RECT 3.48 1.965 3.83 2.315 ;
      RECT 1.035 2.025 3.83 2.195 ;
      RECT 3.505 6.655 3.83 6.98 ;
      RECT 2.39 6.745 3.83 6.915 ;
      RECT 2.39 2.395 2.55 6.915 ;
      RECT 0.565 3.055 2.55 3.23 ;
      RECT 0.565 2.345 0.74 3.23 ;
      RECT 2.705 2.365 3.025 2.685 ;
      RECT -3.91 2.205 -3.63 2.575 ;
      RECT 2.39 2.395 3.025 2.565 ;
      RECT -3.91 2.345 0.74 2.52 ;
      RECT 1.66 5.855 1.985 6.18 ;
      RECT 1.73 3.495 1.9 6.18 ;
      RECT 1.66 3.495 1.985 3.82 ;
      RECT -4.57 7.295 0.95 7.46 ;
      RECT 0.785 3.815 0.95 7.46 ;
      RECT -4.57 5.77 -4.405 7.46 ;
      RECT -4.59 5.77 -4.31 6.14 ;
      RECT 0.95 3.655 1.275 3.98 ;
      RECT -0.84 6.48 -0.58 6.8 ;
      RECT -0.78 2.74 -0.64 6.8 ;
      RECT -0.84 2.74 -0.58 3.06 ;
      RECT -1.52 4.78 -1.26 5.1 ;
      RECT -1.46 3.76 -1.32 5.1 ;
      RECT -1.52 3.76 -1.26 4.08 ;
      RECT -2.54 6.48 -2.28 6.8 ;
      RECT -2.48 5.21 -2.34 6.8 ;
      RECT -3.16 5.21 -2.34 5.35 ;
      RECT -3.16 2.74 -3.02 5.35 ;
      RECT -3.23 4.135 -2.95 4.505 ;
      RECT -3.22 2.74 -2.96 3.06 ;
      RECT -5.27 4.135 -4.99 4.505 ;
      RECT -5.2 2.4 -5.06 4.505 ;
      RECT -5.26 2.4 -5 2.72 ;
      RECT -5.94 4.78 -5.68 5.1 ;
      RECT -5.88 2.74 -5.74 5.1 ;
      RECT -5.94 2.74 -5.68 3.06 ;
      RECT -1.86 5.77 -1.58 6.14 ;
      RECT -2.21 3.735 -1.93 4.105 ;
      RECT -2.55 3.055 -2.27 3.425 ;
      RECT -2.9 5.77 -2.62 6.14 ;
      RECT -3.58 3.395 -3.3 3.765 ;
      RECT -3.91 6.46 -3.63 6.83 ;
    LAYER via1 ;
      RECT 3.595 6.74 3.745 6.89 ;
      RECT 3.58 2.065 3.73 2.215 ;
      RECT 2.79 2.45 2.94 2.6 ;
      RECT 2.79 6.37 2.94 6.52 ;
      RECT 1.75 3.58 1.9 3.73 ;
      RECT 1.75 5.94 1.9 6.09 ;
      RECT 1.125 2.08 1.275 2.23 ;
      RECT 1.04 3.74 1.19 3.89 ;
      RECT -0.785 2.825 -0.635 2.975 ;
      RECT -0.785 6.565 -0.635 6.715 ;
      RECT -1.465 3.845 -1.315 3.995 ;
      RECT -1.465 4.865 -1.315 5.015 ;
      RECT -1.805 5.885 -1.655 6.035 ;
      RECT -2.145 3.845 -1.995 3.995 ;
      RECT -2.485 3.165 -2.335 3.315 ;
      RECT -2.485 6.565 -2.335 6.715 ;
      RECT -2.835 5.885 -2.685 6.035 ;
      RECT -3.165 2.825 -3.015 2.975 ;
      RECT -3.505 3.505 -3.355 3.655 ;
      RECT -3.845 2.315 -3.695 2.465 ;
      RECT -3.845 6.565 -3.695 6.715 ;
      RECT -4.525 5.885 -4.375 6.035 ;
      RECT -5.205 2.485 -5.055 2.635 ;
      RECT -5.885 2.825 -5.735 2.975 ;
      RECT -5.885 4.865 -5.735 5.015 ;
    LAYER met1 ;
      RECT -7 0 0.36 1.95 ;
      RECT -7 0 0.655 1.795 ;
      RECT -7.005 0 0.655 1.635 ;
      RECT -8.035 0 6.435 0.305 ;
      RECT 0.45 4.135 6.435 4.745 ;
      RECT -8.035 4.19 -6.625 4.74 ;
      RECT -8.035 4.19 6.435 4.67 ;
      RECT 0.445 4.135 6.435 4.67 ;
      RECT -8.035 4.13 -6.645 4.74 ;
      RECT -8.035 8.575 6.435 8.88 ;
      RECT -6.73 7.18 0.47 8.88 ;
      RECT -7 6.91 0.36 7.39 ;
      RECT 5.835 2.365 6.125 2.595 ;
      RECT 5.895 0.885 6.065 2.595 ;
      RECT 5.835 0.885 6.125 1.115 ;
      RECT 5.835 7.765 6.125 7.995 ;
      RECT 5.895 6.285 6.065 7.995 ;
      RECT 5.835 6.285 6.125 6.515 ;
      RECT 5.425 2.735 5.755 2.965 ;
      RECT 5.425 2.765 5.925 2.935 ;
      RECT 5.425 2.395 5.615 2.965 ;
      RECT 4.845 2.365 5.135 2.595 ;
      RECT 4.845 2.395 5.615 2.565 ;
      RECT 4.905 0.885 5.075 2.595 ;
      RECT 4.845 0.885 5.135 1.115 ;
      RECT 4.845 7.765 5.135 7.995 ;
      RECT 4.905 6.285 5.075 7.995 ;
      RECT 4.845 6.285 5.135 6.515 ;
      RECT 4.845 6.325 5.695 6.485 ;
      RECT 5.525 5.915 5.695 6.485 ;
      RECT 4.845 6.32 5.235 6.485 ;
      RECT 5.465 5.915 5.755 6.145 ;
      RECT 5.465 5.945 5.925 6.115 ;
      RECT 4.475 2.735 4.765 2.965 ;
      RECT 4.475 2.765 4.935 2.935 ;
      RECT 4.535 1.655 4.7 2.965 ;
      RECT 3.05 1.625 3.34 1.855 ;
      RECT 3.05 1.655 4.7 1.825 ;
      RECT 3.11 0.885 3.28 1.855 ;
      RECT 3.05 0.885 3.34 1.115 ;
      RECT 3.05 7.765 3.34 7.995 ;
      RECT 3.11 7.025 3.28 7.995 ;
      RECT 3.11 7.12 4.7 7.29 ;
      RECT 4.53 5.915 4.7 7.29 ;
      RECT 3.05 7.025 3.34 7.255 ;
      RECT 4.475 5.915 4.765 6.145 ;
      RECT 4.475 5.945 4.935 6.115 ;
      RECT 3.48 1.965 3.83 2.315 ;
      RECT 3.31 2.025 3.83 2.195 ;
      RECT 3.505 6.655 3.83 6.98 ;
      RECT 3.48 6.655 3.83 6.885 ;
      RECT 3.31 6.685 3.83 6.855 ;
      RECT 2.705 2.365 3.025 2.685 ;
      RECT 2.675 2.365 3.025 2.595 ;
      RECT 2.39 2.395 3.025 2.565 ;
      RECT 2.705 6.28 3.025 6.605 ;
      RECT 2.675 6.285 3.025 6.515 ;
      RECT 2.505 6.315 3.025 6.485 ;
      RECT 1.66 3.495 1.985 3.82 ;
      RECT 1.74 2.735 1.91 3.82 ;
      RECT 1.68 2.735 1.97 2.965 ;
      RECT 1.68 2.765 2.14 2.935 ;
      RECT 1.66 5.855 1.985 6.18 ;
      RECT 1.66 5.945 2.14 6.115 ;
      RECT 0.95 3.655 1.275 3.98 ;
      RECT 1.075 1.995 1.24 3.98 ;
      RECT 1.035 1.995 1.36 2.32 ;
      RECT -1.55 3.79 -1.23 4.05 ;
      RECT -0.515 3.805 -0.225 4.035 ;
      RECT -1.55 3.85 -0.225 3.99 ;
      RECT -1.89 5.83 -1.57 6.09 ;
      RECT -0.515 5.845 -0.225 6.075 ;
      RECT -0.44 5.55 -0.3 6.075 ;
      RECT -1.8 5.55 -1.66 6.09 ;
      RECT -1.8 5.55 -0.3 5.69 ;
      RECT -0.87 2.77 -0.55 3.03 ;
      RECT -1.145 2.83 -0.55 2.97 ;
      RECT -3.93 6.51 -3.61 6.77 ;
      RECT -4.935 6.525 -4.645 6.755 ;
      RECT -4.935 6.57 -3.02 6.71 ;
      RECT -3.16 6.23 -3.02 6.71 ;
      RECT -3.16 6.23 -1.15 6.37 ;
      RECT -1.29 5.845 -1.15 6.37 ;
      RECT -1.365 5.845 -1.075 6.075 ;
      RECT -1.55 4.81 -1.23 5.07 ;
      RECT -3.695 4.825 -3.405 5.055 ;
      RECT -3.695 4.87 -1.23 5.01 ;
      RECT -2.23 3.79 -1.91 4.05 ;
      RECT -4.595 3.805 -4.305 4.035 ;
      RECT -4.595 3.85 -1.91 3.99 ;
      RECT -2.57 6.51 -2.25 6.77 ;
      RECT -2.57 6.57 -1.975 6.71 ;
      RECT -2.57 3.11 -2.25 3.37 ;
      RECT -2.845 3.17 -2.25 3.31 ;
      RECT -3.25 2.77 -2.93 3.03 ;
      RECT -3.525 2.83 -2.93 2.97 ;
      RECT -3.59 3.45 -3.27 3.71 ;
      RECT -6.465 3.465 -6.175 3.695 ;
      RECT -6.465 3.51 -3.27 3.65 ;
      RECT -4.01 2.79 -3.87 3.65 ;
      RECT -4.085 2.79 -3.795 3.02 ;
      RECT -3.93 2.26 -3.61 2.52 ;
      RECT -3.93 2.275 -3.425 2.505 ;
      RECT -4.02 2.32 -3.425 2.46 ;
      RECT -4.61 5.83 -4.29 6.09 ;
      RECT -6.975 5.845 -6.685 6.075 ;
      RECT -6.975 5.89 -4.29 6.03 ;
      RECT -4.595 2.79 -4.305 3.02 ;
      RECT -5.2 2.835 -4.305 2.975 ;
      RECT -5.2 2.43 -5.06 2.975 ;
      RECT -5.29 2.43 -4.97 2.69 ;
      RECT -5.97 2.77 -5.65 3.03 ;
      RECT -6.245 2.83 -5.65 2.97 ;
      RECT -5.97 4.81 -5.65 5.07 ;
      RECT -6.245 4.87 -5.65 5.01 ;
      RECT -1.195 6.51 -0.55 6.77 ;
      RECT -3.245 5.83 -2.6 6.09 ;
    LAYER mcon ;
      RECT 5.895 0.915 6.065 1.085 ;
      RECT 5.895 2.395 6.065 2.565 ;
      RECT 5.895 6.315 6.065 6.485 ;
      RECT 5.895 7.795 6.065 7.965 ;
      RECT 5.545 0.105 5.715 0.275 ;
      RECT 5.545 4.165 5.715 4.335 ;
      RECT 5.545 4.545 5.715 4.715 ;
      RECT 5.545 8.605 5.715 8.775 ;
      RECT 5.525 2.765 5.695 2.935 ;
      RECT 5.525 5.945 5.695 6.115 ;
      RECT 4.905 0.915 5.075 1.085 ;
      RECT 4.905 2.395 5.075 2.565 ;
      RECT 4.905 6.315 5.075 6.485 ;
      RECT 4.905 7.795 5.075 7.965 ;
      RECT 4.555 0.105 4.725 0.275 ;
      RECT 4.555 4.165 4.725 4.335 ;
      RECT 4.555 4.545 4.725 4.715 ;
      RECT 4.555 8.605 4.725 8.775 ;
      RECT 4.535 2.765 4.705 2.935 ;
      RECT 4.535 5.945 4.705 6.115 ;
      RECT 3.85 0.105 4.02 0.275 ;
      RECT 3.85 4.165 4.02 4.335 ;
      RECT 3.85 4.545 4.02 4.715 ;
      RECT 3.85 8.605 4.02 8.775 ;
      RECT 3.54 2.025 3.71 2.195 ;
      RECT 3.54 6.685 3.71 6.855 ;
      RECT 3.17 0.105 3.34 0.275 ;
      RECT 3.17 8.605 3.34 8.775 ;
      RECT 3.11 0.915 3.28 1.085 ;
      RECT 3.11 1.655 3.28 1.825 ;
      RECT 3.11 7.055 3.28 7.225 ;
      RECT 3.11 7.795 3.28 7.965 ;
      RECT 2.735 2.395 2.905 2.565 ;
      RECT 2.735 6.315 2.905 6.485 ;
      RECT 2.49 0.105 2.66 0.275 ;
      RECT 2.49 8.605 2.66 8.775 ;
      RECT 1.81 0.105 1.98 0.275 ;
      RECT 1.81 8.605 1.98 8.775 ;
      RECT 1.74 2.765 1.91 2.935 ;
      RECT 1.74 5.945 1.91 6.115 ;
      RECT 0.045 1.625 0.215 1.795 ;
      RECT 0.045 4.345 0.215 4.515 ;
      RECT 0.045 7.065 0.215 7.235 ;
      RECT -0.415 1.625 -0.245 1.795 ;
      RECT -0.415 4.345 -0.245 4.515 ;
      RECT -0.415 7.065 -0.245 7.235 ;
      RECT -0.455 3.835 -0.285 4.005 ;
      RECT -0.455 5.875 -0.285 6.045 ;
      RECT -0.795 2.815 -0.625 2.985 ;
      RECT -0.875 1.625 -0.705 1.795 ;
      RECT -0.875 4.345 -0.705 4.515 ;
      RECT -0.875 7.065 -0.705 7.235 ;
      RECT -1.135 6.555 -0.965 6.725 ;
      RECT -1.305 5.875 -1.135 6.045 ;
      RECT -1.335 1.625 -1.165 1.795 ;
      RECT -1.335 4.345 -1.165 4.515 ;
      RECT -1.335 7.065 -1.165 7.235 ;
      RECT -1.795 1.625 -1.625 1.795 ;
      RECT -1.795 4.345 -1.625 4.515 ;
      RECT -1.795 7.065 -1.625 7.235 ;
      RECT -1.815 5.875 -1.645 6.045 ;
      RECT -2.255 1.625 -2.085 1.795 ;
      RECT -2.255 4.345 -2.085 4.515 ;
      RECT -2.255 7.065 -2.085 7.235 ;
      RECT -2.495 3.155 -2.325 3.325 ;
      RECT -2.495 6.555 -2.325 6.725 ;
      RECT -2.715 1.625 -2.545 1.795 ;
      RECT -2.715 4.345 -2.545 4.515 ;
      RECT -2.715 7.065 -2.545 7.235 ;
      RECT -3.175 1.625 -3.005 1.795 ;
      RECT -3.175 2.815 -3.005 2.985 ;
      RECT -3.175 4.345 -3.005 4.515 ;
      RECT -3.175 7.065 -3.005 7.235 ;
      RECT -3.185 5.875 -3.015 6.045 ;
      RECT -3.635 1.625 -3.465 1.795 ;
      RECT -3.635 4.345 -3.465 4.515 ;
      RECT -3.635 4.855 -3.465 5.025 ;
      RECT -3.635 7.065 -3.465 7.235 ;
      RECT -3.655 2.305 -3.485 2.475 ;
      RECT -4.025 2.82 -3.855 2.99 ;
      RECT -4.095 1.625 -3.925 1.795 ;
      RECT -4.095 4.345 -3.925 4.515 ;
      RECT -4.095 7.065 -3.925 7.235 ;
      RECT -4.535 2.82 -4.365 2.99 ;
      RECT -4.535 3.835 -4.365 4.005 ;
      RECT -4.535 5.875 -4.365 6.045 ;
      RECT -4.555 1.625 -4.385 1.795 ;
      RECT -4.555 4.345 -4.385 4.515 ;
      RECT -4.555 7.065 -4.385 7.235 ;
      RECT -4.875 6.555 -4.705 6.725 ;
      RECT -5.015 1.625 -4.845 1.795 ;
      RECT -5.015 4.345 -4.845 4.515 ;
      RECT -5.015 7.065 -4.845 7.235 ;
      RECT -5.475 1.625 -5.305 1.795 ;
      RECT -5.475 4.345 -5.305 4.515 ;
      RECT -5.475 7.065 -5.305 7.235 ;
      RECT -5.895 2.815 -5.725 2.985 ;
      RECT -5.895 4.855 -5.725 5.025 ;
      RECT -5.935 1.625 -5.765 1.795 ;
      RECT -5.935 4.345 -5.765 4.515 ;
      RECT -5.935 7.065 -5.765 7.235 ;
      RECT -6.395 1.625 -6.225 1.795 ;
      RECT -6.395 4.345 -6.225 4.515 ;
      RECT -6.395 7.065 -6.225 7.235 ;
      RECT -6.405 3.495 -6.235 3.665 ;
      RECT -6.855 1.625 -6.685 1.795 ;
      RECT -6.855 4.345 -6.685 4.515 ;
      RECT -6.855 7.065 -6.685 7.235 ;
      RECT -6.915 5.875 -6.745 6.045 ;
    LAYER li ;
      RECT -2.775 0 -2.485 2.63 ;
      RECT -5.975 0 -5.745 2.615 ;
      RECT -6.855 0 -6.645 2.615 ;
      RECT -3.225 0 -2.955 2.605 ;
      RECT -4.135 0 -3.895 2.605 ;
      RECT -4.585 0 -4.345 2.605 ;
      RECT -5.525 0 -5.255 2.605 ;
      RECT -0.105 0 0.225 2.185 ;
      RECT -0.945 0 -0.615 2.185 ;
      RECT -7 0 0.655 1.795 ;
      RECT -7.005 0 0.655 1.635 ;
      RECT 5.465 0 5.635 0.935 ;
      RECT 4.475 0 4.645 0.935 ;
      RECT 1.73 0 1.9 0.935 ;
      RECT -8.035 0 6.435 0.305 ;
      RECT -0.465 4.345 -0.185 5.655 ;
      RECT -1.395 4.345 -1.135 5.655 ;
      RECT -1.845 4.345 -1.565 5.655 ;
      RECT -2.775 4.345 -2.515 5.655 ;
      RECT -3.205 4.345 -2.945 5.655 ;
      RECT -4.155 4.345 -3.875 5.655 ;
      RECT -5.505 3.205 -5.245 5.655 ;
      RECT -6.455 4.345 -6.175 5.655 ;
      RECT 5.465 3.405 5.635 5.475 ;
      RECT 4.475 3.405 4.645 5.475 ;
      RECT 1.73 3.405 1.9 5.475 ;
      RECT 0.45 4.135 6.435 4.745 ;
      RECT -8.035 4.345 -6.625 4.74 ;
      RECT -8.035 4.345 6.435 4.515 ;
      RECT 0.445 4.135 6.435 4.515 ;
      RECT -0.865 3.495 -0.695 4.515 ;
      RECT -1.705 3.835 -1.535 4.515 ;
      RECT -3.285 3.205 -2.955 4.515 ;
      RECT -5.525 3.205 -5.195 4.515 ;
      RECT -5.975 3.205 -5.745 4.515 ;
      RECT -8.035 4.13 -6.645 4.74 ;
      RECT -6.855 3.205 -6.645 4.74 ;
      RECT -8.035 8.575 6.435 8.88 ;
      RECT 5.465 7.945 5.635 8.88 ;
      RECT 4.475 7.945 4.645 8.88 ;
      RECT 1.73 7.945 1.9 8.88 ;
      RECT -6.73 7.18 0.47 8.88 ;
      RECT -7 7.065 0.36 7.235 ;
      RECT -0.495 6.265 -0.185 8.88 ;
      RECT -1.875 6.265 -1.565 8.88 ;
      RECT -4.155 6.265 -3.845 8.88 ;
      RECT -6.455 6.265 -6.145 8.88 ;
      RECT 5.525 1.74 5.695 2.935 ;
      RECT 5.525 1.74 5.99 1.91 ;
      RECT 5.525 6.97 5.99 7.14 ;
      RECT 5.525 5.945 5.695 7.14 ;
      RECT 4.535 1.74 4.705 2.935 ;
      RECT 4.535 1.74 5 1.91 ;
      RECT 4.535 6.97 5 7.14 ;
      RECT 4.535 5.945 4.705 7.14 ;
      RECT 2.68 2.635 2.85 3.865 ;
      RECT 2.735 0.855 2.905 2.805 ;
      RECT 2.68 0.575 2.85 1.025 ;
      RECT 2.68 7.855 2.85 8.305 ;
      RECT 2.735 6.075 2.905 8.025 ;
      RECT 2.68 5.015 2.85 6.245 ;
      RECT 2.16 0.575 2.33 3.865 ;
      RECT 2.16 2.075 2.565 2.405 ;
      RECT 2.16 1.235 2.565 1.565 ;
      RECT 2.16 5.015 2.33 8.305 ;
      RECT 2.16 7.315 2.565 7.645 ;
      RECT 2.16 6.475 2.565 6.805 ;
      RECT -0.105 3.495 0.275 4.175 ;
      RECT 0.105 2.365 0.275 4.175 ;
      RECT -1.975 2.365 -1.745 3.035 ;
      RECT -1.975 2.365 0.275 2.535 ;
      RECT -0.445 2.045 -0.275 2.535 ;
      RECT -0.455 3.155 -0.285 4.005 ;
      RECT -1.37 3.155 -0.065 3.325 ;
      RECT -0.31 2.705 -0.065 3.325 ;
      RECT -1.37 2.785 -1.2 3.325 ;
      RECT -1.575 2.785 -1.2 2.955 ;
      RECT -1.395 6.265 -0.7 6.895 ;
      RECT -0.87 4.685 -0.7 6.895 ;
      RECT -0.965 4.685 -0.635 5.665 ;
      RECT -1.365 3.495 -1.035 4.175 ;
      RECT -2.275 3.495 -1.875 4.175 ;
      RECT -2.275 3.495 -1.035 3.665 ;
      RECT -2.775 3.075 -2.455 4.175 ;
      RECT -2.775 3.075 -2.325 3.325 ;
      RECT -2.775 3.075 -2.145 3.245 ;
      RECT -2.315 2.025 -2.145 3.245 ;
      RECT -2.315 2.025 -1.36 2.195 ;
      RECT -2.775 6.265 -2.08 6.895 ;
      RECT -2.25 4.685 -2.08 6.895 ;
      RECT -2.345 4.685 -2.015 5.665 ;
      RECT -2.755 5.825 -2.42 6.075 ;
      RECT -3.3 5.825 -2.965 6.075 ;
      RECT -3.3 5.875 -2.42 6.045 ;
      RECT -3.64 6.265 -2.945 6.895 ;
      RECT -3.64 4.685 -3.47 6.895 ;
      RECT -3.705 4.685 -3.375 5.665 ;
      RECT -4.145 3.205 -3.815 4.16 ;
      RECT -4.145 3.205 -3.465 3.375 ;
      RECT -3.635 1.965 -3.465 3.375 ;
      RECT -3.725 1.965 -3.395 2.605 ;
      RECT -4.145 5.825 -3.81 6.095 ;
      RECT -4.535 5.875 -3.81 6.045 ;
      RECT -4.665 3.205 -4.335 4.16 ;
      RECT -5.015 3.205 -4.335 3.375 ;
      RECT -5.015 1.965 -4.845 3.375 ;
      RECT -5.085 1.965 -4.755 2.605 ;
      RECT -4.875 5.875 -4.705 6.725 ;
      RECT -5.6 5.825 -5.265 6.075 ;
      RECT -5.6 5.875 -4.705 6.045 ;
      RECT -5.535 2.785 -5.185 3.035 ;
      RECT -6.055 2.785 -5.725 3.035 ;
      RECT -6.055 2.815 -5.185 2.985 ;
      RECT -5.94 6.265 -5.245 6.895 ;
      RECT -5.94 4.685 -5.77 6.895 ;
      RECT -6.005 4.685 -5.675 5.665 ;
      RECT -6.445 5.825 -6.11 6.095 ;
      RECT -6.915 5.875 -6.11 6.045 ;
      RECT -6.475 3.195 -6.145 4.175 ;
      RECT -6.475 1.965 -6.225 4.175 ;
      RECT -6.475 1.965 -6.145 2.595 ;
      RECT 5.895 0.575 6.065 1.085 ;
      RECT 5.895 2.395 6.065 3.865 ;
      RECT 5.895 5.015 6.065 6.485 ;
      RECT 5.895 7.795 6.065 8.305 ;
      RECT 4.905 0.575 5.075 1.085 ;
      RECT 4.905 2.395 5.075 3.865 ;
      RECT 4.905 5.015 5.075 6.485 ;
      RECT 4.905 7.795 5.075 8.305 ;
      RECT 3.54 0.575 3.71 3.865 ;
      RECT 3.54 5.015 3.71 8.305 ;
      RECT 3.11 0.575 3.28 1.085 ;
      RECT 3.11 1.655 3.28 3.865 ;
      RECT 3.11 5.015 3.28 7.225 ;
      RECT 3.11 7.795 3.28 8.305 ;
      RECT 1.74 1.66 1.91 2.935 ;
      RECT 1.74 5.945 1.91 7.22 ;
      RECT -0.53 5.825 -0.195 6.095 ;
      RECT -1.03 2.785 -0.48 2.985 ;
      RECT -1.375 5.825 -1.04 6.075 ;
      RECT -1.91 5.825 -1.575 6.095 ;
      RECT -3.295 2.785 -2.945 3.035 ;
      RECT -4.155 2.785 -3.805 3.035 ;
      RECT -4.675 2.785 -4.325 3.035 ;
  END
END sky130_osu_single_mpr2ct_8

MACRO sky130_osu_single_mpr2ea_8
  CLASS CORE ;
  ORIGIN 9.9 0 ;
  FOREIGN sky130_osu_single_mpr2ea_8 -9.9 0 ;
  SIZE 16.335 BY 8.88 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT -4.28 3.535 -3.95 3.865 ;
      RECT -5.485 3.55 -3.95 3.85 ;
      RECT -5.485 2.43 -5.185 3.85 ;
      RECT -5.74 2.415 -5.41 2.745 ;
      RECT -0.26 2.975 0.07 3.705 ;
      RECT -0.74 1.85 -0.41 2.58 ;
      RECT -2.34 2.575 -2.01 3.305 ;
      RECT -3.9 2.015 -3.57 2.745 ;
      RECT -4.78 2.015 -4.45 2.745 ;
      RECT -6.46 2.415 -6.13 3.145 ;
      RECT -7.46 1.855 -7.13 2.585 ;
      RECT -8.9 2.575 -8.57 3.305 ;
    LAYER via2 ;
      RECT -0.195 3.04 0.005 3.24 ;
      RECT -0.675 2.315 -0.475 2.515 ;
      RECT -2.275 3.04 -2.075 3.24 ;
      RECT -3.835 2.48 -3.635 2.68 ;
      RECT -4.215 3.6 -4.015 3.8 ;
      RECT -4.715 2.48 -4.515 2.68 ;
      RECT -5.675 2.48 -5.475 2.68 ;
      RECT -6.395 2.48 -6.195 2.68 ;
      RECT -7.395 1.92 -7.195 2.12 ;
      RECT -8.835 3.04 -8.635 3.24 ;
    LAYER met2 ;
      RECT 2.705 6.28 3.025 6.605 ;
      RECT 2.735 5.695 2.905 6.605 ;
      RECT 2.735 5.695 2.91 6.045 ;
      RECT 2.735 5.695 3.71 5.87 ;
      RECT 3.535 1.965 3.71 5.87 ;
      RECT -0.235 2.955 0.045 3.325 ;
      RECT -0.235 3.01 0.655 3.175 ;
      RECT 0.49 2.025 0.655 3.175 ;
      RECT -0.225 2.7 0.035 3.325 ;
      RECT 3.48 1.965 3.83 2.315 ;
      RECT 0.49 2.04 3.83 2.195 ;
      RECT 1.435 2.025 3.83 2.195 ;
      RECT 0.49 2.025 1.07 2.195 ;
      RECT 3.505 6.655 3.83 6.98 ;
      RECT 2.39 6.745 3.83 6.915 ;
      RECT 2.39 2.395 2.55 6.915 ;
      RECT 2.705 2.365 3.025 2.685 ;
      RECT 2.39 2.395 3.025 2.565 ;
      RECT 1.655 5.84 1.995 6.19 ;
      RECT 1.74 2.705 1.91 6.19 ;
      RECT 1.665 2.705 2.005 3.055 ;
      RECT -8.875 2.955 -8.595 3.325 ;
      RECT -8.865 1.29 -8.695 3.325 ;
      RECT 1.175 1.29 1.345 1.815 ;
      RECT 1.085 1.46 1.425 1.81 ;
      RECT -8.865 1.29 1.345 1.46 ;
      RECT -2.195 2.395 -1.915 2.765 ;
      RECT -3.265 2.42 -3.005 2.74 ;
      RECT -0.715 2.23 -0.435 2.6 ;
      RECT -0.105 2.14 0.155 2.46 ;
      RECT -3.205 1.58 -3.065 2.74 ;
      RECT -2.125 1.58 -1.985 2.765 ;
      RECT -1.005 2.23 0.155 2.37 ;
      RECT -1.005 1.58 -0.865 2.37 ;
      RECT -3.205 1.58 -0.865 1.72 ;
      RECT -3.175 3.72 -1 3.885 ;
      RECT -1.145 2.6 -1 3.885 ;
      RECT -4.255 3.515 -3.975 3.885 ;
      RECT -4.255 3.63 -3.035 3.77 ;
      RECT -1.425 2.6 -1 2.74 ;
      RECT -1.425 2.42 -1.165 2.74 ;
      RECT -8.085 4 -4.425 4.14 ;
      RECT -4.565 3.185 -4.425 4.14 ;
      RECT -8.085 3.07 -7.945 4.14 ;
      RECT -1.545 3.26 -1.285 3.58 ;
      RECT -4.565 3.185 -2.035 3.325 ;
      RECT -2.315 2.955 -2.035 3.325 ;
      RECT -8.085 3.07 -7.635 3.325 ;
      RECT -7.915 2.955 -7.635 3.325 ;
      RECT -1.545 3.07 -1.345 3.58 ;
      RECT -2.315 3.07 -1.345 3.21 ;
      RECT -1.745 1.86 -1.605 3.21 ;
      RECT -1.805 1.86 -1.545 2.18 ;
      RECT -7.905 2.42 -7.645 2.74 ;
      RECT -7.905 2.51 -6.865 2.65 ;
      RECT -7.005 1.72 -6.865 2.65 ;
      RECT -4.245 1.86 -3.985 2.18 ;
      RECT -7.005 1.72 -4.045 1.86 ;
      RECT -4.865 2.7 -4.605 3.02 ;
      RECT -4.865 2.7 -4.545 2.93 ;
      RECT -4.755 2.395 -4.475 2.765 ;
      RECT -5.165 3.26 -4.845 3.58 ;
      RECT -5.165 2.14 -5.025 3.58 ;
      RECT -5.225 2.14 -4.965 2.46 ;
      RECT -7.665 3.54 -7.405 3.86 ;
      RECT -7.665 3.63 -5.985 3.77 ;
      RECT -6.125 3.35 -5.985 3.77 ;
      RECT -6.125 3.35 -5.685 3.58 ;
      RECT -5.945 3.26 -5.685 3.58 ;
      RECT -6.625 2.42 -6.225 2.93 ;
      RECT -6.435 2.395 -6.155 2.765 ;
      RECT -6.685 2.42 -6.155 2.74 ;
      RECT -3.875 2.395 -3.595 2.765 ;
      RECT -5.715 2.395 -5.435 2.765 ;
      RECT -7.435 1.835 -7.155 2.205 ;
    LAYER via1 ;
      RECT 3.595 6.74 3.745 6.89 ;
      RECT 3.58 2.065 3.73 2.215 ;
      RECT 2.79 2.45 2.94 2.6 ;
      RECT 2.79 6.37 2.94 6.52 ;
      RECT 1.765 2.805 1.915 2.955 ;
      RECT 1.755 5.94 1.905 6.09 ;
      RECT 1.185 1.56 1.335 1.71 ;
      RECT -0.05 2.225 0.1 2.375 ;
      RECT -0.17 2.785 -0.02 2.935 ;
      RECT -1.37 2.505 -1.22 2.655 ;
      RECT -1.49 3.345 -1.34 3.495 ;
      RECT -1.75 1.945 -1.6 2.095 ;
      RECT -3.21 2.505 -3.06 2.655 ;
      RECT -3.81 2.505 -3.66 2.655 ;
      RECT -4.19 1.945 -4.04 2.095 ;
      RECT -4.81 2.785 -4.66 2.935 ;
      RECT -5.05 3.345 -4.9 3.495 ;
      RECT -5.17 2.225 -5.02 2.375 ;
      RECT -5.65 2.505 -5.5 2.655 ;
      RECT -5.89 3.345 -5.74 3.495 ;
      RECT -6.63 2.505 -6.48 2.655 ;
      RECT -7.37 1.945 -7.22 2.095 ;
      RECT -7.61 3.625 -7.46 3.775 ;
      RECT -7.85 2.505 -7.7 2.655 ;
      RECT -7.85 3.065 -7.7 3.215 ;
      RECT -8.81 3.065 -8.66 3.215 ;
    LAYER met1 ;
      RECT -9.15 0 0.51 1.74 ;
      RECT -9.15 0 0.665 1.585 ;
      RECT -9.895 0 6.435 0.305 ;
      RECT -9.895 4.135 6.435 4.745 ;
      RECT -9.15 3.98 0.51 4.745 ;
      RECT 5.835 2.365 6.125 2.595 ;
      RECT 5.895 0.885 6.065 2.595 ;
      RECT 5.835 0.885 6.125 1.115 ;
      RECT 5.835 7.765 6.125 7.995 ;
      RECT 5.895 6.285 6.065 7.995 ;
      RECT 5.835 6.285 6.125 6.515 ;
      RECT 5.425 2.735 5.755 2.965 ;
      RECT 5.425 2.765 5.925 2.935 ;
      RECT 5.425 2.395 5.615 2.965 ;
      RECT 4.845 2.365 5.135 2.595 ;
      RECT 4.845 2.395 5.615 2.565 ;
      RECT 4.905 0.885 5.075 2.595 ;
      RECT 4.845 0.885 5.135 1.115 ;
      RECT 4.845 7.765 5.135 7.995 ;
      RECT 4.905 6.285 5.075 7.995 ;
      RECT 4.845 6.285 5.135 6.515 ;
      RECT 4.845 6.325 5.695 6.485 ;
      RECT 5.525 5.915 5.695 6.485 ;
      RECT 4.845 6.32 5.235 6.485 ;
      RECT 5.465 5.915 5.755 6.145 ;
      RECT 5.465 5.945 5.925 6.115 ;
      RECT 4.475 2.735 4.765 2.965 ;
      RECT 4.475 2.765 4.935 2.935 ;
      RECT 4.535 1.655 4.7 2.965 ;
      RECT 3.05 1.625 3.34 1.855 ;
      RECT 3.05 1.655 4.7 1.825 ;
      RECT 3.11 0.885 3.28 1.855 ;
      RECT 3.05 0.885 3.34 1.115 ;
      RECT 3.05 7.765 3.34 7.995 ;
      RECT 3.11 7.025 3.28 7.995 ;
      RECT 3.11 7.12 4.7 7.29 ;
      RECT 4.53 5.915 4.7 7.29 ;
      RECT 3.05 7.025 3.34 7.255 ;
      RECT 4.475 5.915 4.765 6.145 ;
      RECT 4.475 5.945 4.935 6.115 ;
      RECT 3.48 1.965 3.83 2.315 ;
      RECT 3.31 2.025 3.83 2.195 ;
      RECT 3.505 6.655 3.83 6.98 ;
      RECT 3.48 6.655 3.83 6.885 ;
      RECT 3.31 6.685 3.83 6.855 ;
      RECT 2.705 2.365 3.025 2.685 ;
      RECT 2.675 2.365 3.025 2.595 ;
      RECT 1.175 2.395 3.025 2.565 ;
      RECT 1.175 1.46 1.345 2.565 ;
      RECT 1.085 1.46 1.425 1.81 ;
      RECT 2.705 6.28 3.025 6.605 ;
      RECT 2.675 6.285 3.025 6.515 ;
      RECT 2.505 6.315 3.025 6.485 ;
      RECT 1.665 2.705 2.005 3.055 ;
      RECT 1.665 2.765 2.14 2.935 ;
      RECT 1.655 5.84 1.995 6.19 ;
      RECT 1.655 5.945 2.14 6.115 ;
      RECT -0.84 2.465 -0.55 2.695 ;
      RECT -0.84 2.465 -0.385 2.65 ;
      RECT -0.525 2.37 0.095 2.51 ;
      RECT -0.135 2.17 0.185 2.43 ;
      RECT -1.745 2.93 -0.145 3.07 ;
      RECT -1.745 2.93 0.02 3.055 ;
      RECT -0.255 2.73 0.065 2.99 ;
      RECT -0.3 2.745 0.17 2.975 ;
      RECT -2.08 2.79 -1.605 2.975 ;
      RECT -2.08 2.745 -1.79 2.975 ;
      RECT -0.3 2.735 0.065 2.99 ;
      RECT -1.455 2.45 -1.135 2.71 ;
      RECT -1.455 2.45 -0.99 2.695 ;
      RECT -1.13 2.07 -0.99 2.695 ;
      RECT -1.13 2.07 -0.865 2.21 ;
      RECT -0.6 1.905 -0.31 2.135 ;
      RECT -1.005 1.95 -0.31 2.09 ;
      RECT -1.56 3.29 -1.27 3.815 ;
      RECT -1.575 3.29 -1.255 3.55 ;
      RECT -1.835 1.89 -1.515 2.15 ;
      RECT -1.835 1.905 -1.27 2.135 ;
      RECT -2.56 3.585 -2.27 3.815 ;
      RECT -2.365 2.23 -2.225 3.77 ;
      RECT -2.32 2.185 -2.03 2.415 ;
      RECT -2.725 2.23 -2.03 2.37 ;
      RECT -2.725 2.07 -2.585 2.37 ;
      RECT -4.185 2.07 -2.585 2.21 ;
      RECT -4.275 1.89 -3.955 2.15 ;
      RECT -4.275 1.905 -3.71 2.15 ;
      RECT -5.165 2.93 -2.585 3.07 ;
      RECT -2.8 2.745 -2.51 2.975 ;
      RECT -5.24 2.745 -4.575 2.975 ;
      RECT -4.895 2.73 -4.575 3.07 ;
      RECT -3.895 2.45 -3.575 2.71 ;
      RECT -3.895 2.465 -3.47 2.695 ;
      RECT -5.255 2.17 -4.935 2.43 ;
      RECT -4.76 2.185 -4.47 2.415 ;
      RECT -5.255 2.23 -4.47 2.37 ;
      RECT -5.135 3.29 -4.815 3.55 ;
      RECT -5.975 3.29 -5.655 3.55 ;
      RECT -5.135 3.305 -4.71 3.535 ;
      RECT -5.975 3.35 -4.71 3.49 ;
      RECT -6.44 3.025 -6.15 3.255 ;
      RECT -6.365 1.95 -6.225 3.255 ;
      RECT -6.715 2.45 -6.225 2.71 ;
      RECT -6.96 2.465 -6.225 2.695 ;
      RECT -5.96 1.905 -5.67 2.135 ;
      RECT -6.365 1.95 -5.67 2.09 ;
      RECT -7.2 3.305 -6.91 3.535 ;
      RECT -7.2 3.305 -6.745 3.49 ;
      RECT -6.885 2.93 -6.745 3.49 ;
      RECT -7.245 2.93 -6.745 3.07 ;
      RECT -7.245 1.95 -7.105 3.07 ;
      RECT -7.455 1.89 -7.135 2.15 ;
      RECT -7.695 3.57 -7.375 3.83 ;
      RECT -8.4 3.585 -8.11 3.815 ;
      RECT -8.4 3.63 -7.375 3.77 ;
      RECT -8.325 3.58 -8.065 3.77 ;
      RECT -7.935 2.45 -7.615 2.71 ;
      RECT -7.935 2.465 -7.39 2.695 ;
      RECT -7.935 3.01 -7.615 3.27 ;
      RECT -7.935 3.025 -7.39 3.255 ;
      RECT -8.895 3.01 -8.575 3.27 ;
      RECT -8.805 1.95 -8.665 3.27 ;
      RECT -8.4 1.905 -8.11 2.135 ;
      RECT -8.805 1.95 -8.11 2.09 ;
      RECT -9.89 8.575 6.435 8.88 ;
      RECT -3.295 2.45 -2.975 2.71 ;
      RECT -5.735 2.45 -5.415 2.71 ;
    LAYER mcon ;
      RECT 5.895 0.915 6.065 1.085 ;
      RECT 5.895 2.395 6.065 2.565 ;
      RECT 5.895 6.315 6.065 6.485 ;
      RECT 5.895 7.795 6.065 7.965 ;
      RECT 5.545 0.105 5.715 0.275 ;
      RECT 5.545 4.165 5.715 4.335 ;
      RECT 5.545 4.545 5.715 4.715 ;
      RECT 5.545 8.605 5.715 8.775 ;
      RECT 5.525 2.765 5.695 2.935 ;
      RECT 5.525 5.945 5.695 6.115 ;
      RECT 4.905 0.915 5.075 1.085 ;
      RECT 4.905 2.395 5.075 2.565 ;
      RECT 4.905 6.315 5.075 6.485 ;
      RECT 4.905 7.795 5.075 7.965 ;
      RECT 4.555 0.105 4.725 0.275 ;
      RECT 4.555 4.165 4.725 4.335 ;
      RECT 4.555 4.545 4.725 4.715 ;
      RECT 4.555 8.605 4.725 8.775 ;
      RECT 4.535 2.765 4.705 2.935 ;
      RECT 4.535 5.945 4.705 6.115 ;
      RECT 3.85 0.105 4.02 0.275 ;
      RECT 3.85 4.165 4.02 4.335 ;
      RECT 3.85 4.545 4.02 4.715 ;
      RECT 3.85 8.605 4.02 8.775 ;
      RECT 3.54 2.025 3.71 2.195 ;
      RECT 3.54 6.685 3.71 6.855 ;
      RECT 3.17 0.105 3.34 0.275 ;
      RECT 3.17 8.605 3.34 8.775 ;
      RECT 3.11 0.915 3.28 1.085 ;
      RECT 3.11 1.655 3.28 1.825 ;
      RECT 3.11 7.055 3.28 7.225 ;
      RECT 3.11 7.795 3.28 7.965 ;
      RECT 2.735 2.395 2.905 2.565 ;
      RECT 2.735 6.315 2.905 6.485 ;
      RECT 2.49 0.105 2.66 0.275 ;
      RECT 2.49 8.605 2.66 8.775 ;
      RECT 1.81 0.105 1.98 0.275 ;
      RECT 1.81 8.605 1.98 8.775 ;
      RECT 1.74 2.765 1.91 2.935 ;
      RECT 1.74 5.945 1.91 6.115 ;
      RECT 0.195 1.415 0.365 1.585 ;
      RECT 0.195 4.135 0.365 4.305 ;
      RECT -0.06 2.775 0.11 2.945 ;
      RECT -0.265 1.415 -0.095 1.585 ;
      RECT -0.265 4.135 -0.095 4.305 ;
      RECT -0.54 1.935 -0.37 2.105 ;
      RECT -0.725 1.415 -0.555 1.585 ;
      RECT -0.725 4.135 -0.555 4.305 ;
      RECT -0.78 2.495 -0.61 2.665 ;
      RECT -1.185 1.415 -1.015 1.585 ;
      RECT -1.185 4.135 -1.015 4.305 ;
      RECT -1.26 2.495 -1.09 2.665 ;
      RECT -1.5 1.935 -1.33 2.105 ;
      RECT -1.5 3.615 -1.33 3.785 ;
      RECT -1.645 1.415 -1.475 1.585 ;
      RECT -1.645 4.135 -1.475 4.305 ;
      RECT -2.02 2.775 -1.85 2.945 ;
      RECT -2.105 1.415 -1.935 1.585 ;
      RECT -2.105 4.135 -1.935 4.305 ;
      RECT -2.26 2.215 -2.09 2.385 ;
      RECT -2.5 3.615 -2.33 3.785 ;
      RECT -2.565 1.415 -2.395 1.585 ;
      RECT -2.565 4.135 -2.395 4.305 ;
      RECT -2.74 2.775 -2.57 2.945 ;
      RECT -3.025 1.415 -2.855 1.585 ;
      RECT -3.025 4.135 -2.855 4.305 ;
      RECT -3.22 2.495 -3.05 2.665 ;
      RECT -3.485 1.415 -3.315 1.585 ;
      RECT -3.485 4.135 -3.315 4.305 ;
      RECT -3.7 2.495 -3.53 2.665 ;
      RECT -3.94 1.935 -3.77 2.105 ;
      RECT -3.945 1.415 -3.775 1.585 ;
      RECT -3.945 4.135 -3.775 4.305 ;
      RECT -4.405 1.415 -4.235 1.585 ;
      RECT -4.405 4.135 -4.235 4.305 ;
      RECT -4.7 2.215 -4.53 2.385 ;
      RECT -4.865 1.415 -4.695 1.585 ;
      RECT -4.865 4.135 -4.695 4.305 ;
      RECT -4.94 3.335 -4.77 3.505 ;
      RECT -5.18 2.775 -5.01 2.945 ;
      RECT -5.325 1.415 -5.155 1.585 ;
      RECT -5.325 4.135 -5.155 4.305 ;
      RECT -5.66 2.495 -5.49 2.665 ;
      RECT -5.785 1.415 -5.615 1.585 ;
      RECT -5.785 4.135 -5.615 4.305 ;
      RECT -5.9 1.935 -5.73 2.105 ;
      RECT -5.9 3.335 -5.73 3.505 ;
      RECT -6.245 1.415 -6.075 1.585 ;
      RECT -6.245 4.135 -6.075 4.305 ;
      RECT -6.38 3.055 -6.21 3.225 ;
      RECT -6.705 1.415 -6.535 1.585 ;
      RECT -6.705 4.135 -6.535 4.305 ;
      RECT -6.9 2.495 -6.73 2.665 ;
      RECT -7.14 3.335 -6.97 3.505 ;
      RECT -7.165 1.415 -6.995 1.585 ;
      RECT -7.165 4.135 -6.995 4.305 ;
      RECT -7.38 1.935 -7.21 2.105 ;
      RECT -7.62 2.495 -7.45 2.665 ;
      RECT -7.62 3.055 -7.45 3.225 ;
      RECT -7.625 1.415 -7.455 1.585 ;
      RECT -7.625 4.135 -7.455 4.305 ;
      RECT -8.085 1.415 -7.915 1.585 ;
      RECT -8.085 4.135 -7.915 4.305 ;
      RECT -8.34 1.935 -8.17 2.105 ;
      RECT -8.34 3.615 -8.17 3.785 ;
      RECT -8.545 1.415 -8.375 1.585 ;
      RECT -8.545 4.135 -8.375 4.305 ;
      RECT -8.82 3.055 -8.65 3.225 ;
      RECT -9.005 1.415 -8.835 1.585 ;
      RECT -9.005 4.135 -8.835 4.305 ;
    LAYER li ;
      RECT -1.02 0 -0.85 2.085 ;
      RECT -2.98 0 -2.81 2.085 ;
      RECT -5.42 0 -5.25 2.085 ;
      RECT -6.38 0 -6.21 2.085 ;
      RECT -6.9 0 -6.73 2.085 ;
      RECT -7.86 0 -7.69 2.085 ;
      RECT -8.82 0 -8.65 2.085 ;
      RECT -3.05 0 -2.81 1.595 ;
      RECT -4.6 0 -4.405 1.595 ;
      RECT -6.725 0 -6.53 1.595 ;
      RECT -9.025 0 -8.83 1.595 ;
      RECT -9.15 0 0.665 1.585 ;
      RECT 5.465 0 5.635 0.935 ;
      RECT 4.475 0 4.645 0.935 ;
      RECT 1.73 0 1.9 0.935 ;
      RECT -9.895 0 6.435 0.305 ;
      RECT 5.465 3.405 5.635 5.475 ;
      RECT 4.475 3.405 4.645 5.475 ;
      RECT 1.73 3.405 1.9 5.475 ;
      RECT -9.895 4.135 6.435 4.745 ;
      RECT -0.06 3.635 0.11 4.745 ;
      RECT -1.02 3.635 -0.85 4.745 ;
      RECT -3.46 3.635 -3.29 4.745 ;
      RECT -4.46 3.635 -4.29 4.745 ;
      RECT -5.42 3.635 -5.25 4.745 ;
      RECT -7.86 3.635 -7.69 4.745 ;
      RECT -9.89 8.575 6.435 8.88 ;
      RECT 5.465 7.945 5.635 8.88 ;
      RECT 4.475 7.945 4.645 8.88 ;
      RECT 1.73 7.945 1.9 8.88 ;
      RECT 5.525 1.74 5.695 2.935 ;
      RECT 5.525 1.74 5.99 1.91 ;
      RECT 5.525 6.97 5.99 7.14 ;
      RECT 5.525 5.945 5.695 7.14 ;
      RECT 4.535 1.74 4.705 2.935 ;
      RECT 4.535 1.74 5 1.91 ;
      RECT 4.535 6.97 5 7.14 ;
      RECT 4.535 5.945 4.705 7.14 ;
      RECT 2.68 2.635 2.85 3.865 ;
      RECT 2.735 0.855 2.905 2.805 ;
      RECT 2.68 0.575 2.85 1.025 ;
      RECT 2.68 7.855 2.85 8.305 ;
      RECT 2.735 6.075 2.905 8.025 ;
      RECT 2.68 5.015 2.85 6.245 ;
      RECT 2.16 0.575 2.33 3.865 ;
      RECT 2.16 2.075 2.565 2.405 ;
      RECT 2.16 1.235 2.565 1.565 ;
      RECT 2.16 5.015 2.33 8.305 ;
      RECT 2.16 7.315 2.565 7.645 ;
      RECT 2.16 6.475 2.565 6.805 ;
      RECT -0.54 1.835 -0.37 2.105 ;
      RECT -0.54 1.835 0.19 2.005 ;
      RECT -0.06 2.575 0.11 2.945 ;
      RECT -0.38 2.575 0.11 2.745 ;
      RECT -0.62 3.225 -0.29 3.395 ;
      RECT -1.38 3.055 -0.37 3.225 ;
      RECT -1.38 2.575 -1.21 3.225 ;
      RECT -1.26 2.495 -1.09 2.825 ;
      RECT -2.1 3.225 -1.77 3.395 ;
      RECT -4.02 3.225 -2.73 3.395 ;
      RECT -2.98 3.14 -1.85 3.31 ;
      RECT -2.26 2.215 -1.85 2.385 ;
      RECT -2.02 1.755 -1.85 2.385 ;
      RECT -2.02 2.575 -1.85 2.945 ;
      RECT -2.34 2.575 -1.85 2.745 ;
      RECT -4.78 2.575 -3.45 2.745 ;
      RECT -3.7 2.495 -3.53 2.745 ;
      RECT -4.7 2.175 -4.53 2.385 ;
      RECT -4.7 2.175 -4.21 2.345 ;
      RECT -6.02 3.335 -5.73 3.505 ;
      RECT -6.02 2.575 -5.85 3.505 ;
      RECT -6.22 2.575 -5.85 2.745 ;
      RECT -7.22 2.575 -6.73 2.745 ;
      RECT -6.9 2.495 -6.73 2.745 ;
      RECT -7.14 3.335 -6.73 3.505 ;
      RECT -6.9 3.145 -6.73 3.505 ;
      RECT -8.1 3.055 -7.45 3.225 ;
      RECT -8.1 2.495 -7.93 3.225 ;
      RECT -8.46 3.615 -8.17 3.785 ;
      RECT -8.46 2.575 -8.29 3.785 ;
      RECT -8.66 2.575 -8.29 2.745 ;
      RECT 5.895 0.575 6.065 1.085 ;
      RECT 5.895 2.395 6.065 3.865 ;
      RECT 5.895 5.015 6.065 6.485 ;
      RECT 5.895 7.795 6.065 8.305 ;
      RECT 4.905 0.575 5.075 1.085 ;
      RECT 4.905 2.395 5.075 3.865 ;
      RECT 4.905 5.015 5.075 6.485 ;
      RECT 4.905 7.795 5.075 8.305 ;
      RECT 3.54 0.575 3.71 3.865 ;
      RECT 3.54 5.015 3.71 8.305 ;
      RECT 3.11 0.575 3.28 1.085 ;
      RECT 3.11 1.655 3.28 3.865 ;
      RECT 3.11 5.015 3.28 7.225 ;
      RECT 3.11 7.795 3.28 8.305 ;
      RECT 1.74 1.66 1.91 2.935 ;
      RECT 1.74 5.945 1.91 7.22 ;
      RECT -0.78 2.495 -0.61 2.825 ;
      RECT -1.5 1.755 -1.33 2.105 ;
      RECT -1.5 3.485 -1.33 3.815 ;
      RECT -2.5 3.485 -2.33 3.815 ;
      RECT -2.74 2.495 -2.57 2.945 ;
      RECT -3.22 2.495 -3.05 2.825 ;
      RECT -3.94 1.755 -3.77 2.105 ;
      RECT -4.94 3.145 -4.77 3.505 ;
      RECT -5.18 2.495 -5.01 2.945 ;
      RECT -5.66 2.495 -5.49 2.825 ;
      RECT -5.9 1.755 -5.73 2.105 ;
      RECT -6.38 3.055 -6.21 3.475 ;
      RECT -7.38 1.755 -7.21 2.105 ;
      RECT -7.62 2.495 -7.45 2.825 ;
      RECT -8.34 1.755 -8.17 2.105 ;
      RECT -8.82 3.055 -8.65 3.475 ;
  END
END sky130_osu_single_mpr2ea_8

MACRO sky130_osu_single_mpr2et_8
  CLASS CORE ;
  ORIGIN 12.13 0 ;
  FOREIGN sky130_osu_single_mpr2et_8 -12.13 0 ;
  SIZE 18.565 BY 8.88 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT -2.075 3.535 -1.52 3.865 ;
      RECT -2.075 1.87 -1.775 3.865 ;
      RECT -6.01 2.975 -5.455 3.305 ;
      RECT -5.755 1.87 -5.455 3.305 ;
      RECT -5.755 1.87 -1.775 2.17 ;
      RECT -0.89 1.855 -0.16 2.185 ;
      RECT -3.11 3.535 -2.38 3.865 ;
      RECT -4.81 3.535 -4.08 3.865 ;
      RECT -7.25 2.415 -6.52 2.745 ;
      RECT -8.69 2.975 -7.96 3.305 ;
      RECT -9.765 2.415 -9.035 2.745 ;
      RECT -10.8 2.415 -10.07 2.745 ;
      RECT -11.13 3.535 -10.4 3.865 ;
    LAYER via2 ;
      RECT -0.825 1.92 -0.625 2.12 ;
      RECT -1.785 3.6 -1.585 3.8 ;
      RECT -2.785 3.6 -2.585 3.8 ;
      RECT -4.745 3.6 -4.545 3.8 ;
      RECT -5.945 3.04 -5.745 3.24 ;
      RECT -7.185 2.48 -6.985 2.68 ;
      RECT -8.625 3.04 -8.425 3.24 ;
      RECT -9.365 2.48 -9.165 2.68 ;
      RECT -10.585 2.48 -10.385 2.68 ;
      RECT -11.065 3.6 -10.865 3.8 ;
    LAYER met2 ;
      RECT 2.705 6.28 3.025 6.605 ;
      RECT 2.735 5.695 2.905 6.605 ;
      RECT 2.735 5.695 2.91 6.045 ;
      RECT 2.735 5.695 3.71 5.87 ;
      RECT 3.535 1.965 3.71 5.87 ;
      RECT -9.655 2.98 -9.395 3.3 ;
      RECT -9.715 2.51 -9.575 3.21 ;
      RECT -9.405 2.395 -9.125 2.765 ;
      RECT -7.935 2.42 -7.675 2.74 ;
      RECT -9.715 2.51 -7.675 2.65 ;
      RECT -9.31 1.32 -9.14 2.765 ;
      RECT 3.48 1.965 3.83 2.315 ;
      RECT 1.425 2.04 3.83 2.195 ;
      RECT 1.435 2.025 3.83 2.195 ;
      RECT 1.435 1.32 1.605 2.195 ;
      RECT -9.31 1.32 1.605 1.49 ;
      RECT 3.505 6.655 3.83 6.98 ;
      RECT 2.39 6.745 3.83 6.915 ;
      RECT 2.39 2.395 2.55 6.915 ;
      RECT 2.705 2.365 3.025 2.685 ;
      RECT 2.39 2.395 3.025 2.565 ;
      RECT 1.655 5.845 1.995 6.195 ;
      RECT 1.74 2.705 1.91 6.195 ;
      RECT 1.665 2.705 2.005 3.055 ;
      RECT -4.75 4.135 1.36 4.325 ;
      RECT 1.19 3.145 1.36 4.325 ;
      RECT 1.17 3.15 1.36 4.325 ;
      RECT -4.75 3.515 -4.56 4.325 ;
      RECT -4.785 3.515 -4.505 3.885 ;
      RECT -4.715 3.07 -4.575 4.325 ;
      RECT 1.1 3.15 1.44 3.5 ;
      RECT -4.905 2.955 -4.625 3.325 ;
      RECT -5.195 3.07 -4.575 3.21 ;
      RECT -5.195 1.86 -5.055 3.21 ;
      RECT -5.255 1.86 -4.995 2.18 ;
      RECT -2.295 2.98 -2.035 3.3 ;
      RECT -2.235 1.86 -2.095 3.3 ;
      RECT -2.295 1.86 -2.035 2.18 ;
      RECT -3.295 3.54 -3.035 3.86 ;
      RECT -3.295 2.955 -3.095 3.86 ;
      RECT -3.355 1.86 -3.215 3.49 ;
      RECT -3.355 2.955 -2.855 3.325 ;
      RECT -3.415 1.86 -3.155 2.18 ;
      RECT -3.775 3.54 -3.515 3.86 ;
      RECT -3.715 1.95 -3.575 3.86 ;
      RECT -4.015 1.95 -3.575 2.18 ;
      RECT -4.015 1.86 -3.755 2.18 ;
      RECT -4.255 2.42 -3.995 2.74 ;
      RECT -4.835 2.51 -3.995 2.65 ;
      RECT -4.835 1.57 -4.695 2.65 ;
      RECT -8.175 1.86 -7.915 2.18 ;
      RECT -8.175 1.95 -7.135 2.09 ;
      RECT -7.275 1.57 -7.135 2.09 ;
      RECT -7.275 1.57 -4.695 1.71 ;
      RECT -5.985 2.955 -5.705 3.325 ;
      RECT -5.915 1.86 -5.775 3.325 ;
      RECT -5.975 1.86 -5.715 2.18 ;
      RECT -6.335 3.54 -6.075 3.86 ;
      RECT -6.275 1.95 -6.135 3.86 ;
      RECT -6.695 1.86 -6.435 2.18 ;
      RECT -6.695 1.95 -6.135 2.09 ;
      RECT -8.665 2.955 -8.385 3.325 ;
      RECT -6.695 2.98 -6.435 3.3 ;
      RECT -9.015 2.98 -8.385 3.3 ;
      RECT -9.015 3.07 -6.435 3.21 ;
      RECT -7.225 2.395 -6.945 2.765 ;
      RECT -7.225 2.42 -6.695 2.74 ;
      RECT -10.135 2.98 -9.875 3.3 ;
      RECT -10.075 1.86 -9.935 3.3 ;
      RECT -10.135 1.86 -9.875 2.18 ;
      RECT -11.105 3.515 -10.825 3.885 ;
      RECT -11.095 3.26 -10.835 3.885 ;
      RECT -0.865 1.835 -0.585 2.205 ;
      RECT -1.825 3.515 -1.545 3.885 ;
      RECT -2.825 3.515 -2.545 3.885 ;
      RECT -10.625 2.395 -10.345 2.765 ;
    LAYER via1 ;
      RECT 3.595 6.74 3.745 6.89 ;
      RECT 3.58 2.065 3.73 2.215 ;
      RECT 2.79 2.45 2.94 2.6 ;
      RECT 2.79 6.37 2.94 6.52 ;
      RECT 1.765 2.805 1.915 2.955 ;
      RECT 1.755 5.945 1.905 6.095 ;
      RECT 1.2 3.25 1.35 3.4 ;
      RECT -0.8 1.945 -0.65 2.095 ;
      RECT -1.76 3.625 -1.61 3.775 ;
      RECT -2.24 1.945 -2.09 2.095 ;
      RECT -2.24 3.065 -2.09 3.215 ;
      RECT -2.76 3.625 -2.61 3.775 ;
      RECT -3.24 3.625 -3.09 3.775 ;
      RECT -3.36 1.945 -3.21 2.095 ;
      RECT -3.72 3.625 -3.57 3.775 ;
      RECT -3.96 1.945 -3.81 2.095 ;
      RECT -4.2 2.505 -4.05 2.655 ;
      RECT -4.72 3.625 -4.57 3.775 ;
      RECT -5.2 1.945 -5.05 2.095 ;
      RECT -5.92 1.945 -5.77 2.095 ;
      RECT -5.92 3.065 -5.77 3.215 ;
      RECT -6.28 3.625 -6.13 3.775 ;
      RECT -6.64 1.945 -6.49 2.095 ;
      RECT -6.64 3.065 -6.49 3.215 ;
      RECT -6.9 2.505 -6.75 2.655 ;
      RECT -7.88 2.505 -7.73 2.655 ;
      RECT -8.12 1.945 -7.97 2.095 ;
      RECT -8.96 3.065 -8.81 3.215 ;
      RECT -9.6 3.065 -9.45 3.215 ;
      RECT -10.08 1.945 -9.93 2.095 ;
      RECT -10.08 3.065 -9.93 3.215 ;
      RECT -10.56 2.505 -10.41 2.655 ;
      RECT -11.04 3.345 -10.89 3.495 ;
    LAYER met1 ;
      RECT -11.38 0 0.58 1.74 ;
      RECT -11.38 0 0.665 1.585 ;
      RECT -12.13 0 6.435 0.305 ;
      RECT -12.125 4.145 -9.66 4.75 ;
      RECT -11.38 4.135 6.435 4.745 ;
      RECT -11.38 3.98 0.58 4.745 ;
      RECT 5.835 2.365 6.125 2.595 ;
      RECT 5.895 0.885 6.065 2.595 ;
      RECT 5.835 0.885 6.125 1.115 ;
      RECT 5.835 7.765 6.125 7.995 ;
      RECT 5.895 6.285 6.065 7.995 ;
      RECT 5.835 6.285 6.125 6.515 ;
      RECT 5.425 2.735 5.755 2.965 ;
      RECT 5.425 2.765 5.925 2.935 ;
      RECT 5.425 2.395 5.615 2.965 ;
      RECT 4.845 2.365 5.135 2.595 ;
      RECT 4.845 2.395 5.615 2.565 ;
      RECT 4.905 0.885 5.075 2.595 ;
      RECT 4.845 0.885 5.135 1.115 ;
      RECT 4.845 7.765 5.135 7.995 ;
      RECT 4.905 6.285 5.075 7.995 ;
      RECT 4.845 6.285 5.135 6.515 ;
      RECT 4.845 6.325 5.695 6.485 ;
      RECT 5.525 5.915 5.695 6.485 ;
      RECT 4.845 6.32 5.235 6.485 ;
      RECT 5.465 5.915 5.755 6.145 ;
      RECT 5.465 5.945 5.925 6.115 ;
      RECT 4.475 2.735 4.765 2.965 ;
      RECT 4.475 2.765 4.935 2.935 ;
      RECT 4.535 1.655 4.7 2.965 ;
      RECT 3.05 1.625 3.34 1.855 ;
      RECT 3.05 1.655 4.7 1.825 ;
      RECT 3.11 0.885 3.28 1.855 ;
      RECT 3.05 0.885 3.34 1.115 ;
      RECT 3.05 7.765 3.34 7.995 ;
      RECT 3.11 7.025 3.28 7.995 ;
      RECT 3.11 7.12 4.7 7.29 ;
      RECT 4.53 5.915 4.7 7.29 ;
      RECT 3.05 7.025 3.34 7.255 ;
      RECT 4.475 5.915 4.765 6.145 ;
      RECT 4.475 5.945 4.935 6.115 ;
      RECT 3.48 1.965 3.83 2.315 ;
      RECT 3.31 2.025 3.83 2.195 ;
      RECT 3.505 6.655 3.83 6.98 ;
      RECT 3.48 6.655 3.83 6.885 ;
      RECT 3.31 6.685 3.83 6.855 ;
      RECT 1.1 3.15 1.44 3.5 ;
      RECT 1.19 2.395 1.36 3.5 ;
      RECT 2.705 2.365 3.025 2.685 ;
      RECT 2.675 2.365 3.025 2.595 ;
      RECT 1.19 2.395 3.025 2.565 ;
      RECT 2.705 6.28 3.025 6.605 ;
      RECT 2.675 6.285 3.025 6.515 ;
      RECT 2.505 6.315 3.025 6.485 ;
      RECT 1.665 2.705 2.005 3.055 ;
      RECT 1.665 2.765 2.14 2.935 ;
      RECT 1.655 5.845 1.995 6.195 ;
      RECT 1.655 5.945 2.14 6.115 ;
      RECT -1.845 3.57 -1.525 3.83 ;
      RECT -0.555 2.745 -0.415 3.605 ;
      RECT -1.755 3.465 -0.415 3.605 ;
      RECT -1.755 3.025 -1.615 3.83 ;
      RECT -1.83 3.025 -1.54 3.255 ;
      RECT -0.63 2.745 -0.34 2.975 ;
      RECT -1.11 3.025 -0.82 3.255 ;
      RECT -0.915 1.95 -0.775 3.21 ;
      RECT -0.885 1.89 -0.565 2.15 ;
      RECT -4.285 2.45 -3.965 2.71 ;
      RECT -1.59 2.465 -1.3 2.695 ;
      RECT -4.195 2.37 -1.375 2.51 ;
      RECT -2.325 1.89 -2.005 2.15 ;
      RECT -1.83 1.905 -1.54 2.135 ;
      RECT -2.325 1.95 -1.54 2.09 ;
      RECT -2.325 3.01 -2.005 3.27 ;
      RECT -2.325 2.79 -2.095 3.27 ;
      RECT -2.83 2.745 -2.54 2.975 ;
      RECT -2.83 2.79 -2.095 2.93 ;
      RECT -3.805 3.57 -3.485 3.83 ;
      RECT -4.27 3.585 -3.98 3.815 ;
      RECT -4.27 3.63 -3.485 3.77 ;
      RECT -5.51 2.465 -5.22 2.695 ;
      RECT -5.51 2.51 -4.575 2.65 ;
      RECT -4.715 1.95 -4.575 2.65 ;
      RECT -4.045 1.89 -3.725 2.15 ;
      RECT -4.27 1.905 -3.725 2.135 ;
      RECT -4.715 1.95 -3.725 2.09 ;
      RECT -6.365 3.57 -6.045 3.83 ;
      RECT -6.365 3.63 -5.295 3.77 ;
      RECT -5.435 3.07 -5.295 3.77 ;
      RECT -4.27 3.025 -3.98 3.255 ;
      RECT -5.435 3.07 -3.98 3.21 ;
      RECT -6.005 1.89 -5.685 2.15 ;
      RECT -6.23 1.905 -5.685 2.135 ;
      RECT -6.985 2.45 -6.665 2.71 ;
      RECT -5.99 2.465 -5.7 2.695 ;
      RECT -7.23 2.465 -6.665 2.695 ;
      RECT -7.23 2.51 -5.7 2.65 ;
      RECT -7.71 3.025 -7.42 3.255 ;
      RECT -7.515 1.95 -7.375 3.21 ;
      RECT -6.725 1.89 -6.405 2.15 ;
      RECT -7.71 1.905 -7.42 2.135 ;
      RECT -7.71 1.95 -6.405 2.09 ;
      RECT -8.115 3.465 -7.015 3.605 ;
      RECT -7.23 3.305 -6.94 3.535 ;
      RECT -8.19 3.305 -7.9 3.535 ;
      RECT -7.95 2.37 -7.66 2.74 ;
      RECT -8.715 2.37 -7.66 2.51 ;
      RECT -8.205 1.89 -7.885 2.15 ;
      RECT -10.165 1.89 -9.845 2.15 ;
      RECT -10.165 1.95 -7.885 2.09 ;
      RECT -9.045 3.01 -8.725 3.27 ;
      RECT -9.045 3.01 -8.215 3.15 ;
      RECT -8.43 2.745 -8.215 3.15 ;
      RECT -8.43 2.745 -8.14 2.975 ;
      RECT -10.645 2.45 -10.325 2.71 ;
      RECT -9.235 2.465 -8.945 2.695 ;
      RECT -10.645 2.465 -10.1 2.695 ;
      RECT -10.645 2.55 -9.695 2.69 ;
      RECT -9.835 2.37 -9.695 2.69 ;
      RECT -9.335 2.465 -8.945 2.65 ;
      RECT -9.835 2.37 -9.195 2.51 ;
      RECT -11.125 3.26 -10.805 3.675 ;
      RECT -11.045 1.905 -10.89 3.675 ;
      RECT -11.11 1.905 -10.82 2.135 ;
      RECT -12.125 8.575 6.435 8.88 ;
      RECT -0.3 2.735 0.02 3.055 ;
      RECT -2.845 3.57 -2.525 3.83 ;
      RECT -3.445 1.89 -2.765 2.15 ;
      RECT -3.325 3.57 -3.005 3.83 ;
      RECT -4.805 3.57 -4.485 3.83 ;
      RECT -5.285 1.89 -4.965 2.15 ;
      RECT -6.005 3.01 -5.685 3.27 ;
      RECT -6.725 3.01 -6.405 3.27 ;
      RECT -9.685 3.01 -9.365 3.27 ;
      RECT -10.165 3.01 -9.845 3.27 ;
    LAYER mcon ;
      RECT 5.895 0.915 6.065 1.085 ;
      RECT 5.895 2.395 6.065 2.565 ;
      RECT 5.895 6.315 6.065 6.485 ;
      RECT 5.895 7.795 6.065 7.965 ;
      RECT 5.545 0.105 5.715 0.275 ;
      RECT 5.545 4.165 5.715 4.335 ;
      RECT 5.545 4.545 5.715 4.715 ;
      RECT 5.545 8.605 5.715 8.775 ;
      RECT 5.525 2.765 5.695 2.935 ;
      RECT 5.525 5.945 5.695 6.115 ;
      RECT 4.905 0.915 5.075 1.085 ;
      RECT 4.905 2.395 5.075 2.565 ;
      RECT 4.905 6.315 5.075 6.485 ;
      RECT 4.905 7.795 5.075 7.965 ;
      RECT 4.555 0.105 4.725 0.275 ;
      RECT 4.555 4.165 4.725 4.335 ;
      RECT 4.555 4.545 4.725 4.715 ;
      RECT 4.555 8.605 4.725 8.775 ;
      RECT 4.535 2.765 4.705 2.935 ;
      RECT 4.535 5.945 4.705 6.115 ;
      RECT 3.85 0.105 4.02 0.275 ;
      RECT 3.85 4.165 4.02 4.335 ;
      RECT 3.85 4.545 4.02 4.715 ;
      RECT 3.85 8.605 4.02 8.775 ;
      RECT 3.54 2.025 3.71 2.195 ;
      RECT 3.54 6.685 3.71 6.855 ;
      RECT 3.17 0.105 3.34 0.275 ;
      RECT 3.17 8.605 3.34 8.775 ;
      RECT 3.11 0.915 3.28 1.085 ;
      RECT 3.11 1.655 3.28 1.825 ;
      RECT 3.11 7.055 3.28 7.225 ;
      RECT 3.11 7.795 3.28 7.965 ;
      RECT 2.735 2.395 2.905 2.565 ;
      RECT 2.735 6.315 2.905 6.485 ;
      RECT 2.49 0.105 2.66 0.275 ;
      RECT 2.49 8.605 2.66 8.775 ;
      RECT 1.81 0.105 1.98 0.275 ;
      RECT 1.81 8.605 1.98 8.775 ;
      RECT 1.74 2.765 1.91 2.935 ;
      RECT 1.74 5.945 1.91 6.115 ;
      RECT 0.265 1.415 0.435 1.585 ;
      RECT 0.265 4.135 0.435 4.305 ;
      RECT -0.195 1.415 -0.025 1.585 ;
      RECT -0.195 4.135 -0.025 4.305 ;
      RECT -0.57 2.775 -0.4 2.945 ;
      RECT -0.655 1.415 -0.485 1.585 ;
      RECT -0.655 4.135 -0.485 4.305 ;
      RECT -0.81 1.935 -0.64 2.105 ;
      RECT -1.05 3.055 -0.88 3.225 ;
      RECT -1.115 1.415 -0.945 1.585 ;
      RECT -1.115 4.135 -0.945 4.305 ;
      RECT -1.53 2.495 -1.36 2.665 ;
      RECT -1.575 1.415 -1.405 1.585 ;
      RECT -1.575 4.135 -1.405 4.305 ;
      RECT -1.77 1.935 -1.6 2.105 ;
      RECT -1.77 3.055 -1.6 3.225 ;
      RECT -1.77 3.615 -1.6 3.785 ;
      RECT -2.035 1.415 -1.865 1.585 ;
      RECT -2.035 4.135 -1.865 4.305 ;
      RECT -2.25 3.055 -2.08 3.225 ;
      RECT -2.495 1.415 -2.325 1.585 ;
      RECT -2.495 4.135 -2.325 4.305 ;
      RECT -2.77 2.775 -2.6 2.945 ;
      RECT -2.77 3.615 -2.6 3.785 ;
      RECT -2.955 1.415 -2.785 1.585 ;
      RECT -2.955 4.135 -2.785 4.305 ;
      RECT -3.25 1.935 -3.08 2.105 ;
      RECT -3.25 3.615 -3.08 3.785 ;
      RECT -3.415 1.415 -3.245 1.585 ;
      RECT -3.415 4.135 -3.245 4.305 ;
      RECT -3.875 1.415 -3.705 1.585 ;
      RECT -3.875 4.135 -3.705 4.305 ;
      RECT -4.21 1.935 -4.04 2.105 ;
      RECT -4.21 2.495 -4.04 2.665 ;
      RECT -4.21 3.055 -4.04 3.225 ;
      RECT -4.21 3.615 -4.04 3.785 ;
      RECT -4.335 1.415 -4.165 1.585 ;
      RECT -4.335 4.135 -4.165 4.305 ;
      RECT -4.73 3.615 -4.56 3.785 ;
      RECT -4.795 1.415 -4.625 1.585 ;
      RECT -4.795 4.135 -4.625 4.305 ;
      RECT -5.21 1.935 -5.04 2.105 ;
      RECT -5.255 1.415 -5.085 1.585 ;
      RECT -5.255 4.135 -5.085 4.305 ;
      RECT -5.45 2.495 -5.28 2.665 ;
      RECT -5.715 1.415 -5.545 1.585 ;
      RECT -5.715 4.135 -5.545 4.305 ;
      RECT -5.93 2.495 -5.76 2.665 ;
      RECT -5.93 3.055 -5.76 3.225 ;
      RECT -6.17 1.935 -6 2.105 ;
      RECT -6.175 1.415 -6.005 1.585 ;
      RECT -6.175 4.135 -6.005 4.305 ;
      RECT -6.635 1.415 -6.465 1.585 ;
      RECT -6.635 4.135 -6.465 4.305 ;
      RECT -6.65 3.055 -6.48 3.225 ;
      RECT -7.095 1.415 -6.925 1.585 ;
      RECT -7.095 4.135 -6.925 4.305 ;
      RECT -7.17 2.495 -7 2.665 ;
      RECT -7.17 3.335 -7 3.505 ;
      RECT -7.555 1.415 -7.385 1.585 ;
      RECT -7.555 4.135 -7.385 4.305 ;
      RECT -7.65 1.935 -7.48 2.105 ;
      RECT -7.65 3.055 -7.48 3.225 ;
      RECT -7.89 2.495 -7.72 2.665 ;
      RECT -8.015 1.415 -7.845 1.585 ;
      RECT -8.015 4.135 -7.845 4.305 ;
      RECT -8.13 3.335 -7.96 3.505 ;
      RECT -8.37 2.775 -8.2 2.945 ;
      RECT -8.475 1.415 -8.305 1.585 ;
      RECT -8.475 4.135 -8.305 4.305 ;
      RECT -8.935 1.415 -8.765 1.585 ;
      RECT -8.935 4.135 -8.765 4.305 ;
      RECT -9.175 2.495 -9.005 2.665 ;
      RECT -9.395 1.415 -9.225 1.585 ;
      RECT -9.395 4.135 -9.225 4.305 ;
      RECT -9.61 3.055 -9.44 3.225 ;
      RECT -9.855 1.415 -9.685 1.585 ;
      RECT -9.855 4.135 -9.685 4.305 ;
      RECT -10.09 1.935 -9.92 2.105 ;
      RECT -10.09 3.055 -9.92 3.225 ;
      RECT -10.315 1.415 -10.145 1.585 ;
      RECT -10.315 4.135 -10.145 4.305 ;
      RECT -10.33 2.495 -10.16 2.665 ;
      RECT -10.775 1.415 -10.605 1.585 ;
      RECT -10.775 4.135 -10.605 4.305 ;
      RECT -11.05 1.935 -10.88 2.105 ;
      RECT -11.05 3.475 -10.88 3.645 ;
      RECT -11.235 1.415 -11.065 1.585 ;
      RECT -11.235 4.135 -11.065 4.305 ;
    LAYER li ;
      RECT -0.33 0 -0.16 2.085 ;
      RECT -1.29 0 -1.12 2.085 ;
      RECT -2.25 0 -2.08 2.085 ;
      RECT -2.77 0 -2.6 2.085 ;
      RECT -3.73 0 -3.56 2.085 ;
      RECT -4.73 0 -4.56 2.085 ;
      RECT -5.69 0 -5.52 2.085 ;
      RECT -7.17 0 -7 2.085 ;
      RECT -9.09 0 -8.92 2.085 ;
      RECT -10.57 0 -10.4 2.085 ;
      RECT -3.05 0 -2.855 1.595 ;
      RECT -6.725 0 -6.53 1.595 ;
      RECT -9.09 0 -8.83 1.595 ;
      RECT -11.38 0 0.665 1.585 ;
      RECT 5.465 0 5.635 0.935 ;
      RECT 4.475 0 4.645 0.935 ;
      RECT 1.73 0 1.9 0.935 ;
      RECT -12.13 0 6.435 0.305 ;
      RECT 5.465 3.405 5.635 5.475 ;
      RECT 4.475 3.405 4.645 5.475 ;
      RECT 1.73 3.405 1.9 5.475 ;
      RECT -12.125 4.145 -9.66 4.75 ;
      RECT -11.38 4.135 6.435 4.745 ;
      RECT -1.29 3.635 -1.12 4.745 ;
      RECT -3.73 3.635 -3.56 4.745 ;
      RECT -5.69 3.635 -5.52 4.745 ;
      RECT -6.65 3.635 -6.48 4.745 ;
      RECT -8.61 3.635 -8.44 4.745 ;
      RECT -9.61 3.635 -9.44 4.745 ;
      RECT -10.57 3.635 -10.4 4.75 ;
      RECT -12.125 8.575 6.435 8.88 ;
      RECT 5.465 7.945 5.635 8.88 ;
      RECT 4.475 7.945 4.645 8.88 ;
      RECT 1.73 7.945 1.9 8.88 ;
      RECT 5.525 1.74 5.695 2.935 ;
      RECT 5.525 1.74 5.99 1.91 ;
      RECT 5.525 6.97 5.99 7.14 ;
      RECT 5.525 5.945 5.695 7.14 ;
      RECT 4.535 1.74 4.705 2.935 ;
      RECT 4.535 1.74 5 1.91 ;
      RECT 4.535 6.97 5 7.14 ;
      RECT 4.535 5.945 4.705 7.14 ;
      RECT 2.68 2.635 2.85 3.865 ;
      RECT 2.735 0.855 2.905 2.805 ;
      RECT 2.68 0.575 2.85 1.025 ;
      RECT 2.68 7.855 2.85 8.305 ;
      RECT 2.735 6.075 2.905 8.025 ;
      RECT 2.68 5.015 2.85 6.245 ;
      RECT 2.16 0.575 2.33 3.865 ;
      RECT 2.16 2.075 2.565 2.405 ;
      RECT 2.16 1.235 2.565 1.565 ;
      RECT 2.16 5.015 2.33 8.305 ;
      RECT 2.16 7.315 2.565 7.645 ;
      RECT 2.16 6.475 2.565 6.805 ;
      RECT -1.05 3.225 -0.08 3.395 ;
      RECT -1.05 3.055 -0.88 3.395 ;
      RECT -1.53 2.495 -1.36 2.825 ;
      RECT -1.53 2.575 -0.8 2.745 ;
      RECT -1.89 3.615 -1.6 3.785 ;
      RECT -1.89 2.575 -1.72 3.785 ;
      RECT -1.89 3.055 -1.6 3.225 ;
      RECT -2.09 2.575 -1.72 2.745 ;
      RECT -2.77 2.675 -2.6 2.945 ;
      RECT -3.01 2.675 -2.6 2.845 ;
      RECT -3.09 2.575 -2.76 2.745 ;
      RECT -3.25 3.615 -2.6 3.785 ;
      RECT -2.77 3.145 -2.6 3.785 ;
      RECT -2.89 3.225 -2.6 3.785 ;
      RECT -4.21 2.915 -4.04 3.225 ;
      RECT -4.21 2.915 -3.32 3.085 ;
      RECT -3.49 2.495 -3.32 3.085 ;
      RECT -4.21 2.575 -3.72 2.745 ;
      RECT -4.21 2.495 -4.04 2.745 ;
      RECT -6.25 3.225 -5.76 3.395 ;
      RECT -5.09 2.575 -4.92 3.225 ;
      RECT -5.93 3.055 -4.92 3.225 ;
      RECT -4.97 2.495 -4.8 2.825 ;
      RECT -6.17 1.835 -6 2.105 ;
      RECT -6.73 1.835 -6 2.005 ;
      RECT -6.65 2.575 -6.48 3.225 ;
      RECT -6.65 2.575 -6.16 2.745 ;
      RECT -7.49 2.575 -7 2.745 ;
      RECT -7.17 2.495 -7 2.745 ;
      RECT -7.65 1.835 -7.48 2.105 ;
      RECT -8.21 1.835 -7.48 2.005 ;
      RECT -8.13 3.225 -7.96 3.505 ;
      RECT -9.17 3.225 -7.88 3.395 ;
      RECT -9.175 2.575 -8.6 2.745 ;
      RECT -9.175 2.495 -9.005 2.745 ;
      RECT -10.09 1.835 -9.92 2.105 ;
      RECT -10.09 1.835 -9.36 2.005 ;
      RECT -9.73 3.055 -9.44 3.225 ;
      RECT -9.73 2.575 -9.56 3.225 ;
      RECT -9.93 2.575 -9.56 2.745 ;
      RECT -10.09 3.055 -9.92 3.475 ;
      RECT -10.71 3.14 -9.92 3.31 ;
      RECT -10.71 2.915 -10.54 3.31 ;
      RECT -10.81 2.495 -10.64 3.085 ;
      RECT -11.05 2.575 -10.64 2.845 ;
      RECT 5.895 0.575 6.065 1.085 ;
      RECT 5.895 2.395 6.065 3.865 ;
      RECT 5.895 5.015 6.065 6.485 ;
      RECT 5.895 7.795 6.065 8.305 ;
      RECT 4.905 0.575 5.075 1.085 ;
      RECT 4.905 2.395 5.075 3.865 ;
      RECT 4.905 5.015 5.075 6.485 ;
      RECT 4.905 7.795 5.075 8.305 ;
      RECT 3.54 0.575 3.71 3.865 ;
      RECT 3.54 5.015 3.71 8.305 ;
      RECT 3.11 0.575 3.28 1.085 ;
      RECT 3.11 1.655 3.28 3.865 ;
      RECT 3.11 5.015 3.28 7.225 ;
      RECT 3.11 7.795 3.28 8.305 ;
      RECT 1.74 1.66 1.91 2.935 ;
      RECT 1.74 5.945 1.91 7.22 ;
      RECT -0.57 2.495 -0.4 2.945 ;
      RECT -0.81 1.755 -0.64 2.105 ;
      RECT -1.77 1.755 -1.6 2.105 ;
      RECT -2.25 3.055 -2.08 3.475 ;
      RECT -3.25 1.755 -3.08 2.105 ;
      RECT -4.21 1.755 -4.04 2.105 ;
      RECT -4.21 3.485 -4.04 3.815 ;
      RECT -4.73 3.145 -4.56 3.785 ;
      RECT -5.21 1.755 -5.04 2.105 ;
      RECT -5.45 2.495 -5.28 2.825 ;
      RECT -5.93 2.495 -5.76 2.825 ;
      RECT -7.17 3.145 -7 3.505 ;
      RECT -7.65 3.055 -7.48 3.475 ;
      RECT -7.89 2.495 -7.72 2.825 ;
      RECT -8.37 2.495 -8.2 2.945 ;
      RECT -10.33 2.495 -10.16 2.825 ;
      RECT -11.05 1.755 -10.88 2.105 ;
      RECT -11.05 3.285 -10.88 3.645 ;
  END
END sky130_osu_single_mpr2et_8

MACRO sky130_osu_single_mpr2xa_8
  CLASS CORE ;
  ORIGIN 8.825 0 ;
  FOREIGN sky130_osu_single_mpr2xa_8 -8.825 0 ;
  SIZE 15.26 BY 8.88 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met4 ;
      RECT -5.925 2.975 -5.595 3.305 ;
      RECT -5.91 2.5 -5.595 3.305 ;
      RECT -3.765 2.485 -3.435 2.84 ;
      RECT -5.91 2.5 -3.435 2.8 ;
    LAYER via3 ;
      RECT -3.7 2.575 -3.5 2.775 ;
      RECT -5.86 3.04 -5.66 3.24 ;
    LAYER met3 ;
      RECT -3.285 3.51 -2.955 3.865 ;
      RECT -5.19 3.55 -2.955 3.85 ;
      RECT -5.19 2.415 -4.89 3.85 ;
      RECT -5.205 2.415 -4.875 2.745 ;
      RECT -4.215 2.52 -3.435 2.865 ;
      RECT -3.74 2.485 -3.435 2.865 ;
      RECT -3.76 2.515 -3.435 2.865 ;
      RECT -4.64 1.88 -3.91 2.21 ;
      RECT -4.495 1.06 -4.19 2.21 ;
      RECT -4.525 1.06 -4.15 1.43 ;
      RECT -5.92 2.415 -5.6 3.33 ;
      RECT -5.92 2.415 -5.59 2.95 ;
      RECT -0.365 1.855 0.365 2.185 ;
      RECT -2.055 1.87 -1.325 2.2 ;
      RECT -3.09 1.855 -2.36 2.205 ;
      RECT -7.11 2.975 -6.38 3.305 ;
      RECT -7.245 1.855 -6.515 2.185 ;
    LAYER via2 ;
      RECT -0.13 1.92 0.07 2.12 ;
      RECT -1.99 1.935 -1.79 2.135 ;
      RECT -3.01 1.94 -2.81 2.14 ;
      RECT -3.22 3.575 -3.02 3.775 ;
      RECT -3.7 2.575 -3.5 2.775 ;
      RECT -4.435 1.145 -4.235 1.345 ;
      RECT -4.45 1.945 -4.25 2.145 ;
      RECT -5.14 2.48 -4.94 2.68 ;
      RECT -5.855 2.48 -5.655 2.68 ;
      RECT -6.82 3.04 -6.62 3.24 ;
      RECT -7.06 1.92 -6.86 2.12 ;
    LAYER met2 ;
      RECT 2.705 6.28 3.025 6.605 ;
      RECT 2.735 5.695 2.905 6.605 ;
      RECT 2.735 5.695 2.91 6.045 ;
      RECT 2.735 5.695 3.71 5.87 ;
      RECT 3.535 1.965 3.71 5.87 ;
      RECT 3.48 1.965 3.83 2.315 ;
      RECT -7.1 1.835 -6.82 2.205 ;
      RECT 1.07 2.025 3.83 2.195 ;
      RECT -7.1 1.86 -6.71 2.18 ;
      RECT 1.07 0.745 1.24 2.195 ;
      RECT -6.95 0.745 -6.78 2.18 ;
      RECT -6.95 0.745 1.24 0.915 ;
      RECT 3.505 6.655 3.83 6.98 ;
      RECT 2.39 6.745 3.83 6.915 ;
      RECT 2.39 2.395 2.55 6.915 ;
      RECT 2.705 2.365 3.025 2.685 ;
      RECT 2.39 2.395 3.025 2.565 ;
      RECT 1.66 5.86 2 6.21 ;
      RECT 1.74 2.705 1.91 6.21 ;
      RECT 1.66 2.705 2 3.055 ;
      RECT 1.1 2.7 1.44 3.05 ;
      RECT 0.59 2.77 1.44 2.97 ;
      RECT 0.59 1.18 0.79 2.97 ;
      RECT 1.19 2.695 1.36 3.05 ;
      RECT -4.525 1.06 -4.15 1.43 ;
      RECT -4.525 1.18 0.79 1.38 ;
      RECT -0.16 3.54 0.1 3.86 ;
      RECT -0.1 1.835 0.04 3.86 ;
      RECT -0.275 2.395 0.04 2.765 ;
      RECT -0.205 1.95 0.04 2.765 ;
      RECT -0.17 1.835 0.11 2.205 ;
      RECT -0.85 2.42 -0.59 2.74 ;
      RECT -1.51 2.51 -0.59 2.65 ;
      RECT -1.51 1.57 -1.37 2.65 ;
      RECT -5.05 1.86 -4.79 2.18 ;
      RECT -4.87 1.57 -4.73 2.09 ;
      RECT -4.87 1.57 -1.37 1.71 ;
      RECT -2.02 3.26 -1.76 3.58 ;
      RECT -1.96 1.85 -1.82 3.58 ;
      RECT -2.03 1.85 -1.75 2.22 ;
      RECT -4.63 4.01 -2.195 4.15 ;
      RECT -2.335 2.7 -2.195 4.15 ;
      RECT -4.63 3.63 -4.49 4.15 ;
      RECT -4.93 3.63 -4.49 3.86 ;
      RECT -7.27 3.63 -4.49 3.77 ;
      RECT -4.93 3.54 -4.67 3.86 ;
      RECT -7.27 3.35 -7.13 3.77 ;
      RECT -7.78 3.26 -7.52 3.58 ;
      RECT -7.78 3.35 -7.13 3.49 ;
      RECT -7.72 1.86 -7.58 3.58 ;
      RECT -2.395 2.7 -2.135 3.02 ;
      RECT -7.78 1.86 -7.52 2.18 ;
      RECT -2.77 3.54 -2.51 3.86 ;
      RECT -2.71 1.95 -2.57 3.86 ;
      RECT -3.05 1.95 -2.57 2.225 ;
      RECT -3.25 1.855 -2.77 2.2 ;
      RECT -3.26 3.49 -2.98 3.86 ;
      RECT -3.19 2.395 -3.05 3.86 ;
      RECT -3.25 2.395 -2.99 3.02 ;
      RECT -3.26 2.395 -2.98 2.765 ;
      RECT -4.33 3.54 -4.07 3.86 ;
      RECT -4.33 3.35 -4.13 3.86 ;
      RECT -4.525 3.35 -4.13 3.49 ;
      RECT -4.525 1.86 -4.385 3.49 ;
      RECT -4.525 1.86 -4.21 2.23 ;
      RECT -4.585 1.86 -4.21 2.18 ;
      RECT -6.86 2.955 -6.58 3.325 ;
      RECT -5.41 2.98 -5.15 3.3 ;
      RECT -7.03 3.07 -5.15 3.21 ;
      RECT -7.03 2.955 -6.58 3.21 ;
      RECT -7.09 2.395 -6.83 3.02 ;
      RECT -7.1 2.395 -6.82 2.765 ;
      RECT -6.02 2.395 -5.61 2.765 ;
      RECT -6.61 2.42 -6.35 2.74 ;
      RECT -6.61 2.51 -5.61 2.65 ;
      RECT -3.74 2.395 -3.46 2.86 ;
      RECT -3.98 1.86 -3.7 2.205 ;
      RECT -5.18 2.395 -4.9 2.765 ;
    LAYER via1 ;
      RECT 3.595 6.74 3.745 6.89 ;
      RECT 3.58 2.065 3.73 2.215 ;
      RECT 2.79 2.45 2.94 2.6 ;
      RECT 2.79 6.37 2.94 6.52 ;
      RECT 1.76 2.805 1.91 2.955 ;
      RECT 1.76 5.96 1.91 6.11 ;
      RECT 1.2 2.8 1.35 2.95 ;
      RECT -0.105 1.945 0.045 2.095 ;
      RECT -0.105 3.625 0.045 3.775 ;
      RECT -0.795 2.505 -0.645 2.655 ;
      RECT -1.965 1.945 -1.815 2.095 ;
      RECT -1.965 3.345 -1.815 3.495 ;
      RECT -2.34 2.785 -2.19 2.935 ;
      RECT -2.715 3.625 -2.565 3.775 ;
      RECT -3.195 1.945 -3.045 2.095 ;
      RECT -3.195 2.785 -3.045 2.935 ;
      RECT -3.675 2.505 -3.525 2.655 ;
      RECT -3.915 1.945 -3.765 2.095 ;
      RECT -4.275 3.625 -4.125 3.775 ;
      RECT -4.53 1.945 -4.38 2.095 ;
      RECT -4.875 3.625 -4.725 3.775 ;
      RECT -4.995 1.945 -4.845 2.095 ;
      RECT -5.115 2.505 -4.965 2.655 ;
      RECT -5.355 3.065 -5.205 3.215 ;
      RECT -6.555 2.505 -6.405 2.655 ;
      RECT -6.915 1.945 -6.765 2.095 ;
      RECT -7.035 2.785 -6.885 2.935 ;
      RECT -7.725 1.945 -7.575 2.095 ;
      RECT -7.725 3.345 -7.575 3.495 ;
    LAYER met1 ;
      RECT -8.075 0 0.665 1.74 ;
      RECT -8.825 0 6.435 0.305 ;
      RECT -8.825 4.14 6.435 4.745 ;
      RECT -8.075 4.135 6.435 4.745 ;
      RECT -8.075 3.98 0.665 4.745 ;
      RECT 5.835 2.365 6.125 2.595 ;
      RECT 5.895 0.885 6.065 2.595 ;
      RECT 5.835 0.885 6.125 1.115 ;
      RECT 5.835 7.765 6.125 7.995 ;
      RECT 5.895 6.285 6.065 7.995 ;
      RECT 5.835 6.285 6.125 6.515 ;
      RECT 5.425 2.735 5.755 2.965 ;
      RECT 5.425 2.765 5.925 2.935 ;
      RECT 5.425 2.395 5.615 2.965 ;
      RECT 4.845 2.365 5.135 2.595 ;
      RECT 4.845 2.395 5.615 2.565 ;
      RECT 4.905 0.885 5.075 2.595 ;
      RECT 4.845 0.885 5.135 1.115 ;
      RECT 4.845 7.765 5.135 7.995 ;
      RECT 4.905 6.285 5.075 7.995 ;
      RECT 4.845 6.285 5.135 6.515 ;
      RECT 4.845 6.325 5.695 6.485 ;
      RECT 5.525 5.915 5.695 6.485 ;
      RECT 4.845 6.32 5.235 6.485 ;
      RECT 5.465 5.915 5.755 6.145 ;
      RECT 5.465 5.945 5.925 6.115 ;
      RECT 4.475 2.735 4.765 2.965 ;
      RECT 4.475 2.765 4.935 2.935 ;
      RECT 4.535 1.655 4.7 2.965 ;
      RECT 3.05 1.625 3.34 1.855 ;
      RECT 3.05 1.655 4.7 1.825 ;
      RECT 3.11 0.885 3.28 1.855 ;
      RECT 3.05 0.885 3.34 1.115 ;
      RECT 3.05 7.765 3.34 7.995 ;
      RECT 3.11 7.025 3.28 7.995 ;
      RECT 3.11 7.12 4.7 7.29 ;
      RECT 4.53 5.915 4.7 7.29 ;
      RECT 3.05 7.025 3.34 7.255 ;
      RECT 4.475 5.915 4.765 6.145 ;
      RECT 4.475 5.945 4.935 6.115 ;
      RECT 3.48 1.965 3.83 2.315 ;
      RECT 3.31 2.025 3.83 2.195 ;
      RECT 3.505 6.655 3.83 6.98 ;
      RECT 3.48 6.655 3.83 6.885 ;
      RECT 3.31 6.685 3.83 6.855 ;
      RECT 1.1 2.7 1.44 3.05 ;
      RECT 1.19 2.395 1.36 3.05 ;
      RECT 2.705 2.365 3.025 2.685 ;
      RECT 2.675 2.365 3.025 2.595 ;
      RECT 1.19 2.395 3.025 2.565 ;
      RECT 2.705 6.28 3.025 6.605 ;
      RECT 2.675 6.285 3.025 6.515 ;
      RECT 2.505 6.315 3.025 6.485 ;
      RECT 1.66 2.705 2 3.055 ;
      RECT 1.66 2.765 2.14 2.935 ;
      RECT 1.66 5.86 2 6.21 ;
      RECT 1.66 5.945 2.14 6.115 ;
      RECT -0.19 1.89 0.13 2.15 ;
      RECT -0.625 1.905 -0.335 2.135 ;
      RECT -0.625 1.95 0.13 2.09 ;
      RECT -0.19 3.57 0.13 3.83 ;
      RECT -0.625 3.585 -0.335 3.815 ;
      RECT -0.625 3.63 0.13 3.77 ;
      RECT -0.865 3.025 -0.575 3.255 ;
      RECT -0.865 3.07 -0.29 3.21 ;
      RECT -0.43 2.93 -0.17 3.07 ;
      RECT -0.385 2.745 -0.29 3.21 ;
      RECT -0.3 2.735 0.02 3.055 ;
      RECT -2.23 2.93 -1.13 3.07 ;
      RECT -2.425 2.73 -2.105 2.99 ;
      RECT -1.345 2.745 -1.055 2.975 ;
      RECT -2.425 2.745 -2.015 2.99 ;
      RECT -2.05 1.89 -1.73 2.15 ;
      RECT -1.585 1.905 -1.295 2.135 ;
      RECT -2.05 1.95 -1.295 2.09 ;
      RECT -4.75 3.155 -2.57 3.295 ;
      RECT -2.71 2.165 -2.57 3.295 ;
      RECT -4.75 3.07 -3.455 3.295 ;
      RECT -3.745 3.025 -3.455 3.295 ;
      RECT -4.75 2.79 -4.415 3.295 ;
      RECT -4.705 2.745 -4.415 3.295 ;
      RECT -1.825 2.465 -1.535 2.695 ;
      RECT -2.71 2.37 -1.61 2.51 ;
      RECT -2.785 2.165 -2.495 2.415 ;
      RECT -2.8 3.57 -2.48 3.83 ;
      RECT -2.8 3.585 -2.285 3.815 ;
      RECT -4.225 2.465 -3.935 2.695 ;
      RECT -4.075 2.07 -3.935 2.695 ;
      RECT -4.075 2.07 -3.77 2.21 ;
      RECT -3.28 1.89 -2.96 2.15 ;
      RECT -4 1.89 -3.68 2.15 ;
      RECT -3.505 1.905 -2.96 2.135 ;
      RECT -4 1.95 -2.96 2.09 ;
      RECT -4.36 3.57 -4.04 3.83 ;
      RECT -4.465 3.585 -4.04 3.815 ;
      RECT -6.385 3.025 -6.095 3.255 ;
      RECT -6.385 3.025 -5.93 3.21 ;
      RECT -6.07 2.55 -5.93 3.21 ;
      RECT -5.95 1.95 -5.81 2.69 ;
      RECT -5.08 1.89 -4.76 2.15 ;
      RECT -5.905 1.905 -5.615 2.135 ;
      RECT -5.95 1.95 -4.76 2.09 ;
      RECT -5.2 2.45 -4.88 2.71 ;
      RECT -5.665 2.465 -5.375 2.695 ;
      RECT -5.665 2.51 -4.88 2.65 ;
      RECT -5.44 3.01 -5.12 3.27 ;
      RECT -5.44 3.025 -4.895 3.255 ;
      RECT -5.905 3.585 -5.615 3.815 ;
      RECT -6.79 3.465 -5.69 3.605 ;
      RECT -6.865 3.305 -6.575 3.535 ;
      RECT -7.585 2.745 -7.295 2.975 ;
      RECT -7.51 2.37 -7.37 2.975 ;
      RECT -7.51 2.37 -6.89 2.51 ;
      RECT -7.03 1.95 -6.89 2.51 ;
      RECT -7.27 1.95 -6.89 2.21 ;
      RECT -7 1.89 -6.68 2.15 ;
      RECT -6.385 1.905 -6.095 2.135 ;
      RECT -7.27 1.95 -6.095 2.09 ;
      RECT -8.825 8.575 6.435 8.88 ;
      RECT -0.88 2.45 -0.56 2.71 ;
      RECT -2.05 3.29 -1.73 3.55 ;
      RECT -3.28 2.73 -2.96 2.99 ;
      RECT -3.76 2.45 -3.44 2.71 ;
      RECT -4.615 1.89 -4.215 2.15 ;
      RECT -4.96 3.57 -4.64 3.83 ;
      RECT -6.64 2.45 -6.32 2.71 ;
      RECT -7.12 2.73 -6.8 2.99 ;
      RECT -7.81 1.89 -7.49 2.15 ;
      RECT -7.81 3.29 -7.49 3.55 ;
    LAYER mcon ;
      RECT 5.895 0.915 6.065 1.085 ;
      RECT 5.895 2.395 6.065 2.565 ;
      RECT 5.895 6.315 6.065 6.485 ;
      RECT 5.895 7.795 6.065 7.965 ;
      RECT 5.545 0.105 5.715 0.275 ;
      RECT 5.545 4.165 5.715 4.335 ;
      RECT 5.545 4.545 5.715 4.715 ;
      RECT 5.545 8.605 5.715 8.775 ;
      RECT 5.525 2.765 5.695 2.935 ;
      RECT 5.525 5.945 5.695 6.115 ;
      RECT 4.905 0.915 5.075 1.085 ;
      RECT 4.905 2.395 5.075 2.565 ;
      RECT 4.905 6.315 5.075 6.485 ;
      RECT 4.905 7.795 5.075 7.965 ;
      RECT 4.555 0.105 4.725 0.275 ;
      RECT 4.555 4.165 4.725 4.335 ;
      RECT 4.555 4.545 4.725 4.715 ;
      RECT 4.555 8.605 4.725 8.775 ;
      RECT 4.535 2.765 4.705 2.935 ;
      RECT 4.535 5.945 4.705 6.115 ;
      RECT 3.85 0.105 4.02 0.275 ;
      RECT 3.85 4.165 4.02 4.335 ;
      RECT 3.85 4.545 4.02 4.715 ;
      RECT 3.85 8.605 4.02 8.775 ;
      RECT 3.54 2.025 3.71 2.195 ;
      RECT 3.54 6.685 3.71 6.855 ;
      RECT 3.17 0.105 3.34 0.275 ;
      RECT 3.17 8.605 3.34 8.775 ;
      RECT 3.11 0.915 3.28 1.085 ;
      RECT 3.11 1.655 3.28 1.825 ;
      RECT 3.11 7.055 3.28 7.225 ;
      RECT 3.11 7.795 3.28 7.965 ;
      RECT 2.735 2.395 2.905 2.565 ;
      RECT 2.735 6.315 2.905 6.485 ;
      RECT 2.49 0.105 2.66 0.275 ;
      RECT 2.49 8.605 2.66 8.775 ;
      RECT 1.81 0.105 1.98 0.275 ;
      RECT 1.81 8.605 1.98 8.775 ;
      RECT 1.74 2.765 1.91 2.935 ;
      RECT 1.74 5.945 1.91 6.115 ;
      RECT 0.35 1.415 0.52 1.585 ;
      RECT 0.35 4.135 0.52 4.305 ;
      RECT -0.11 1.415 0.06 1.585 ;
      RECT -0.11 4.135 0.06 4.305 ;
      RECT -0.325 2.775 -0.155 2.945 ;
      RECT -0.565 1.935 -0.395 2.105 ;
      RECT -0.565 3.615 -0.395 3.785 ;
      RECT -0.57 1.415 -0.4 1.585 ;
      RECT -0.57 4.135 -0.4 4.305 ;
      RECT -0.805 2.495 -0.635 2.665 ;
      RECT -0.805 3.055 -0.635 3.225 ;
      RECT -1.03 1.415 -0.86 1.585 ;
      RECT -1.03 4.135 -0.86 4.305 ;
      RECT -1.285 2.775 -1.115 2.945 ;
      RECT -1.49 1.415 -1.32 1.585 ;
      RECT -1.49 4.135 -1.32 4.305 ;
      RECT -1.525 1.935 -1.355 2.105 ;
      RECT -1.765 2.495 -1.595 2.665 ;
      RECT -1.95 1.415 -1.78 1.585 ;
      RECT -1.95 4.135 -1.78 4.305 ;
      RECT -1.975 3.335 -1.805 3.505 ;
      RECT -2.245 2.775 -2.075 2.945 ;
      RECT -2.41 1.415 -2.24 1.585 ;
      RECT -2.41 4.135 -2.24 4.305 ;
      RECT -2.515 3.615 -2.345 3.785 ;
      RECT -2.725 2.195 -2.555 2.365 ;
      RECT -2.87 1.415 -2.7 1.585 ;
      RECT -2.87 4.135 -2.7 4.305 ;
      RECT -3.205 2.775 -3.035 2.945 ;
      RECT -3.33 1.415 -3.16 1.585 ;
      RECT -3.33 4.135 -3.16 4.305 ;
      RECT -3.445 1.935 -3.275 2.105 ;
      RECT -3.685 2.495 -3.515 2.665 ;
      RECT -3.685 3.055 -3.515 3.225 ;
      RECT -3.79 1.415 -3.62 1.585 ;
      RECT -3.79 4.135 -3.62 4.305 ;
      RECT -4.165 2.495 -3.995 2.665 ;
      RECT -4.25 1.415 -4.08 1.585 ;
      RECT -4.25 4.135 -4.08 4.305 ;
      RECT -4.405 3.615 -4.235 3.785 ;
      RECT -4.445 1.935 -4.275 2.105 ;
      RECT -4.645 2.775 -4.475 2.945 ;
      RECT -4.71 1.415 -4.54 1.585 ;
      RECT -4.71 4.135 -4.54 4.305 ;
      RECT -4.885 3.615 -4.715 3.785 ;
      RECT -5.125 3.055 -4.955 3.225 ;
      RECT -5.17 1.415 -5 1.585 ;
      RECT -5.17 4.135 -5 4.305 ;
      RECT -5.605 2.495 -5.435 2.665 ;
      RECT -5.63 1.415 -5.46 1.585 ;
      RECT -5.63 4.135 -5.46 4.305 ;
      RECT -5.845 1.935 -5.675 2.105 ;
      RECT -5.845 3.615 -5.675 3.785 ;
      RECT -6.09 1.415 -5.92 1.585 ;
      RECT -6.09 4.135 -5.92 4.305 ;
      RECT -6.325 1.935 -6.155 2.105 ;
      RECT -6.325 3.055 -6.155 3.225 ;
      RECT -6.55 1.415 -6.38 1.585 ;
      RECT -6.55 4.135 -6.38 4.305 ;
      RECT -6.565 2.495 -6.395 2.665 ;
      RECT -6.805 3.335 -6.635 3.505 ;
      RECT -7.01 1.415 -6.84 1.585 ;
      RECT -7.01 4.135 -6.84 4.305 ;
      RECT -7.045 2.775 -6.875 2.945 ;
      RECT -7.47 1.415 -7.3 1.585 ;
      RECT -7.47 4.135 -7.3 4.305 ;
      RECT -7.525 2.775 -7.355 2.945 ;
      RECT -7.735 1.935 -7.565 2.105 ;
      RECT -7.735 3.335 -7.565 3.505 ;
      RECT -7.93 1.415 -7.76 1.585 ;
      RECT -7.93 4.135 -7.76 4.305 ;
    LAYER li ;
      RECT -0.105 0 0.065 2.085 ;
      RECT -1.045 0 -0.875 2.085 ;
      RECT -2.005 0 -1.835 2.085 ;
      RECT -3.925 0 -3.755 2.085 ;
      RECT -4.885 0 -4.715 2.085 ;
      RECT -6.805 0 -6.635 2.085 ;
      RECT -3.05 0 -2.855 1.595 ;
      RECT -6.805 0 -6.53 1.595 ;
      RECT -8.075 0 0.665 1.585 ;
      RECT 5.465 0 5.635 0.935 ;
      RECT 4.475 0 4.645 0.935 ;
      RECT 1.73 0 1.9 0.935 ;
      RECT -8.825 0 6.435 0.305 ;
      RECT 5.465 3.405 5.635 5.475 ;
      RECT 4.475 3.405 4.645 5.475 ;
      RECT 1.73 3.405 1.9 5.475 ;
      RECT -8.825 4.14 6.435 4.745 ;
      RECT -8.075 4.135 6.435 4.745 ;
      RECT -1.045 3.635 -0.875 4.745 ;
      RECT -2.965 3.635 -2.795 4.745 ;
      RECT -3.905 3.635 -3.735 4.745 ;
      RECT -5.365 3.635 -5.195 4.745 ;
      RECT -7.285 3.635 -7.115 4.745 ;
      RECT -8.825 8.575 6.435 8.88 ;
      RECT 5.465 7.945 5.635 8.88 ;
      RECT 4.475 7.945 4.645 8.88 ;
      RECT 1.73 7.945 1.9 8.88 ;
      RECT 5.525 1.74 5.695 2.935 ;
      RECT 5.525 1.74 5.99 1.91 ;
      RECT 5.525 6.97 5.99 7.14 ;
      RECT 5.525 5.945 5.695 7.14 ;
      RECT 4.535 1.74 4.705 2.935 ;
      RECT 4.535 1.74 5 1.91 ;
      RECT 4.535 6.97 5 7.14 ;
      RECT 4.535 5.945 4.705 7.14 ;
      RECT 2.68 2.635 2.85 3.865 ;
      RECT 2.735 0.855 2.905 2.805 ;
      RECT 2.68 0.575 2.85 1.025 ;
      RECT 2.68 7.855 2.85 8.305 ;
      RECT 2.735 6.075 2.905 8.025 ;
      RECT 2.68 5.015 2.85 6.245 ;
      RECT 2.16 0.575 2.33 3.865 ;
      RECT 2.16 2.075 2.565 2.405 ;
      RECT 2.16 1.235 2.565 1.565 ;
      RECT 2.16 5.015 2.33 8.305 ;
      RECT 2.16 7.315 2.565 7.645 ;
      RECT 2.16 6.475 2.565 6.805 ;
      RECT -0.565 3.615 -0.05 3.785 ;
      RECT -0.22 3.225 -0.05 3.785 ;
      RECT -0.115 3.145 0.055 3.475 ;
      RECT -0.325 2.535 -0.05 2.945 ;
      RECT -0.445 2.535 -0.05 2.745 ;
      RECT -1.975 3.145 -1.805 3.505 ;
      RECT -1.975 3.225 -0.635 3.395 ;
      RECT -0.805 3.055 -0.635 3.395 ;
      RECT -2.245 2.575 -2.075 2.945 ;
      RECT -2.725 2.575 -2.075 2.845 ;
      RECT -2.805 2.575 -1.995 2.745 ;
      RECT -3.445 1.815 -3.275 2.105 ;
      RECT -3.445 1.815 -2.205 1.985 ;
      RECT -2.725 2.155 -2.555 2.365 ;
      RECT -3.085 2.155 -2.555 2.325 ;
      RECT -3.685 3.225 -3.195 3.395 ;
      RECT -3.685 3.055 -3.515 3.395 ;
      RECT -4.405 3.225 -4.235 3.785 ;
      RECT -4.515 3.225 -4.185 3.395 ;
      RECT -4.445 1.835 -4.275 2.105 ;
      RECT -4.405 1.755 -4.235 2.085 ;
      RECT -4.54 1.835 -4.235 2.055 ;
      RECT -5.965 3.225 -5.675 3.785 ;
      RECT -5.845 3.145 -5.675 3.785 ;
      RECT -6.205 2.575 -5.835 2.745 ;
      RECT -6.205 1.935 -6.035 2.745 ;
      RECT -6.325 1.935 -6.035 2.105 ;
      RECT 5.895 0.575 6.065 1.085 ;
      RECT 5.895 2.395 6.065 3.865 ;
      RECT 5.895 5.015 6.065 6.485 ;
      RECT 5.895 7.795 6.065 8.305 ;
      RECT 4.905 0.575 5.075 1.085 ;
      RECT 4.905 2.395 5.075 3.865 ;
      RECT 4.905 5.015 5.075 6.485 ;
      RECT 4.905 7.795 5.075 8.305 ;
      RECT 3.54 0.575 3.71 3.865 ;
      RECT 3.54 5.015 3.71 8.305 ;
      RECT 3.11 0.575 3.28 1.085 ;
      RECT 3.11 1.655 3.28 3.865 ;
      RECT 3.11 5.015 3.28 7.225 ;
      RECT 3.11 7.795 3.28 8.305 ;
      RECT 1.74 1.66 1.91 2.935 ;
      RECT 1.74 5.945 1.91 7.22 ;
      RECT -0.565 1.755 -0.395 2.105 ;
      RECT -0.805 2.495 -0.635 2.825 ;
      RECT -1.285 2.495 -1.115 2.945 ;
      RECT -1.525 1.755 -1.355 2.105 ;
      RECT -1.765 2.495 -1.595 2.825 ;
      RECT -2.515 3.485 -2.345 3.815 ;
      RECT -3.205 2.495 -3.035 2.945 ;
      RECT -3.685 2.495 -3.515 2.825 ;
      RECT -4.165 2.495 -3.995 2.825 ;
      RECT -4.645 2.495 -4.475 2.945 ;
      RECT -4.885 3.485 -4.715 3.815 ;
      RECT -5.125 2.495 -4.955 3.225 ;
      RECT -5.605 2.495 -5.435 2.825 ;
      RECT -5.845 1.755 -5.675 2.105 ;
      RECT -6.325 3.055 -6.155 3.475 ;
      RECT -6.565 2.495 -6.395 2.825 ;
      RECT -6.805 3.145 -6.635 3.505 ;
      RECT -7.045 2.495 -6.875 2.945 ;
      RECT -7.525 2.495 -7.355 2.945 ;
      RECT -7.735 1.755 -7.565 2.105 ;
      RECT -7.735 3.145 -7.565 3.505 ;
  END
END sky130_osu_single_mpr2xa_8

MACRO sky130_osu_single_mpr2ya_8
  CLASS CORE ;
  ORIGIN 8.825 0 ;
  FOREIGN sky130_osu_single_mpr2ya_8 -8.825 0 ;
  SIZE 15.26 BY 8.88 ;
  SYMMETRY X Y ;
  SITE b0r2 ;
  OBS
    LAYER met3 ;
      RECT -4.965 1.855 -4.635 2.585 ;
      RECT -4.935 1.04 -4.625 1.985 ;
      RECT -4.96 1.04 -4.585 1.41 ;
      RECT -0.525 2.015 -0.195 2.745 ;
      RECT -1.725 2.88 -1.395 3.61 ;
      RECT -2.565 1.855 -1.835 2.185 ;
      RECT -4.005 1.855 -3.275 2.185 ;
      RECT -3.645 2.76 -3.315 3.49 ;
      RECT -6.165 2.015 -5.835 2.745 ;
      RECT -6.885 2.015 -6.555 2.745 ;
    LAYER via2 ;
      RECT -0.46 2.48 -0.26 2.68 ;
      RECT -1.66 3.04 -1.46 3.24 ;
      RECT -2.5 1.92 -2.3 2.12 ;
      RECT -3.58 2.825 -3.38 3.025 ;
      RECT -3.94 1.92 -3.74 2.12 ;
      RECT -4.87 1.125 -4.67 1.325 ;
      RECT -4.9 1.92 -4.7 2.12 ;
      RECT -6.1 2.48 -5.9 2.68 ;
      RECT -6.82 2.48 -6.62 2.68 ;
    LAYER met2 ;
      RECT 2.705 6.28 3.025 6.605 ;
      RECT 2.735 5.695 2.905 6.605 ;
      RECT 2.735 5.695 2.91 6.045 ;
      RECT 2.735 5.695 3.71 5.87 ;
      RECT 3.535 1.965 3.71 5.87 ;
      RECT -6.14 2.44 -5.86 2.72 ;
      RECT -6.14 2.44 -5.84 2.615 ;
      RECT -6.05 2.33 -5.79 2.59 ;
      RECT -6.085 2.425 -5.79 2.59 ;
      RECT -5.95 0.73 -5.795 2.59 ;
      RECT 3.48 1.965 3.83 2.315 ;
      RECT 1.07 2.025 3.83 2.195 ;
      RECT 1.07 0.73 1.24 2.195 ;
      RECT -5.95 0.73 1.24 0.9 ;
      RECT 3.505 6.655 3.83 6.98 ;
      RECT 2.39 6.745 3.83 6.915 ;
      RECT 2.39 2.395 2.55 6.915 ;
      RECT 2.705 2.365 3.025 2.685 ;
      RECT 2.39 2.395 3.025 2.565 ;
      RECT 1.655 5.86 1.995 6.21 ;
      RECT 1.735 2.705 1.91 6.21 ;
      RECT 1.66 2.705 2 3.055 ;
      RECT 1.1 2.705 1.44 3.055 ;
      RECT 0.4 2.77 1.44 2.97 ;
      RECT 0.4 2.765 0.71 2.97 ;
      RECT 0.4 1.04 0.605 2.97 ;
      RECT 1.19 2.7 1.36 3.055 ;
      RECT -4.96 1.04 -4.585 1.41 ;
      RECT -4.96 1.04 0.605 1.245 ;
      RECT -0.5 2.44 -0.22 2.72 ;
      RECT -0.505 2.44 -0.22 2.673 ;
      RECT -0.525 2.44 -0.22 2.65 ;
      RECT -0.535 2.44 -0.22 2.63 ;
      RECT -0.545 2.44 -0.22 2.615 ;
      RECT -0.57 2.44 -0.22 2.588 ;
      RECT -0.58 2.44 -0.22 2.563 ;
      RECT -0.625 2.295 -0.345 2.555 ;
      RECT -0.625 2.39 -0.245 2.555 ;
      RECT -0.625 2.335 -0.3 2.555 ;
      RECT -0.625 2.327 -0.305 2.555 ;
      RECT -0.625 2.317 -0.31 2.555 ;
      RECT -0.625 2.305 -0.315 2.555 ;
      RECT -1.7 3 -1.42 3.28 ;
      RECT -1.7 3 -1.385 3.26 ;
      RECT -1.665 2.42 -1.615 2.68 ;
      RECT -1.875 2.42 -1.87 2.68 ;
      RECT -2.68 1.975 -2.65 2.235 ;
      RECT -2.91 1.975 -2.835 2.235 ;
      RECT -1.69 2.37 -1.665 2.68 ;
      RECT -1.695 2.327 -1.69 2.68 ;
      RECT -1.7 2.31 -1.695 2.68 ;
      RECT -1.705 2.297 -1.7 2.68 ;
      RECT -1.78 2.18 -1.705 2.68 ;
      RECT -1.825 1.997 -1.78 2.68 ;
      RECT -1.83 1.925 -1.825 2.68 ;
      RECT -1.845 1.9 -1.83 2.68 ;
      RECT -1.87 1.862 -1.845 2.68 ;
      RECT -1.88 1.842 -1.87 2.402 ;
      RECT -1.895 1.834 -1.88 2.357 ;
      RECT -1.9 1.826 -1.895 2.328 ;
      RECT -1.905 1.823 -1.9 2.308 ;
      RECT -1.91 1.82 -1.905 2.288 ;
      RECT -1.915 1.817 -1.91 2.268 ;
      RECT -1.945 1.806 -1.915 2.205 ;
      RECT -1.965 1.791 -1.945 2.12 ;
      RECT -1.97 1.783 -1.965 2.083 ;
      RECT -1.98 1.777 -1.97 2.05 ;
      RECT -1.995 1.769 -1.98 2.01 ;
      RECT -2 1.762 -1.995 1.97 ;
      RECT -2.005 1.759 -2 1.948 ;
      RECT -2.01 1.756 -2.005 1.935 ;
      RECT -2.015 1.755 -2.01 1.925 ;
      RECT -2.03 1.749 -2.015 1.915 ;
      RECT -2.055 1.736 -2.03 1.9 ;
      RECT -2.105 1.711 -2.055 1.871 ;
      RECT -2.12 1.69 -2.105 1.846 ;
      RECT -2.13 1.683 -2.12 1.835 ;
      RECT -2.185 1.664 -2.13 1.808 ;
      RECT -2.21 1.642 -2.185 1.781 ;
      RECT -2.215 1.635 -2.21 1.776 ;
      RECT -2.23 1.635 -2.215 1.774 ;
      RECT -2.255 1.627 -2.23 1.77 ;
      RECT -2.27 1.625 -2.255 1.766 ;
      RECT -2.3 1.625 -2.27 1.763 ;
      RECT -2.31 1.625 -2.3 1.758 ;
      RECT -2.355 1.625 -2.31 1.756 ;
      RECT -2.384 1.625 -2.355 1.757 ;
      RECT -2.47 1.625 -2.384 1.759 ;
      RECT -2.484 1.626 -2.47 1.761 ;
      RECT -2.57 1.627 -2.484 1.763 ;
      RECT -2.585 1.628 -2.57 1.773 ;
      RECT -2.59 1.629 -2.585 1.782 ;
      RECT -2.61 1.632 -2.59 1.792 ;
      RECT -2.625 1.64 -2.61 1.807 ;
      RECT -2.645 1.658 -2.625 1.822 ;
      RECT -2.655 1.67 -2.645 1.845 ;
      RECT -2.665 1.679 -2.655 1.875 ;
      RECT -2.68 1.691 -2.665 1.92 ;
      RECT -2.735 1.724 -2.68 2.235 ;
      RECT -2.74 1.752 -2.735 2.235 ;
      RECT -2.76 1.767 -2.74 2.235 ;
      RECT -2.795 1.827 -2.76 2.235 ;
      RECT -2.797 1.877 -2.795 2.235 ;
      RECT -2.8 1.885 -2.797 2.235 ;
      RECT -2.81 1.9 -2.8 2.235 ;
      RECT -2.815 1.912 -2.81 2.235 ;
      RECT -2.825 1.937 -2.815 2.235 ;
      RECT -2.835 1.965 -2.825 2.235 ;
      RECT -4.93 3.47 -4.88 3.73 ;
      RECT -2.02 3.02 -1.96 3.28 ;
      RECT -2.035 3.02 -2.02 3.29 ;
      RECT -2.054 3.02 -2.035 3.323 ;
      RECT -2.14 3.02 -2.054 3.448 ;
      RECT -2.22 3.02 -2.14 3.63 ;
      RECT -2.225 3.257 -2.22 3.715 ;
      RECT -2.25 3.327 -2.225 3.743 ;
      RECT -2.255 3.397 -2.25 3.77 ;
      RECT -2.275 3.469 -2.255 3.792 ;
      RECT -2.28 3.536 -2.275 3.815 ;
      RECT -2.29 3.565 -2.28 3.83 ;
      RECT -2.3 3.587 -2.29 3.847 ;
      RECT -2.305 3.597 -2.3 3.858 ;
      RECT -2.31 3.605 -2.305 3.866 ;
      RECT -2.32 3.613 -2.31 3.878 ;
      RECT -2.325 3.625 -2.32 3.888 ;
      RECT -2.33 3.633 -2.325 3.893 ;
      RECT -2.35 3.651 -2.33 3.903 ;
      RECT -2.355 3.668 -2.35 3.91 ;
      RECT -2.36 3.676 -2.355 3.911 ;
      RECT -2.365 3.687 -2.36 3.913 ;
      RECT -2.405 3.725 -2.365 3.923 ;
      RECT -2.41 3.76 -2.405 3.934 ;
      RECT -2.415 3.765 -2.41 3.937 ;
      RECT -2.44 3.775 -2.415 3.944 ;
      RECT -2.45 3.789 -2.44 3.953 ;
      RECT -2.47 3.801 -2.45 3.956 ;
      RECT -2.52 3.82 -2.47 3.96 ;
      RECT -2.565 3.835 -2.52 3.965 ;
      RECT -2.63 3.838 -2.565 3.971 ;
      RECT -2.645 3.836 -2.63 3.978 ;
      RECT -2.675 3.835 -2.645 3.978 ;
      RECT -2.714 3.834 -2.675 3.974 ;
      RECT -2.8 3.831 -2.714 3.97 ;
      RECT -2.817 3.829 -2.8 3.967 ;
      RECT -2.903 3.827 -2.817 3.964 ;
      RECT -2.989 3.824 -2.903 3.958 ;
      RECT -3.075 3.82 -2.989 3.953 ;
      RECT -3.153 3.817 -3.075 3.949 ;
      RECT -3.239 3.814 -3.153 3.947 ;
      RECT -3.325 3.811 -3.239 3.944 ;
      RECT -3.383 3.809 -3.325 3.941 ;
      RECT -3.469 3.806 -3.383 3.939 ;
      RECT -3.555 3.802 -3.469 3.937 ;
      RECT -3.641 3.799 -3.555 3.934 ;
      RECT -3.727 3.795 -3.641 3.932 ;
      RECT -3.813 3.791 -3.727 3.929 ;
      RECT -3.899 3.788 -3.813 3.927 ;
      RECT -3.985 3.784 -3.899 3.924 ;
      RECT -4.071 3.781 -3.985 3.922 ;
      RECT -4.157 3.777 -4.071 3.919 ;
      RECT -4.243 3.774 -4.157 3.917 ;
      RECT -4.329 3.77 -4.243 3.914 ;
      RECT -4.415 3.767 -4.329 3.912 ;
      RECT -4.425 3.765 -4.415 3.908 ;
      RECT -4.43 3.765 -4.425 3.906 ;
      RECT -4.47 3.76 -4.43 3.9 ;
      RECT -4.484 3.751 -4.47 3.893 ;
      RECT -4.57 3.721 -4.484 3.878 ;
      RECT -4.59 3.687 -4.57 3.863 ;
      RECT -4.66 3.656 -4.59 3.85 ;
      RECT -4.665 3.631 -4.66 3.839 ;
      RECT -4.67 3.625 -4.665 3.837 ;
      RECT -4.739 3.47 -4.67 3.825 ;
      RECT -4.825 3.47 -4.739 3.799 ;
      RECT -4.85 3.47 -4.825 3.778 ;
      RECT -4.855 3.47 -4.85 3.768 ;
      RECT -4.86 3.47 -4.855 3.76 ;
      RECT -4.88 3.47 -4.86 3.743 ;
      RECT -2.46 2.04 -2.2 2.3 ;
      RECT -2.475 2.04 -2.2 2.203 ;
      RECT -2.505 2.04 -2.2 2.178 ;
      RECT -2.54 1.88 -2.26 2.16 ;
      RECT -2.57 3.37 -2.51 3.63 ;
      RECT -3.545 2.06 -3.49 2.32 ;
      RECT -2.61 3.327 -2.57 3.63 ;
      RECT -2.639 3.248 -2.61 3.63 ;
      RECT -2.725 3.12 -2.639 3.63 ;
      RECT -2.745 3 -2.725 3.63 ;
      RECT -2.77 2.951 -2.745 3.63 ;
      RECT -2.775 2.916 -2.77 3.48 ;
      RECT -2.805 2.876 -2.775 3.418 ;
      RECT -2.83 2.813 -2.805 3.333 ;
      RECT -2.84 2.775 -2.83 3.27 ;
      RECT -2.855 2.75 -2.84 3.231 ;
      RECT -2.898 2.708 -2.855 3.137 ;
      RECT -2.9 2.681 -2.898 3.064 ;
      RECT -2.905 2.676 -2.9 3.055 ;
      RECT -2.91 2.669 -2.905 3.03 ;
      RECT -2.915 2.663 -2.91 3.015 ;
      RECT -2.92 2.657 -2.915 3.003 ;
      RECT -2.93 2.648 -2.92 2.985 ;
      RECT -2.935 2.639 -2.93 2.963 ;
      RECT -2.96 2.62 -2.935 2.913 ;
      RECT -2.965 2.601 -2.96 2.863 ;
      RECT -2.98 2.587 -2.965 2.823 ;
      RECT -2.985 2.573 -2.98 2.79 ;
      RECT -2.99 2.566 -2.985 2.783 ;
      RECT -3.005 2.553 -2.99 2.775 ;
      RECT -3.05 2.515 -3.005 2.748 ;
      RECT -3.08 2.468 -3.05 2.713 ;
      RECT -3.1 2.437 -3.08 2.69 ;
      RECT -3.18 2.37 -3.1 2.643 ;
      RECT -3.21 2.3 -3.18 2.59 ;
      RECT -3.215 2.277 -3.21 2.573 ;
      RECT -3.245 2.255 -3.215 2.558 ;
      RECT -3.275 2.214 -3.245 2.53 ;
      RECT -3.28 2.189 -3.275 2.515 ;
      RECT -3.285 2.183 -3.28 2.508 ;
      RECT -3.295 2.06 -3.285 2.5 ;
      RECT -3.305 2.06 -3.295 2.493 ;
      RECT -3.31 2.06 -3.305 2.485 ;
      RECT -3.33 2.06 -3.31 2.473 ;
      RECT -3.38 2.06 -3.33 2.443 ;
      RECT -3.435 2.06 -3.38 2.393 ;
      RECT -3.465 2.06 -3.435 2.353 ;
      RECT -3.49 2.06 -3.465 2.33 ;
      RECT -3.62 2.785 -3.34 3.065 ;
      RECT -3.655 2.7 -3.395 2.96 ;
      RECT -3.655 2.782 -3.385 2.96 ;
      RECT -5.455 2.155 -5.45 2.64 ;
      RECT -5.565 2.34 -5.56 2.64 ;
      RECT -5.655 2.38 -5.59 2.64 ;
      RECT -3.98 1.88 -3.89 2.51 ;
      RECT -4.015 1.93 -4.01 2.51 ;
      RECT -4.07 1.955 -4.06 2.51 ;
      RECT -4.115 1.955 -4.105 2.51 ;
      RECT -3.745 1.88 -3.7 2.16 ;
      RECT -4.895 1.61 -4.695 1.75 ;
      RECT -3.779 1.88 -3.745 2.172 ;
      RECT -3.865 1.88 -3.779 2.212 ;
      RECT -3.88 1.88 -3.865 2.253 ;
      RECT -3.885 1.88 -3.88 2.273 ;
      RECT -3.89 1.88 -3.885 2.293 ;
      RECT -4.01 1.922 -3.98 2.51 ;
      RECT -4.06 1.942 -4.015 2.51 ;
      RECT -4.075 1.957 -4.07 2.51 ;
      RECT -4.105 1.957 -4.075 2.51 ;
      RECT -4.15 1.942 -4.115 2.51 ;
      RECT -4.155 1.93 -4.15 2.29 ;
      RECT -4.16 1.927 -4.155 2.27 ;
      RECT -4.175 1.917 -4.16 2.223 ;
      RECT -4.18 1.91 -4.175 2.186 ;
      RECT -4.185 1.907 -4.18 2.169 ;
      RECT -4.2 1.897 -4.185 2.125 ;
      RECT -4.205 1.888 -4.2 2.085 ;
      RECT -4.21 1.884 -4.205 2.07 ;
      RECT -4.22 1.878 -4.21 2.053 ;
      RECT -4.26 1.859 -4.22 2.028 ;
      RECT -4.265 1.841 -4.26 2.008 ;
      RECT -4.275 1.835 -4.265 2.003 ;
      RECT -4.305 1.819 -4.275 1.99 ;
      RECT -4.32 1.801 -4.305 1.973 ;
      RECT -4.335 1.789 -4.32 1.96 ;
      RECT -4.34 1.781 -4.335 1.953 ;
      RECT -4.37 1.767 -4.34 1.94 ;
      RECT -4.375 1.752 -4.37 1.928 ;
      RECT -4.385 1.746 -4.375 1.92 ;
      RECT -4.405 1.734 -4.385 1.908 ;
      RECT -4.415 1.722 -4.405 1.895 ;
      RECT -4.445 1.706 -4.415 1.88 ;
      RECT -4.465 1.686 -4.445 1.863 ;
      RECT -4.47 1.676 -4.465 1.853 ;
      RECT -4.495 1.664 -4.47 1.84 ;
      RECT -4.5 1.652 -4.495 1.828 ;
      RECT -4.505 1.647 -4.5 1.824 ;
      RECT -4.52 1.64 -4.505 1.816 ;
      RECT -4.53 1.627 -4.52 1.806 ;
      RECT -4.535 1.625 -4.53 1.8 ;
      RECT -4.56 1.618 -4.535 1.789 ;
      RECT -4.565 1.611 -4.56 1.778 ;
      RECT -4.59 1.61 -4.565 1.765 ;
      RECT -4.609 1.61 -4.59 1.755 ;
      RECT -4.695 1.61 -4.609 1.752 ;
      RECT -4.925 1.61 -4.895 1.755 ;
      RECT -4.965 1.617 -4.925 1.768 ;
      RECT -4.99 1.627 -4.965 1.781 ;
      RECT -5.005 1.636 -4.99 1.791 ;
      RECT -5.035 1.641 -5.005 1.81 ;
      RECT -5.04 1.647 -5.035 1.828 ;
      RECT -5.06 1.657 -5.04 1.843 ;
      RECT -5.07 1.67 -5.06 1.863 ;
      RECT -5.085 1.682 -5.07 1.88 ;
      RECT -5.09 1.692 -5.085 1.89 ;
      RECT -5.095 1.697 -5.09 1.895 ;
      RECT -5.105 1.705 -5.095 1.908 ;
      RECT -5.155 1.737 -5.105 1.945 ;
      RECT -5.17 1.772 -5.155 1.986 ;
      RECT -5.175 1.782 -5.17 2.001 ;
      RECT -5.18 1.787 -5.175 2.008 ;
      RECT -5.205 1.803 -5.18 2.028 ;
      RECT -5.22 1.824 -5.205 2.053 ;
      RECT -5.245 1.845 -5.22 2.078 ;
      RECT -5.255 1.864 -5.245 2.101 ;
      RECT -5.28 1.882 -5.255 2.124 ;
      RECT -5.295 1.902 -5.28 2.148 ;
      RECT -5.3 1.912 -5.295 2.16 ;
      RECT -5.315 1.924 -5.3 2.18 ;
      RECT -5.325 1.939 -5.315 2.22 ;
      RECT -5.33 1.947 -5.325 2.248 ;
      RECT -5.34 1.957 -5.33 2.268 ;
      RECT -5.345 1.97 -5.34 2.293 ;
      RECT -5.35 1.983 -5.345 2.313 ;
      RECT -5.355 1.989 -5.35 2.335 ;
      RECT -5.365 1.998 -5.355 2.355 ;
      RECT -5.37 2.018 -5.365 2.378 ;
      RECT -5.375 2.024 -5.37 2.398 ;
      RECT -5.38 2.031 -5.375 2.42 ;
      RECT -5.385 2.042 -5.38 2.433 ;
      RECT -5.395 2.052 -5.385 2.458 ;
      RECT -5.415 2.077 -5.395 2.64 ;
      RECT -5.445 2.117 -5.415 2.64 ;
      RECT -5.45 2.147 -5.445 2.64 ;
      RECT -5.475 2.175 -5.455 2.64 ;
      RECT -5.505 2.22 -5.475 2.64 ;
      RECT -5.51 2.247 -5.505 2.64 ;
      RECT -5.53 2.265 -5.51 2.64 ;
      RECT -5.54 2.29 -5.53 2.64 ;
      RECT -5.545 2.302 -5.54 2.64 ;
      RECT -5.56 2.325 -5.545 2.64 ;
      RECT -5.58 2.352 -5.565 2.64 ;
      RECT -5.59 2.375 -5.58 2.64 ;
      RECT -3.8 3.26 -3.72 3.52 ;
      RECT -4.565 2.48 -4.495 2.74 ;
      RECT -3.834 3.227 -3.8 3.52 ;
      RECT -3.92 3.13 -3.834 3.52 ;
      RECT -3.94 3.042 -3.92 3.52 ;
      RECT -3.95 3.012 -3.94 3.52 ;
      RECT -3.96 2.992 -3.95 3.52 ;
      RECT -3.98 2.979 -3.96 3.52 ;
      RECT -3.995 2.969 -3.98 3.348 ;
      RECT -4 2.962 -3.995 3.303 ;
      RECT -4.01 2.956 -4 3.293 ;
      RECT -4.02 2.948 -4.01 3.275 ;
      RECT -4.025 2.942 -4.02 3.263 ;
      RECT -4.035 2.937 -4.025 3.25 ;
      RECT -4.055 2.927 -4.035 3.223 ;
      RECT -4.095 2.906 -4.055 3.175 ;
      RECT -4.11 2.887 -4.095 3.133 ;
      RECT -4.135 2.873 -4.11 3.103 ;
      RECT -4.145 2.861 -4.135 3.07 ;
      RECT -4.15 2.856 -4.145 3.06 ;
      RECT -4.18 2.842 -4.15 3.04 ;
      RECT -4.19 2.826 -4.18 3.013 ;
      RECT -4.195 2.821 -4.19 3.003 ;
      RECT -4.22 2.812 -4.195 2.983 ;
      RECT -4.23 2.8 -4.22 2.963 ;
      RECT -4.3 2.768 -4.23 2.938 ;
      RECT -4.305 2.737 -4.3 2.915 ;
      RECT -4.354 2.48 -4.305 2.898 ;
      RECT -4.44 2.48 -4.354 2.857 ;
      RECT -4.495 2.48 -4.44 2.785 ;
      RECT -4.405 3.265 -4.245 3.525 ;
      RECT -4.88 1.88 -4.83 2.565 ;
      RECT -5.09 2.305 -5.055 2.565 ;
      RECT -4.775 1.88 -4.77 2.34 ;
      RECT -4.685 1.88 -4.66 2.16 ;
      RECT -4.41 3.262 -4.405 3.525 ;
      RECT -4.445 3.25 -4.41 3.525 ;
      RECT -4.505 3.223 -4.445 3.525 ;
      RECT -4.51 3.206 -4.505 3.379 ;
      RECT -4.515 3.203 -4.51 3.366 ;
      RECT -4.535 3.196 -4.515 3.353 ;
      RECT -4.57 3.179 -4.535 3.335 ;
      RECT -4.61 3.158 -4.57 3.315 ;
      RECT -4.615 3.146 -4.61 3.303 ;
      RECT -4.655 3.132 -4.615 3.289 ;
      RECT -4.675 3.115 -4.655 3.271 ;
      RECT -4.685 3.107 -4.675 3.263 ;
      RECT -4.7 1.88 -4.685 2.178 ;
      RECT -4.715 3.097 -4.685 3.25 ;
      RECT -4.73 1.88 -4.7 2.223 ;
      RECT -4.725 3.087 -4.715 3.237 ;
      RECT -4.755 3.072 -4.725 3.224 ;
      RECT -4.77 1.88 -4.73 2.29 ;
      RECT -4.77 3.04 -4.755 3.21 ;
      RECT -4.775 3.012 -4.77 3.204 ;
      RECT -4.78 1.88 -4.775 2.345 ;
      RECT -4.79 2.982 -4.775 3.198 ;
      RECT -4.785 1.88 -4.78 2.358 ;
      RECT -4.795 1.88 -4.785 2.378 ;
      RECT -4.83 2.895 -4.79 3.183 ;
      RECT -4.83 1.88 -4.795 2.418 ;
      RECT -4.835 2.827 -4.83 3.171 ;
      RECT -4.85 2.782 -4.835 3.166 ;
      RECT -4.855 2.72 -4.85 3.161 ;
      RECT -4.88 2.627 -4.855 3.154 ;
      RECT -4.885 1.88 -4.88 3.146 ;
      RECT -4.9 1.88 -4.885 3.133 ;
      RECT -4.92 1.88 -4.9 3.09 ;
      RECT -4.93 1.88 -4.92 3.04 ;
      RECT -4.935 1.88 -4.93 3.013 ;
      RECT -4.94 1.88 -4.935 2.991 ;
      RECT -4.945 2.106 -4.94 2.974 ;
      RECT -4.95 2.128 -4.945 2.952 ;
      RECT -4.955 2.17 -4.95 2.935 ;
      RECT -4.985 2.22 -4.955 2.879 ;
      RECT -4.99 2.247 -4.985 2.821 ;
      RECT -5.005 2.265 -4.99 2.785 ;
      RECT -5.01 2.283 -5.005 2.749 ;
      RECT -5.016 2.29 -5.01 2.73 ;
      RECT -5.02 2.297 -5.016 2.713 ;
      RECT -5.025 2.302 -5.02 2.682 ;
      RECT -5.035 2.305 -5.025 2.657 ;
      RECT -5.045 2.305 -5.035 2.623 ;
      RECT -5.05 2.305 -5.045 2.6 ;
      RECT -5.055 2.305 -5.05 2.58 ;
      RECT -6.435 3.47 -6.175 3.73 ;
      RECT -6.415 3.397 -6.235 3.73 ;
      RECT -6.415 3.14 -6.24 3.73 ;
      RECT -6.415 2.932 -6.25 3.73 ;
      RECT -6.41 2.85 -6.25 3.73 ;
      RECT -6.41 2.615 -6.26 3.73 ;
      RECT -6.41 2.462 -6.265 3.73 ;
      RECT -6.405 2.447 -6.265 3.73 ;
      RECT -6.355 2.162 -6.265 3.73 ;
      RECT -6.4 2.397 -6.265 3.73 ;
      RECT -6.37 2.215 -6.265 3.73 ;
      RECT -6.385 2.327 -6.265 3.73 ;
      RECT -6.38 2.285 -6.265 3.73 ;
      RECT -6.385 2.327 -6.25 2.39 ;
      RECT -6.35 1.915 -6.245 2.335 ;
      RECT -6.35 1.915 -6.23 2.318 ;
      RECT -6.35 1.915 -6.195 2.28 ;
      RECT -6.355 2.162 -6.145 2.213 ;
      RECT -6.35 1.915 -6.09 2.175 ;
      RECT -7.09 2.62 -6.83 2.88 ;
      RECT -7.09 2.62 -6.82 2.838 ;
      RECT -7.09 2.62 -6.734 2.809 ;
      RECT -7.09 2.62 -6.665 2.761 ;
      RECT -7.09 2.62 -6.63 2.73 ;
      RECT -6.86 2.44 -6.58 2.72 ;
      RECT -7.025 2.605 -6.58 2.72 ;
      RECT -6.935 2.482 -6.83 2.88 ;
      RECT -7.005 2.545 -6.58 2.72 ;
    LAYER via1 ;
      RECT 3.595 6.74 3.745 6.89 ;
      RECT 3.58 2.065 3.73 2.215 ;
      RECT 2.79 2.45 2.94 2.6 ;
      RECT 2.79 6.37 2.94 6.52 ;
      RECT 1.76 2.805 1.91 2.955 ;
      RECT 1.755 5.96 1.905 6.11 ;
      RECT 1.2 2.805 1.35 2.955 ;
      RECT -0.57 2.35 -0.42 2.5 ;
      RECT -1.59 3.055 -1.44 3.205 ;
      RECT -1.82 2.475 -1.67 2.625 ;
      RECT -2.165 3.075 -2.015 3.225 ;
      RECT -2.405 2.095 -2.255 2.245 ;
      RECT -2.715 3.425 -2.565 3.575 ;
      RECT -2.855 2.03 -2.705 2.18 ;
      RECT -3.49 2.115 -3.34 2.265 ;
      RECT -3.6 2.755 -3.45 2.905 ;
      RECT -3.925 3.315 -3.775 3.465 ;
      RECT -4.095 2.305 -3.945 2.455 ;
      RECT -4.45 3.32 -4.3 3.47 ;
      RECT -4.51 2.535 -4.36 2.685 ;
      RECT -4.875 3.525 -4.725 3.675 ;
      RECT -5.035 2.36 -4.885 2.51 ;
      RECT -5.6 2.435 -5.45 2.585 ;
      RECT -5.995 2.385 -5.845 2.535 ;
      RECT -6.295 1.97 -6.145 2.12 ;
      RECT -6.38 3.525 -6.23 3.675 ;
      RECT -7.035 2.675 -6.885 2.825 ;
    LAYER met1 ;
      RECT -8.075 0 0.665 1.74 ;
      RECT -8.825 0 6.435 0.305 ;
      RECT -8.825 4.14 6.435 4.745 ;
      RECT -8.075 4.135 6.435 4.745 ;
      RECT -8.075 3.98 0.665 4.745 ;
      RECT 5.835 2.365 6.125 2.595 ;
      RECT 5.895 0.885 6.065 2.595 ;
      RECT 5.835 0.885 6.125 1.115 ;
      RECT 5.835 7.765 6.125 7.995 ;
      RECT 5.895 6.285 6.065 7.995 ;
      RECT 5.835 6.285 6.125 6.515 ;
      RECT 5.425 2.735 5.755 2.965 ;
      RECT 5.425 2.765 5.925 2.935 ;
      RECT 5.425 2.395 5.615 2.965 ;
      RECT 4.845 2.365 5.135 2.595 ;
      RECT 4.845 2.395 5.615 2.565 ;
      RECT 4.905 0.885 5.075 2.595 ;
      RECT 4.845 0.885 5.135 1.115 ;
      RECT 4.845 7.765 5.135 7.995 ;
      RECT 4.905 6.285 5.075 7.995 ;
      RECT 4.845 6.285 5.135 6.515 ;
      RECT 4.845 6.325 5.695 6.485 ;
      RECT 5.525 5.915 5.695 6.485 ;
      RECT 4.845 6.32 5.235 6.485 ;
      RECT 5.465 5.915 5.755 6.145 ;
      RECT 5.465 5.945 5.925 6.115 ;
      RECT 4.475 2.735 4.765 2.965 ;
      RECT 4.475 2.765 4.935 2.935 ;
      RECT 4.535 1.655 4.7 2.965 ;
      RECT 3.05 1.625 3.34 1.855 ;
      RECT 3.05 1.655 4.7 1.825 ;
      RECT 3.11 0.885 3.28 1.855 ;
      RECT 3.05 0.885 3.34 1.115 ;
      RECT 3.05 7.765 3.34 7.995 ;
      RECT 3.11 7.025 3.28 7.995 ;
      RECT 3.11 7.12 4.7 7.29 ;
      RECT 4.53 5.915 4.7 7.29 ;
      RECT 3.05 7.025 3.34 7.255 ;
      RECT 4.475 5.915 4.765 6.145 ;
      RECT 4.475 5.945 4.935 6.115 ;
      RECT 3.48 1.965 3.83 2.315 ;
      RECT 3.31 2.025 3.83 2.195 ;
      RECT 3.505 6.655 3.83 6.98 ;
      RECT 3.48 6.655 3.83 6.885 ;
      RECT 3.31 6.685 3.83 6.855 ;
      RECT 1.1 2.705 1.44 3.055 ;
      RECT 1.19 2.395 1.36 3.055 ;
      RECT 2.705 2.365 3.025 2.685 ;
      RECT 2.675 2.365 3.025 2.595 ;
      RECT 1.19 2.395 3.025 2.565 ;
      RECT 2.705 6.28 3.025 6.605 ;
      RECT 2.675 6.285 3.025 6.515 ;
      RECT 2.505 6.315 3.025 6.485 ;
      RECT 1.66 2.705 2 3.055 ;
      RECT 1.66 2.765 2.14 2.935 ;
      RECT 1.655 5.86 1.995 6.21 ;
      RECT 1.655 5.945 2.14 6.115 ;
      RECT -1.605 2.985 -1.455 3.26 ;
      RECT -1.065 2.065 -1.06 2.285 ;
      RECT 0.085 2.265 0.1 2.463 ;
      RECT 0.05 2.257 0.085 2.47 ;
      RECT 0.02 2.25 0.05 2.47 ;
      RECT -0.035 2.215 0.02 2.47 ;
      RECT -0.1 2.152 -0.035 2.47 ;
      RECT -0.105 2.117 -0.1 2.468 ;
      RECT -0.11 2.112 -0.105 2.46 ;
      RECT -0.115 2.107 -0.11 2.446 ;
      RECT -0.12 2.104 -0.115 2.439 ;
      RECT -0.165 2.094 -0.12 2.39 ;
      RECT -0.185 2.081 -0.165 2.325 ;
      RECT -0.19 2.076 -0.185 2.298 ;
      RECT -0.195 2.075 -0.19 2.291 ;
      RECT -0.2 2.074 -0.195 2.284 ;
      RECT -0.285 2.059 -0.2 2.23 ;
      RECT -0.315 2.04 -0.285 2.18 ;
      RECT -0.395 2.023 -0.315 2.165 ;
      RECT -0.43 2.01 -0.395 2.15 ;
      RECT -0.438 2.01 -0.43 2.145 ;
      RECT -0.524 2.011 -0.438 2.145 ;
      RECT -0.61 2.013 -0.524 2.145 ;
      RECT -0.635 2.014 -0.61 2.149 ;
      RECT -0.71 2.02 -0.635 2.164 ;
      RECT -0.793 2.032 -0.71 2.188 ;
      RECT -0.879 2.045 -0.793 2.214 ;
      RECT -0.965 2.058 -0.879 2.24 ;
      RECT -1 2.067 -0.965 2.259 ;
      RECT -1.05 2.067 -1 2.272 ;
      RECT -1.06 2.065 -1.05 2.283 ;
      RECT -1.075 2.062 -1.065 2.285 ;
      RECT -1.09 2.054 -1.075 2.293 ;
      RECT -1.105 2.046 -1.09 2.313 ;
      RECT -1.11 2.041 -1.105 2.37 ;
      RECT -1.125 2.036 -1.11 2.443 ;
      RECT -1.13 2.031 -1.125 2.485 ;
      RECT -1.135 2.029 -1.13 2.513 ;
      RECT -1.14 2.027 -1.135 2.535 ;
      RECT -1.15 2.023 -1.14 2.578 ;
      RECT -1.155 2.02 -1.15 2.603 ;
      RECT -1.16 2.018 -1.155 2.623 ;
      RECT -1.165 2.016 -1.16 2.647 ;
      RECT -1.17 2.012 -1.165 2.67 ;
      RECT -1.175 2.008 -1.17 2.693 ;
      RECT -1.21 1.998 -1.175 2.8 ;
      RECT -1.215 1.988 -1.21 2.898 ;
      RECT -1.22 1.986 -1.215 2.925 ;
      RECT -1.225 1.985 -1.22 2.945 ;
      RECT -1.23 1.977 -1.225 2.965 ;
      RECT -1.235 1.972 -1.23 3 ;
      RECT -1.24 1.97 -1.235 3.018 ;
      RECT -1.245 1.97 -1.24 3.043 ;
      RECT -1.25 1.97 -1.245 3.065 ;
      RECT -1.285 1.97 -1.25 3.108 ;
      RECT -1.31 1.97 -1.285 3.137 ;
      RECT -1.32 1.97 -1.31 2.323 ;
      RECT -1.317 2.38 -1.31 3.147 ;
      RECT -1.32 2.437 -1.317 3.15 ;
      RECT -1.325 1.97 -1.32 2.295 ;
      RECT -1.325 2.487 -1.32 3.153 ;
      RECT -1.335 1.97 -1.325 2.285 ;
      RECT -1.33 2.54 -1.325 3.156 ;
      RECT -1.335 2.625 -1.33 3.16 ;
      RECT -1.345 1.97 -1.335 2.273 ;
      RECT -1.34 2.672 -1.335 3.164 ;
      RECT -1.345 2.747 -1.34 3.168 ;
      RECT -1.38 1.97 -1.345 2.248 ;
      RECT -1.355 2.83 -1.345 3.173 ;
      RECT -1.365 2.897 -1.355 3.18 ;
      RECT -1.37 2.925 -1.365 3.185 ;
      RECT -1.38 2.938 -1.37 3.191 ;
      RECT -1.425 1.97 -1.38 2.205 ;
      RECT -1.385 2.943 -1.38 3.198 ;
      RECT -1.425 2.96 -1.385 3.26 ;
      RECT -1.43 1.972 -1.425 2.178 ;
      RECT -1.455 2.98 -1.425 3.26 ;
      RECT -1.435 1.977 -1.43 2.15 ;
      RECT -1.645 2.989 -1.605 3.26 ;
      RECT -1.67 2.997 -1.645 3.23 ;
      RECT -1.715 3.005 -1.67 3.23 ;
      RECT -1.73 3.01 -1.715 3.225 ;
      RECT -1.74 3.01 -1.73 3.219 ;
      RECT -1.75 3.017 -1.74 3.216 ;
      RECT -1.755 3.055 -1.75 3.205 ;
      RECT -1.76 3.117 -1.755 3.183 ;
      RECT -0.49 2.992 -0.305 3.215 ;
      RECT -0.49 3.007 -0.3 3.211 ;
      RECT -0.5 2.28 -0.415 3.21 ;
      RECT -0.5 3.007 -0.295 3.204 ;
      RECT -0.505 3.015 -0.295 3.203 ;
      RECT -0.3 2.735 0.02 3.055 ;
      RECT -0.505 2.907 -0.335 2.998 ;
      RECT -0.51 2.907 -0.335 2.98 ;
      RECT -0.52 2.715 -0.385 2.955 ;
      RECT -0.525 2.715 -0.385 2.9 ;
      RECT -0.565 2.295 -0.395 2.8 ;
      RECT -0.58 2.295 -0.395 2.67 ;
      RECT -0.585 2.295 -0.395 2.623 ;
      RECT -0.59 2.295 -0.395 2.603 ;
      RECT -0.595 2.295 -0.395 2.578 ;
      RECT -0.625 2.295 -0.365 2.555 ;
      RECT -0.615 2.292 -0.405 2.555 ;
      RECT -0.49 2.287 -0.405 3.215 ;
      RECT -0.605 2.28 -0.415 2.555 ;
      RECT -0.61 2.285 -0.415 2.555 ;
      RECT -1.78 2.497 -1.595 2.71 ;
      RECT -1.78 2.505 -1.585 2.703 ;
      RECT -1.8 2.505 -1.585 2.7 ;
      RECT -1.805 2.505 -1.585 2.685 ;
      RECT -1.875 2.42 -1.615 2.68 ;
      RECT -1.875 2.565 -1.58 2.593 ;
      RECT -2.22 3.02 -1.96 3.28 ;
      RECT -2.195 2.965 -2 3.28 ;
      RECT -2.2 2.714 -2.02 3.008 ;
      RECT -2.2 2.72 -2.01 3.008 ;
      RECT -2.22 2.722 -2.01 2.953 ;
      RECT -2.225 2.732 -2.01 2.82 ;
      RECT -2.195 2.712 -2.02 3.28 ;
      RECT -2.109 2.71 -2.02 3.28 ;
      RECT -2.25 1.93 -2.215 2.3 ;
      RECT -2.46 2.04 -2.455 2.3 ;
      RECT -2.215 1.937 -2.2 2.3 ;
      RECT -2.325 1.93 -2.25 2.378 ;
      RECT -2.335 1.93 -2.325 2.463 ;
      RECT -2.36 1.93 -2.335 2.498 ;
      RECT -2.4 1.93 -2.36 2.566 ;
      RECT -2.41 1.937 -2.4 2.618 ;
      RECT -2.44 2.04 -2.41 2.659 ;
      RECT -2.445 2.04 -2.44 2.698 ;
      RECT -2.455 2.04 -2.445 2.718 ;
      RECT -2.46 2.335 -2.455 2.755 ;
      RECT -2.465 2.352 -2.46 2.775 ;
      RECT -2.48 2.415 -2.465 2.815 ;
      RECT -2.485 2.458 -2.48 2.85 ;
      RECT -2.49 2.466 -2.485 2.863 ;
      RECT -2.5 2.48 -2.49 2.885 ;
      RECT -2.525 2.515 -2.5 2.95 ;
      RECT -2.535 2.55 -2.525 3.013 ;
      RECT -2.555 2.58 -2.535 3.074 ;
      RECT -2.57 2.616 -2.555 3.141 ;
      RECT -2.58 2.644 -2.57 3.18 ;
      RECT -2.59 2.666 -2.58 3.2 ;
      RECT -2.595 2.676 -2.59 3.211 ;
      RECT -2.6 2.685 -2.595 3.214 ;
      RECT -2.61 2.703 -2.6 3.218 ;
      RECT -2.62 2.721 -2.61 3.219 ;
      RECT -2.645 2.76 -2.62 3.216 ;
      RECT -2.665 2.802 -2.645 3.213 ;
      RECT -2.68 2.84 -2.665 3.212 ;
      RECT -2.715 2.875 -2.68 3.209 ;
      RECT -2.72 2.897 -2.715 3.207 ;
      RECT -2.785 2.937 -2.72 3.204 ;
      RECT -2.79 2.977 -2.785 3.2 ;
      RECT -2.805 2.987 -2.79 3.191 ;
      RECT -2.815 3.107 -2.805 3.176 ;
      RECT -2.335 3.52 -2.325 3.78 ;
      RECT -2.335 3.523 -2.315 3.779 ;
      RECT -2.345 3.513 -2.335 3.778 ;
      RECT -2.355 3.528 -2.275 3.774 ;
      RECT -2.37 3.507 -2.355 3.772 ;
      RECT -2.395 3.532 -2.27 3.768 ;
      RECT -2.41 3.492 -2.395 3.763 ;
      RECT -2.41 3.534 -2.26 3.762 ;
      RECT -2.41 3.542 -2.245 3.755 ;
      RECT -2.47 3.479 -2.41 3.745 ;
      RECT -2.48 3.466 -2.47 3.727 ;
      RECT -2.505 3.456 -2.48 3.717 ;
      RECT -2.51 3.446 -2.505 3.709 ;
      RECT -2.575 3.542 -2.245 3.691 ;
      RECT -2.66 3.542 -2.245 3.653 ;
      RECT -2.77 3.37 -2.51 3.63 ;
      RECT -2.395 3.5 -2.37 3.768 ;
      RECT -2.355 3.51 -2.345 3.774 ;
      RECT -2.77 3.518 -2.33 3.63 ;
      RECT -3.555 3.275 -3.525 3.575 ;
      RECT -3.78 3.26 -3.775 3.535 ;
      RECT -3.98 3.26 -3.825 3.52 ;
      RECT -2.68 1.975 -2.65 2.235 ;
      RECT -2.69 1.975 -2.68 2.343 ;
      RECT -2.71 1.975 -2.69 2.353 ;
      RECT -2.725 1.975 -2.71 2.365 ;
      RECT -2.78 1.975 -2.725 2.415 ;
      RECT -2.795 1.975 -2.78 2.463 ;
      RECT -2.825 1.975 -2.795 2.498 ;
      RECT -2.88 1.975 -2.825 2.56 ;
      RECT -2.9 1.975 -2.88 2.628 ;
      RECT -2.905 1.975 -2.9 2.658 ;
      RECT -2.91 1.975 -2.905 2.67 ;
      RECT -2.915 2.092 -2.91 2.688 ;
      RECT -2.935 2.11 -2.915 2.713 ;
      RECT -2.955 2.137 -2.935 2.763 ;
      RECT -2.96 2.157 -2.955 2.794 ;
      RECT -2.965 2.165 -2.96 2.811 ;
      RECT -2.98 2.191 -2.965 2.84 ;
      RECT -2.995 2.233 -2.98 2.875 ;
      RECT -3 2.262 -2.995 2.898 ;
      RECT -3.005 2.277 -3 2.911 ;
      RECT -3.01 2.3 -3.005 2.922 ;
      RECT -3.02 2.32 -3.01 2.94 ;
      RECT -3.03 2.35 -3.02 2.963 ;
      RECT -3.035 2.372 -3.03 2.983 ;
      RECT -3.04 2.387 -3.035 2.998 ;
      RECT -3.055 2.417 -3.04 3.025 ;
      RECT -3.06 2.447 -3.055 3.051 ;
      RECT -3.065 2.465 -3.06 3.063 ;
      RECT -3.075 2.495 -3.065 3.082 ;
      RECT -3.085 2.52 -3.075 3.107 ;
      RECT -3.09 2.54 -3.085 3.126 ;
      RECT -3.095 2.557 -3.09 3.139 ;
      RECT -3.105 2.583 -3.095 3.158 ;
      RECT -3.115 2.621 -3.105 3.185 ;
      RECT -3.12 2.647 -3.115 3.205 ;
      RECT -3.125 2.657 -3.12 3.215 ;
      RECT -3.13 2.67 -3.125 3.23 ;
      RECT -3.135 2.685 -3.13 3.24 ;
      RECT -3.14 2.707 -3.135 3.255 ;
      RECT -3.145 2.725 -3.14 3.266 ;
      RECT -3.15 2.735 -3.145 3.277 ;
      RECT -3.155 2.743 -3.15 3.289 ;
      RECT -3.16 2.751 -3.155 3.3 ;
      RECT -3.165 2.777 -3.16 3.313 ;
      RECT -3.175 2.805 -3.165 3.326 ;
      RECT -3.18 2.835 -3.175 3.335 ;
      RECT -3.185 2.85 -3.18 3.342 ;
      RECT -3.2 2.875 -3.185 3.349 ;
      RECT -3.205 2.897 -3.2 3.355 ;
      RECT -3.21 2.922 -3.205 3.358 ;
      RECT -3.219 2.95 -3.21 3.362 ;
      RECT -3.225 2.967 -3.219 3.367 ;
      RECT -3.23 2.985 -3.225 3.371 ;
      RECT -3.235 2.997 -3.23 3.374 ;
      RECT -3.24 3.018 -3.235 3.378 ;
      RECT -3.245 3.036 -3.24 3.381 ;
      RECT -3.25 3.05 -3.245 3.384 ;
      RECT -3.255 3.067 -3.25 3.387 ;
      RECT -3.26 3.08 -3.255 3.39 ;
      RECT -3.285 3.117 -3.26 3.398 ;
      RECT -3.29 3.162 -3.285 3.407 ;
      RECT -3.295 3.19 -3.29 3.41 ;
      RECT -3.305 3.21 -3.295 3.414 ;
      RECT -3.31 3.23 -3.305 3.419 ;
      RECT -3.315 3.245 -3.31 3.422 ;
      RECT -3.335 3.255 -3.315 3.429 ;
      RECT -3.4 3.262 -3.335 3.455 ;
      RECT -3.435 3.265 -3.4 3.483 ;
      RECT -3.45 3.268 -3.435 3.498 ;
      RECT -3.46 3.269 -3.45 3.513 ;
      RECT -3.47 3.27 -3.46 3.53 ;
      RECT -3.475 3.27 -3.47 3.545 ;
      RECT -3.48 3.27 -3.475 3.553 ;
      RECT -3.495 3.271 -3.48 3.568 ;
      RECT -3.525 3.273 -3.495 3.575 ;
      RECT -3.635 3.28 -3.555 3.575 ;
      RECT -3.68 3.285 -3.635 3.575 ;
      RECT -3.69 3.286 -3.68 3.565 ;
      RECT -3.7 3.287 -3.69 3.558 ;
      RECT -3.72 3.289 -3.7 3.553 ;
      RECT -3.73 3.26 -3.72 3.548 ;
      RECT -3.775 3.26 -3.73 3.54 ;
      RECT -3.805 3.26 -3.78 3.53 ;
      RECT -3.825 3.26 -3.805 3.523 ;
      RECT -3.545 2.06 -3.285 2.32 ;
      RECT -3.665 2.075 -3.655 2.24 ;
      RECT -3.68 2.075 -3.675 2.235 ;
      RECT -6.315 1.915 -6.13 2.205 ;
      RECT -4.5 2.04 -4.485 2.195 ;
      RECT -6.35 1.915 -6.325 2.175 ;
      RECT -3.935 1.965 -3.93 2.107 ;
      RECT -4.02 1.96 -3.995 2.1 ;
      RECT -3.62 2.077 -3.545 2.27 ;
      RECT -3.635 2.075 -3.62 2.253 ;
      RECT -3.655 2.075 -3.635 2.245 ;
      RECT -3.675 2.075 -3.665 2.238 ;
      RECT -3.72 2.07 -3.68 2.228 ;
      RECT -3.76 2.045 -3.72 2.213 ;
      RECT -3.775 2.02 -3.76 2.203 ;
      RECT -3.78 2.014 -3.775 2.201 ;
      RECT -3.815 2.006 -3.78 2.184 ;
      RECT -3.82 1.999 -3.815 2.172 ;
      RECT -3.84 1.994 -3.82 2.16 ;
      RECT -3.85 1.988 -3.84 2.145 ;
      RECT -3.87 1.983 -3.85 2.13 ;
      RECT -3.88 1.978 -3.87 2.123 ;
      RECT -3.885 1.976 -3.88 2.118 ;
      RECT -3.89 1.975 -3.885 2.115 ;
      RECT -3.93 1.97 -3.89 2.111 ;
      RECT -3.95 1.964 -3.935 2.106 ;
      RECT -3.985 1.961 -3.95 2.103 ;
      RECT -3.995 1.96 -3.985 2.101 ;
      RECT -4.055 1.96 -4.02 2.098 ;
      RECT -4.1 1.96 -4.055 2.098 ;
      RECT -4.15 1.96 -4.1 2.101 ;
      RECT -4.165 1.962 -4.15 2.103 ;
      RECT -4.18 1.965 -4.165 2.104 ;
      RECT -4.19 1.97 -4.18 2.105 ;
      RECT -4.22 1.975 -4.19 2.11 ;
      RECT -4.23 1.981 -4.22 2.118 ;
      RECT -4.24 1.983 -4.23 2.122 ;
      RECT -4.25 1.987 -4.24 2.126 ;
      RECT -4.275 1.993 -4.25 2.134 ;
      RECT -4.285 1.998 -4.275 2.142 ;
      RECT -4.3 2.002 -4.285 2.146 ;
      RECT -4.335 2.008 -4.3 2.154 ;
      RECT -4.355 2.013 -4.335 2.164 ;
      RECT -4.385 2.02 -4.355 2.173 ;
      RECT -4.43 2.029 -4.385 2.187 ;
      RECT -4.435 2.034 -4.43 2.198 ;
      RECT -4.455 2.037 -4.435 2.199 ;
      RECT -4.485 2.04 -4.455 2.197 ;
      RECT -4.52 2.04 -4.5 2.193 ;
      RECT -4.59 2.04 -4.52 2.184 ;
      RECT -4.605 2.037 -4.59 2.176 ;
      RECT -4.645 2.03 -4.605 2.171 ;
      RECT -4.67 2.02 -4.645 2.164 ;
      RECT -4.675 2.014 -4.67 2.161 ;
      RECT -4.715 2.008 -4.675 2.158 ;
      RECT -4.73 2.001 -4.715 2.153 ;
      RECT -4.75 1.997 -4.73 2.148 ;
      RECT -4.765 1.992 -4.75 2.144 ;
      RECT -4.78 1.987 -4.765 2.142 ;
      RECT -4.795 1.983 -4.78 2.141 ;
      RECT -4.81 1.981 -4.795 2.137 ;
      RECT -4.82 1.979 -4.81 2.132 ;
      RECT -4.835 1.976 -4.82 2.128 ;
      RECT -4.845 1.974 -4.835 2.123 ;
      RECT -4.865 1.971 -4.845 2.119 ;
      RECT -4.91 1.97 -4.865 2.117 ;
      RECT -4.97 1.972 -4.91 2.118 ;
      RECT -4.99 1.974 -4.97 2.12 ;
      RECT -5.02 1.977 -4.99 2.121 ;
      RECT -5.07 1.982 -5.02 2.123 ;
      RECT -5.075 1.985 -5.07 2.125 ;
      RECT -5.085 1.987 -5.075 2.128 ;
      RECT -5.09 1.989 -5.085 2.131 ;
      RECT -5.14 1.992 -5.09 2.138 ;
      RECT -5.16 1.996 -5.14 2.15 ;
      RECT -5.17 1.999 -5.16 2.156 ;
      RECT -5.18 2 -5.17 2.159 ;
      RECT -5.219 2.003 -5.18 2.161 ;
      RECT -5.305 2.01 -5.219 2.164 ;
      RECT -5.379 2.02 -5.305 2.168 ;
      RECT -5.465 2.031 -5.379 2.173 ;
      RECT -5.48 2.038 -5.465 2.175 ;
      RECT -5.535 2.042 -5.48 2.176 ;
      RECT -5.549 2.045 -5.535 2.178 ;
      RECT -5.635 2.045 -5.549 2.18 ;
      RECT -5.675 2.042 -5.635 2.183 ;
      RECT -5.699 2.038 -5.675 2.185 ;
      RECT -5.785 2.028 -5.699 2.188 ;
      RECT -5.815 2.017 -5.785 2.189 ;
      RECT -5.834 2.013 -5.815 2.188 ;
      RECT -5.92 2.006 -5.834 2.185 ;
      RECT -5.98 1.995 -5.92 2.182 ;
      RECT -6 1.987 -5.98 2.18 ;
      RECT -6.035 1.982 -6 2.179 ;
      RECT -6.06 1.977 -6.035 2.178 ;
      RECT -6.09 1.972 -6.06 2.177 ;
      RECT -6.115 1.915 -6.09 2.176 ;
      RECT -6.13 1.915 -6.115 2.2 ;
      RECT -6.325 1.915 -6.315 2.2 ;
      RECT -4.55 2.935 -4.545 3.075 ;
      RECT -4.89 2.935 -4.855 3.073 ;
      RECT -5.315 2.92 -5.3 3.065 ;
      RECT -3.485 2.7 -3.395 2.96 ;
      RECT -3.655 2.565 -3.555 2.96 ;
      RECT -6.62 2.54 -6.54 2.75 ;
      RECT -3.53 2.677 -3.485 2.96 ;
      RECT -3.54 2.647 -3.53 2.96 ;
      RECT -3.555 2.57 -3.54 2.96 ;
      RECT -3.74 2.565 -3.655 2.925 ;
      RECT -3.745 2.567 -3.74 2.92 ;
      RECT -3.75 2.572 -3.745 2.92 ;
      RECT -3.785 2.672 -3.75 2.92 ;
      RECT -3.795 2.7 -3.785 2.92 ;
      RECT -3.805 2.715 -3.795 2.92 ;
      RECT -3.815 2.727 -3.805 2.92 ;
      RECT -3.82 2.737 -3.815 2.92 ;
      RECT -3.835 2.747 -3.82 2.922 ;
      RECT -3.84 2.762 -3.835 2.924 ;
      RECT -3.855 2.775 -3.84 2.926 ;
      RECT -3.86 2.79 -3.855 2.929 ;
      RECT -3.88 2.8 -3.86 2.933 ;
      RECT -3.895 2.81 -3.88 2.936 ;
      RECT -3.93 2.817 -3.895 2.941 ;
      RECT -3.974 2.824 -3.93 2.949 ;
      RECT -4.06 2.836 -3.974 2.962 ;
      RECT -4.085 2.847 -4.06 2.973 ;
      RECT -4.115 2.852 -4.085 2.978 ;
      RECT -4.15 2.857 -4.115 2.986 ;
      RECT -4.18 2.862 -4.15 2.993 ;
      RECT -4.205 2.867 -4.18 2.998 ;
      RECT -4.27 2.874 -4.205 3.007 ;
      RECT -4.34 2.887 -4.27 3.023 ;
      RECT -4.37 2.897 -4.34 3.035 ;
      RECT -4.395 2.902 -4.37 3.042 ;
      RECT -4.45 2.909 -4.395 3.05 ;
      RECT -4.455 2.916 -4.45 3.055 ;
      RECT -4.46 2.918 -4.455 3.056 ;
      RECT -4.475 2.92 -4.46 3.058 ;
      RECT -4.48 2.92 -4.475 3.061 ;
      RECT -4.545 2.927 -4.48 3.068 ;
      RECT -4.58 2.937 -4.55 3.078 ;
      RECT -4.597 2.94 -4.58 3.08 ;
      RECT -4.683 2.939 -4.597 3.079 ;
      RECT -4.769 2.937 -4.683 3.076 ;
      RECT -4.855 2.936 -4.769 3.074 ;
      RECT -4.956 2.934 -4.89 3.073 ;
      RECT -5.042 2.931 -4.956 3.071 ;
      RECT -5.128 2.927 -5.042 3.069 ;
      RECT -5.214 2.924 -5.128 3.068 ;
      RECT -5.3 2.921 -5.214 3.066 ;
      RECT -5.4 2.92 -5.315 3.063 ;
      RECT -5.45 2.918 -5.4 3.061 ;
      RECT -5.47 2.915 -5.45 3.059 ;
      RECT -5.49 2.913 -5.47 3.056 ;
      RECT -5.515 2.909 -5.49 3.053 ;
      RECT -5.56 2.903 -5.515 3.048 ;
      RECT -5.6 2.897 -5.56 3.04 ;
      RECT -5.625 2.892 -5.6 3.033 ;
      RECT -5.68 2.885 -5.625 3.025 ;
      RECT -5.704 2.878 -5.68 3.018 ;
      RECT -5.79 2.869 -5.704 3.008 ;
      RECT -5.82 2.861 -5.79 2.998 ;
      RECT -5.85 2.857 -5.82 2.993 ;
      RECT -5.855 2.854 -5.85 2.99 ;
      RECT -5.86 2.853 -5.855 2.99 ;
      RECT -5.935 2.846 -5.86 2.983 ;
      RECT -5.974 2.837 -5.935 2.972 ;
      RECT -6.06 2.827 -5.974 2.96 ;
      RECT -6.1 2.817 -6.06 2.948 ;
      RECT -6.139 2.812 -6.1 2.941 ;
      RECT -6.225 2.802 -6.139 2.93 ;
      RECT -6.265 2.79 -6.225 2.919 ;
      RECT -6.3 2.775 -6.265 2.912 ;
      RECT -6.31 2.765 -6.3 2.909 ;
      RECT -6.33 2.75 -6.31 2.907 ;
      RECT -6.36 2.72 -6.33 2.903 ;
      RECT -6.37 2.7 -6.36 2.898 ;
      RECT -6.375 2.692 -6.37 2.895 ;
      RECT -6.38 2.685 -6.375 2.893 ;
      RECT -6.395 2.672 -6.38 2.886 ;
      RECT -6.4 2.662 -6.395 2.878 ;
      RECT -6.405 2.655 -6.4 2.873 ;
      RECT -6.41 2.65 -6.405 2.869 ;
      RECT -6.425 2.637 -6.41 2.861 ;
      RECT -6.43 2.547 -6.425 2.85 ;
      RECT -6.435 2.542 -6.43 2.843 ;
      RECT -6.51 2.54 -6.435 2.803 ;
      RECT -6.54 2.54 -6.51 2.758 ;
      RECT -6.635 2.545 -6.62 2.745 ;
      RECT -4.15 2.25 -3.89 2.51 ;
      RECT -4.165 2.238 -3.985 2.475 ;
      RECT -4.17 2.239 -3.985 2.473 ;
      RECT -4.185 2.243 -3.975 2.463 ;
      RECT -4.19 2.248 -3.97 2.433 ;
      RECT -4.185 2.245 -3.97 2.463 ;
      RECT -4.17 2.24 -3.975 2.473 ;
      RECT -4.15 2.237 -3.985 2.51 ;
      RECT -4.15 2.236 -3.995 2.51 ;
      RECT -4.125 2.235 -3.995 2.51 ;
      RECT -4.565 2.48 -4.305 2.74 ;
      RECT -4.69 2.525 -4.305 2.735 ;
      RECT -4.7 2.53 -4.305 2.73 ;
      RECT -4.685 3.47 -4.67 3.78 ;
      RECT -6.09 3.24 -6.08 3.37 ;
      RECT -6.31 3.235 -6.205 3.37 ;
      RECT -6.395 3.24 -6.345 3.37 ;
      RECT -7.845 1.975 -7.84 3.08 ;
      RECT -4.59 3.562 -4.585 3.698 ;
      RECT -4.595 3.557 -4.59 3.758 ;
      RECT -4.6 3.555 -4.595 3.771 ;
      RECT -4.615 3.552 -4.6 3.773 ;
      RECT -4.62 3.547 -4.615 3.775 ;
      RECT -4.625 3.543 -4.62 3.778 ;
      RECT -4.64 3.538 -4.625 3.78 ;
      RECT -4.67 3.53 -4.64 3.78 ;
      RECT -4.709 3.47 -4.685 3.78 ;
      RECT -4.795 3.47 -4.709 3.777 ;
      RECT -4.825 3.47 -4.795 3.77 ;
      RECT -4.85 3.47 -4.825 3.763 ;
      RECT -4.875 3.47 -4.85 3.755 ;
      RECT -4.89 3.47 -4.875 3.748 ;
      RECT -4.915 3.47 -4.89 3.74 ;
      RECT -4.93 3.47 -4.915 3.733 ;
      RECT -4.97 3.48 -4.93 3.722 ;
      RECT -4.98 3.475 -4.97 3.712 ;
      RECT -4.984 3.474 -4.98 3.709 ;
      RECT -5.07 3.466 -4.984 3.692 ;
      RECT -5.103 3.455 -5.07 3.669 ;
      RECT -5.189 3.444 -5.103 3.647 ;
      RECT -5.275 3.428 -5.189 3.616 ;
      RECT -5.345 3.413 -5.275 3.588 ;
      RECT -5.355 3.406 -5.345 3.575 ;
      RECT -5.385 3.403 -5.355 3.565 ;
      RECT -5.41 3.399 -5.385 3.558 ;
      RECT -5.425 3.396 -5.41 3.553 ;
      RECT -5.43 3.395 -5.425 3.548 ;
      RECT -5.46 3.39 -5.43 3.541 ;
      RECT -5.465 3.385 -5.46 3.536 ;
      RECT -5.48 3.382 -5.465 3.531 ;
      RECT -5.485 3.377 -5.48 3.526 ;
      RECT -5.505 3.372 -5.485 3.523 ;
      RECT -5.52 3.367 -5.505 3.515 ;
      RECT -5.535 3.361 -5.52 3.51 ;
      RECT -5.565 3.352 -5.535 3.503 ;
      RECT -5.57 3.345 -5.565 3.495 ;
      RECT -5.575 3.343 -5.57 3.493 ;
      RECT -5.58 3.342 -5.575 3.49 ;
      RECT -5.62 3.335 -5.58 3.483 ;
      RECT -5.634 3.325 -5.62 3.473 ;
      RECT -5.685 3.314 -5.634 3.461 ;
      RECT -5.71 3.3 -5.685 3.447 ;
      RECT -5.735 3.289 -5.71 3.439 ;
      RECT -5.755 3.278 -5.735 3.433 ;
      RECT -5.765 3.272 -5.755 3.428 ;
      RECT -5.77 3.27 -5.765 3.424 ;
      RECT -5.79 3.265 -5.77 3.419 ;
      RECT -5.82 3.255 -5.79 3.409 ;
      RECT -5.825 3.247 -5.82 3.402 ;
      RECT -5.84 3.245 -5.825 3.398 ;
      RECT -5.86 3.245 -5.84 3.393 ;
      RECT -5.865 3.244 -5.86 3.391 ;
      RECT -5.87 3.244 -5.865 3.388 ;
      RECT -5.91 3.243 -5.87 3.383 ;
      RECT -5.935 3.242 -5.91 3.378 ;
      RECT -5.995 3.241 -5.935 3.375 ;
      RECT -6.08 3.24 -5.995 3.373 ;
      RECT -6.119 3.239 -6.09 3.37 ;
      RECT -6.205 3.237 -6.119 3.37 ;
      RECT -6.345 3.237 -6.31 3.37 ;
      RECT -6.435 3.241 -6.395 3.373 ;
      RECT -6.45 3.244 -6.435 3.38 ;
      RECT -6.46 3.245 -6.45 3.387 ;
      RECT -6.485 3.248 -6.46 3.392 ;
      RECT -6.49 3.25 -6.485 3.395 ;
      RECT -6.54 3.252 -6.49 3.396 ;
      RECT -6.579 3.256 -6.54 3.398 ;
      RECT -6.665 3.258 -6.579 3.401 ;
      RECT -6.683 3.26 -6.665 3.403 ;
      RECT -6.769 3.263 -6.683 3.405 ;
      RECT -6.855 3.267 -6.769 3.408 ;
      RECT -6.892 3.271 -6.855 3.411 ;
      RECT -6.978 3.274 -6.892 3.414 ;
      RECT -7.064 3.278 -6.978 3.417 ;
      RECT -7.15 3.283 -7.064 3.421 ;
      RECT -7.17 3.285 -7.15 3.424 ;
      RECT -7.19 3.284 -7.17 3.425 ;
      RECT -7.239 3.281 -7.19 3.426 ;
      RECT -7.325 3.276 -7.239 3.429 ;
      RECT -7.375 3.271 -7.325 3.431 ;
      RECT -7.399 3.269 -7.375 3.432 ;
      RECT -7.485 3.264 -7.399 3.434 ;
      RECT -7.51 3.26 -7.485 3.433 ;
      RECT -7.52 3.257 -7.51 3.431 ;
      RECT -7.53 3.25 -7.52 3.428 ;
      RECT -7.535 3.23 -7.53 3.423 ;
      RECT -7.545 3.2 -7.535 3.418 ;
      RECT -7.56 3.07 -7.545 3.409 ;
      RECT -7.565 3.062 -7.56 3.402 ;
      RECT -7.585 3.055 -7.565 3.394 ;
      RECT -7.59 3.037 -7.585 3.386 ;
      RECT -7.6 3.017 -7.59 3.381 ;
      RECT -7.605 2.99 -7.6 3.377 ;
      RECT -7.61 2.967 -7.605 3.374 ;
      RECT -7.63 2.925 -7.61 3.366 ;
      RECT -7.665 2.84 -7.63 3.35 ;
      RECT -7.67 2.772 -7.665 3.338 ;
      RECT -7.685 2.742 -7.67 3.332 ;
      RECT -7.69 1.987 -7.685 2.233 ;
      RECT -7.7 2.712 -7.685 3.323 ;
      RECT -7.695 1.982 -7.69 2.265 ;
      RECT -7.7 1.977 -7.695 2.308 ;
      RECT -7.705 1.975 -7.7 2.343 ;
      RECT -7.72 2.675 -7.7 3.313 ;
      RECT -7.71 1.975 -7.705 2.38 ;
      RECT -7.725 1.975 -7.71 2.478 ;
      RECT -7.725 2.648 -7.72 3.306 ;
      RECT -7.73 1.975 -7.725 2.553 ;
      RECT -7.73 2.636 -7.725 3.303 ;
      RECT -7.735 1.975 -7.73 2.585 ;
      RECT -7.735 2.615 -7.73 3.3 ;
      RECT -7.74 1.975 -7.735 3.297 ;
      RECT -7.775 1.975 -7.74 3.283 ;
      RECT -7.79 1.975 -7.775 3.265 ;
      RECT -7.81 1.975 -7.79 3.255 ;
      RECT -7.835 1.975 -7.81 3.238 ;
      RECT -7.84 1.975 -7.835 3.188 ;
      RECT -7.85 1.975 -7.845 3.018 ;
      RECT -7.855 1.975 -7.85 2.925 ;
      RECT -7.86 1.975 -7.855 2.838 ;
      RECT -7.865 1.975 -7.86 2.77 ;
      RECT -7.87 1.975 -7.865 2.713 ;
      RECT -7.88 1.975 -7.87 2.608 ;
      RECT -7.885 1.975 -7.88 2.48 ;
      RECT -7.89 1.975 -7.885 2.398 ;
      RECT -7.895 1.977 -7.89 2.315 ;
      RECT -7.9 1.982 -7.895 2.248 ;
      RECT -7.905 1.987 -7.9 2.175 ;
      RECT -5.09 2.305 -4.83 2.565 ;
      RECT -5.07 2.272 -4.86 2.565 ;
      RECT -5.07 2.27 -4.87 2.565 ;
      RECT -5.06 2.257 -4.87 2.565 ;
      RECT -5.06 2.255 -4.945 2.565 ;
      RECT -5.585 2.38 -5.41 2.66 ;
      RECT -5.59 2.38 -5.41 2.658 ;
      RECT -5.59 2.38 -5.395 2.655 ;
      RECT -5.6 2.38 -5.395 2.653 ;
      RECT -5.655 2.38 -5.395 2.64 ;
      RECT -5.655 2.455 -5.39 2.618 ;
      RECT -6.11 2.392 -6.09 2.635 ;
      RECT -6.11 2.392 -6.05 2.634 ;
      RECT -6.115 2.394 -6.05 2.633 ;
      RECT -6.115 2.394 -5.964 2.632 ;
      RECT -6.115 2.394 -5.895 2.631 ;
      RECT -6.115 2.394 -5.875 2.623 ;
      RECT -6.135 2.397 -5.875 2.621 ;
      RECT -6.15 2.407 -5.875 2.606 ;
      RECT -6.15 2.407 -5.86 2.605 ;
      RECT -6.155 2.416 -5.86 2.597 ;
      RECT -6.155 2.416 -5.855 2.593 ;
      RECT -6.05 2.33 -5.79 2.59 ;
      RECT -6.16 2.418 -5.79 2.475 ;
      RECT -6.09 2.385 -5.79 2.59 ;
      RECT -6.125 3.578 -6.12 3.785 ;
      RECT -6.175 3.572 -6.125 3.784 ;
      RECT -6.208 3.586 -6.115 3.783 ;
      RECT -6.294 3.586 -6.115 3.782 ;
      RECT -6.38 3.586 -6.115 3.781 ;
      RECT -6.38 3.685 -6.11 3.778 ;
      RECT -6.385 3.685 -6.11 3.773 ;
      RECT -6.39 3.685 -6.11 3.755 ;
      RECT -6.395 3.685 -6.11 3.738 ;
      RECT -6.435 3.47 -6.175 3.73 ;
      RECT -6.975 2.62 -6.889 3.034 ;
      RECT -6.975 2.62 -6.85 3.031 ;
      RECT -6.975 2.62 -6.83 3.021 ;
      RECT -7.02 2.62 -6.83 3.018 ;
      RECT -7.02 2.772 -6.82 3.008 ;
      RECT -7.02 2.793 -6.815 3.002 ;
      RECT -7.02 2.811 -6.81 2.998 ;
      RECT -7.02 2.831 -6.8 2.993 ;
      RECT -7.045 2.831 -6.8 2.99 ;
      RECT -7.055 2.831 -6.8 2.968 ;
      RECT -7.055 2.847 -6.795 2.938 ;
      RECT -7.09 2.62 -6.83 2.925 ;
      RECT -7.09 2.859 -6.79 2.88 ;
      RECT -8.825 8.575 6.435 8.88 ;
      RECT -4.505 3.265 -4.245 3.525 ;
    LAYER mcon ;
      RECT 5.895 0.915 6.065 1.085 ;
      RECT 5.895 2.395 6.065 2.565 ;
      RECT 5.895 6.315 6.065 6.485 ;
      RECT 5.895 7.795 6.065 7.965 ;
      RECT 5.545 0.105 5.715 0.275 ;
      RECT 5.545 4.165 5.715 4.335 ;
      RECT 5.545 4.545 5.715 4.715 ;
      RECT 5.545 8.605 5.715 8.775 ;
      RECT 5.525 2.765 5.695 2.935 ;
      RECT 5.525 5.945 5.695 6.115 ;
      RECT 4.905 0.915 5.075 1.085 ;
      RECT 4.905 2.395 5.075 2.565 ;
      RECT 4.905 6.315 5.075 6.485 ;
      RECT 4.905 7.795 5.075 7.965 ;
      RECT 4.555 0.105 4.725 0.275 ;
      RECT 4.555 4.165 4.725 4.335 ;
      RECT 4.555 4.545 4.725 4.715 ;
      RECT 4.555 8.605 4.725 8.775 ;
      RECT 4.535 2.765 4.705 2.935 ;
      RECT 4.535 5.945 4.705 6.115 ;
      RECT 3.85 0.105 4.02 0.275 ;
      RECT 3.85 4.165 4.02 4.335 ;
      RECT 3.85 4.545 4.02 4.715 ;
      RECT 3.85 8.605 4.02 8.775 ;
      RECT 3.54 2.025 3.71 2.195 ;
      RECT 3.54 6.685 3.71 6.855 ;
      RECT 3.17 0.105 3.34 0.275 ;
      RECT 3.17 8.605 3.34 8.775 ;
      RECT 3.11 0.915 3.28 1.085 ;
      RECT 3.11 1.655 3.28 1.825 ;
      RECT 3.11 7.055 3.28 7.225 ;
      RECT 3.11 7.795 3.28 7.965 ;
      RECT 2.735 2.395 2.905 2.565 ;
      RECT 2.735 6.315 2.905 6.485 ;
      RECT 2.49 0.105 2.66 0.275 ;
      RECT 2.49 8.605 2.66 8.775 ;
      RECT 1.81 0.105 1.98 0.275 ;
      RECT 1.81 8.605 1.98 8.775 ;
      RECT 1.74 2.765 1.91 2.935 ;
      RECT 1.74 5.945 1.91 6.115 ;
      RECT 0.35 1.415 0.52 1.585 ;
      RECT 0.35 4.135 0.52 4.305 ;
      RECT -0.09 2.28 0.08 2.45 ;
      RECT -0.11 1.415 0.06 1.585 ;
      RECT -0.11 4.135 0.06 4.305 ;
      RECT -0.485 3.025 -0.315 3.195 ;
      RECT -0.57 1.415 -0.4 1.585 ;
      RECT -0.57 4.135 -0.4 4.305 ;
      RECT -0.595 2.3 -0.425 2.47 ;
      RECT -1.03 1.415 -0.86 1.585 ;
      RECT -1.03 4.135 -0.86 4.305 ;
      RECT -1.415 1.99 -1.245 2.16 ;
      RECT -1.49 1.415 -1.32 1.585 ;
      RECT -1.49 4.135 -1.32 4.305 ;
      RECT -1.73 3.03 -1.56 3.2 ;
      RECT -1.775 2.52 -1.605 2.69 ;
      RECT -1.95 1.415 -1.78 1.585 ;
      RECT -1.95 4.135 -1.78 4.305 ;
      RECT -2.2 2.73 -2.03 2.9 ;
      RECT -2.39 1.95 -2.22 2.12 ;
      RECT -2.41 1.415 -2.24 1.585 ;
      RECT -2.41 4.135 -2.24 4.305 ;
      RECT -2.44 3.56 -2.27 3.73 ;
      RECT -2.775 3 -2.605 3.17 ;
      RECT -2.87 1.415 -2.7 1.585 ;
      RECT -2.87 2.16 -2.7 2.33 ;
      RECT -2.87 4.135 -2.7 4.305 ;
      RECT -3.33 1.415 -3.16 1.585 ;
      RECT -3.33 4.135 -3.16 4.305 ;
      RECT -3.67 3.385 -3.5 3.555 ;
      RECT -3.73 2.585 -3.56 2.755 ;
      RECT -3.79 1.415 -3.62 1.585 ;
      RECT -3.79 4.135 -3.62 4.305 ;
      RECT -4.17 2.255 -4 2.425 ;
      RECT -4.25 1.415 -4.08 1.585 ;
      RECT -4.25 4.135 -4.08 4.305 ;
      RECT -4.435 3.305 -4.265 3.475 ;
      RECT -4.68 2.545 -4.51 2.715 ;
      RECT -4.71 1.415 -4.54 1.585 ;
      RECT -4.71 4.135 -4.54 4.305 ;
      RECT -4.775 3.575 -4.605 3.745 ;
      RECT -5.05 2.27 -4.88 2.44 ;
      RECT -5.17 1.415 -5 1.585 ;
      RECT -5.17 4.135 -5 4.305 ;
      RECT -5.58 2.47 -5.41 2.64 ;
      RECT -5.63 1.415 -5.46 1.585 ;
      RECT -5.63 4.135 -5.46 4.305 ;
      RECT -6.09 1.415 -5.92 1.585 ;
      RECT -6.09 4.135 -5.92 4.305 ;
      RECT -6.1 2.415 -5.93 2.585 ;
      RECT -6.305 2.015 -6.135 2.185 ;
      RECT -6.305 3.595 -6.135 3.765 ;
      RECT -6.55 1.415 -6.38 1.585 ;
      RECT -6.55 4.135 -6.38 4.305 ;
      RECT -6.615 2.56 -6.445 2.73 ;
      RECT -7.01 1.415 -6.84 1.585 ;
      RECT -7.01 4.135 -6.84 4.305 ;
      RECT -7.025 2.785 -6.855 2.955 ;
      RECT -7.47 1.415 -7.3 1.585 ;
      RECT -7.47 4.135 -7.3 4.305 ;
      RECT -7.735 3.085 -7.565 3.255 ;
      RECT -7.88 1.995 -7.71 2.165 ;
      RECT -7.93 1.415 -7.76 1.585 ;
      RECT -7.93 4.135 -7.76 4.305 ;
    LAYER li ;
      RECT -0.105 0 0.065 2.085 ;
      RECT -1.045 0 -0.875 2.085 ;
      RECT -2.005 0 -1.835 2.085 ;
      RECT -3.925 0 -3.755 2.085 ;
      RECT -4.885 0 -4.715 2.085 ;
      RECT -6.805 0 -6.635 2.085 ;
      RECT -3.05 0 -2.855 1.595 ;
      RECT -6.805 0 -6.53 1.595 ;
      RECT -8.075 0 0.665 1.585 ;
      RECT 5.465 0 5.635 0.935 ;
      RECT 4.475 0 4.645 0.935 ;
      RECT 1.73 0 1.9 0.935 ;
      RECT -8.825 0 6.435 0.305 ;
      RECT 5.465 3.405 5.635 5.475 ;
      RECT 4.475 3.405 4.645 5.475 ;
      RECT 1.73 3.405 1.9 5.475 ;
      RECT -8.825 4.14 6.435 4.745 ;
      RECT -8.075 4.135 6.435 4.745 ;
      RECT -1.045 3.635 -0.875 4.745 ;
      RECT -2.965 3.635 -2.795 4.745 ;
      RECT -3.905 3.635 -3.735 4.745 ;
      RECT -5.365 3.635 -5.195 4.745 ;
      RECT -7.285 3.635 -7.115 4.745 ;
      RECT -8.825 8.575 6.435 8.88 ;
      RECT 5.465 7.945 5.635 8.88 ;
      RECT 4.475 7.945 4.645 8.88 ;
      RECT 1.73 7.945 1.9 8.88 ;
      RECT 5.525 1.74 5.695 2.935 ;
      RECT 5.525 1.74 5.99 1.91 ;
      RECT 5.525 6.97 5.99 7.14 ;
      RECT 5.525 5.945 5.695 7.14 ;
      RECT 4.535 1.74 4.705 2.935 ;
      RECT 4.535 1.74 5 1.91 ;
      RECT 4.535 6.97 5 7.14 ;
      RECT 4.535 5.945 4.705 7.14 ;
      RECT 2.68 2.635 2.85 3.865 ;
      RECT 2.735 0.855 2.905 2.805 ;
      RECT 2.68 0.575 2.85 1.025 ;
      RECT 2.68 7.855 2.85 8.305 ;
      RECT 2.735 6.075 2.905 8.025 ;
      RECT 2.68 5.015 2.85 6.245 ;
      RECT 2.16 0.575 2.33 3.865 ;
      RECT 2.16 2.075 2.565 2.405 ;
      RECT 2.16 1.235 2.565 1.565 ;
      RECT 2.16 5.015 2.33 8.305 ;
      RECT 2.16 7.315 2.565 7.645 ;
      RECT 2.16 6.475 2.565 6.805 ;
      RECT 0.085 3.126 0.09 3.298 ;
      RECT 0.08 3.119 0.085 3.388 ;
      RECT 0.075 3.113 0.08 3.407 ;
      RECT 0.055 3.107 0.075 3.417 ;
      RECT 0.04 3.102 0.055 3.425 ;
      RECT 0.003 3.096 0.04 3.423 ;
      RECT -0.083 3.082 0.003 3.419 ;
      RECT -0.169 3.064 -0.083 3.414 ;
      RECT -0.255 3.045 -0.169 3.408 ;
      RECT -0.285 3.033 -0.255 3.404 ;
      RECT -0.305 3.027 -0.285 3.403 ;
      RECT -0.37 3.025 -0.305 3.401 ;
      RECT -0.385 3.025 -0.37 3.393 ;
      RECT -0.4 3.025 -0.385 3.38 ;
      RECT -0.405 3.025 -0.4 3.37 ;
      RECT -0.42 3.025 -0.405 3.348 ;
      RECT -0.435 3.025 -0.42 3.315 ;
      RECT -0.44 3.025 -0.435 3.293 ;
      RECT -0.45 3.025 -0.44 3.275 ;
      RECT -0.465 3.025 -0.45 3.253 ;
      RECT -0.485 3.025 -0.465 3.215 ;
      RECT -0.135 2.31 -0.1 2.749 ;
      RECT -0.135 2.31 -0.095 2.748 ;
      RECT -0.19 2.37 -0.095 2.747 ;
      RECT -0.325 2.542 -0.095 2.746 ;
      RECT -0.215 2.42 -0.095 2.746 ;
      RECT -0.325 2.542 -0.07 2.736 ;
      RECT -0.27 2.487 0.01 2.653 ;
      RECT -0.095 2.281 -0.09 2.744 ;
      RECT -0.24 2.457 0.05 2.53 ;
      RECT -0.225 2.44 -0.095 2.746 ;
      RECT -0.09 2.28 0.08 2.468 ;
      RECT -0.1 2.283 0.08 2.468 ;
      RECT -0.595 2.16 -0.425 2.47 ;
      RECT -0.595 2.16 -0.42 2.443 ;
      RECT -0.595 2.16 -0.415 2.42 ;
      RECT -0.595 2.16 -0.405 2.37 ;
      RECT -0.6 2.265 -0.405 2.34 ;
      RECT -0.565 1.835 -0.395 2.313 ;
      RECT -0.565 1.835 -0.38 2.234 ;
      RECT -0.575 2.045 -0.38 2.234 ;
      RECT -0.565 1.845 -0.37 2.149 ;
      RECT -0.635 2.587 -0.63 2.79 ;
      RECT -0.645 2.575 -0.635 2.9 ;
      RECT -0.67 2.575 -0.645 2.94 ;
      RECT -0.75 2.575 -0.67 3.025 ;
      RECT -0.76 2.575 -0.75 3.095 ;
      RECT -0.785 2.575 -0.76 3.118 ;
      RECT -0.805 2.575 -0.785 3.153 ;
      RECT -0.85 2.585 -0.805 3.196 ;
      RECT -0.86 2.597 -0.85 3.233 ;
      RECT -0.88 2.611 -0.86 3.253 ;
      RECT -0.89 2.629 -0.88 3.269 ;
      RECT -0.905 2.655 -0.89 3.279 ;
      RECT -0.92 2.696 -0.905 3.293 ;
      RECT -0.93 2.731 -0.92 3.303 ;
      RECT -0.935 2.747 -0.93 3.308 ;
      RECT -0.945 2.762 -0.935 3.313 ;
      RECT -0.965 2.805 -0.945 3.323 ;
      RECT -0.985 2.842 -0.965 3.336 ;
      RECT -1.02 2.865 -0.985 3.354 ;
      RECT -1.03 2.879 -1.02 3.37 ;
      RECT -1.05 2.889 -1.03 3.38 ;
      RECT -1.055 2.898 -1.05 3.388 ;
      RECT -1.065 2.905 -1.055 3.395 ;
      RECT -1.075 2.912 -1.065 3.403 ;
      RECT -1.09 2.922 -1.075 3.411 ;
      RECT -1.1 2.936 -1.09 3.421 ;
      RECT -1.11 2.948 -1.1 3.433 ;
      RECT -1.125 2.97 -1.11 3.446 ;
      RECT -1.135 2.992 -1.125 3.457 ;
      RECT -1.145 3.012 -1.135 3.466 ;
      RECT -1.15 3.027 -1.145 3.473 ;
      RECT -1.18 3.06 -1.15 3.487 ;
      RECT -1.19 3.095 -1.18 3.502 ;
      RECT -1.195 3.102 -1.19 3.508 ;
      RECT -1.215 3.117 -1.195 3.515 ;
      RECT -1.22 3.132 -1.215 3.523 ;
      RECT -1.225 3.141 -1.22 3.528 ;
      RECT -1.24 3.147 -1.225 3.535 ;
      RECT -1.245 3.153 -1.24 3.543 ;
      RECT -1.25 3.157 -1.245 3.55 ;
      RECT -1.255 3.161 -1.25 3.56 ;
      RECT -1.265 3.166 -1.255 3.57 ;
      RECT -1.285 3.177 -1.265 3.598 ;
      RECT -1.3 3.189 -1.285 3.625 ;
      RECT -1.32 3.202 -1.3 3.65 ;
      RECT -1.34 3.217 -1.32 3.674 ;
      RECT -1.355 3.232 -1.34 3.689 ;
      RECT -1.36 3.243 -1.355 3.698 ;
      RECT -1.425 3.288 -1.36 3.708 ;
      RECT -1.46 3.347 -1.425 3.721 ;
      RECT -1.465 3.37 -1.46 3.727 ;
      RECT -1.47 3.377 -1.465 3.729 ;
      RECT -1.485 3.387 -1.47 3.732 ;
      RECT -1.515 3.412 -1.485 3.736 ;
      RECT -1.52 3.43 -1.515 3.74 ;
      RECT -1.525 3.437 -1.52 3.741 ;
      RECT -1.545 3.445 -1.525 3.745 ;
      RECT -1.555 3.452 -1.545 3.749 ;
      RECT -1.599 3.463 -1.555 3.756 ;
      RECT -1.685 3.491 -1.599 3.772 ;
      RECT -1.745 3.515 -1.685 3.79 ;
      RECT -1.79 3.525 -1.745 3.804 ;
      RECT -1.849 3.533 -1.79 3.818 ;
      RECT -1.935 3.54 -1.849 3.837 ;
      RECT -1.96 3.545 -1.935 3.852 ;
      RECT -2.04 3.548 -1.96 3.855 ;
      RECT -2.12 3.552 -2.04 3.842 ;
      RECT -2.129 3.555 -2.12 3.827 ;
      RECT -2.215 3.555 -2.129 3.812 ;
      RECT -2.275 3.557 -2.215 3.789 ;
      RECT -2.279 3.56 -2.275 3.779 ;
      RECT -2.365 3.56 -2.279 3.764 ;
      RECT -2.44 3.56 -2.365 3.74 ;
      RECT -1.125 2.569 -1.115 2.745 ;
      RECT -1.17 2.536 -1.125 2.745 ;
      RECT -1.215 2.487 -1.17 2.745 ;
      RECT -1.245 2.457 -1.215 2.746 ;
      RECT -1.25 2.44 -1.245 2.747 ;
      RECT -1.275 2.42 -1.25 2.748 ;
      RECT -1.29 2.395 -1.275 2.749 ;
      RECT -1.295 2.382 -1.29 2.75 ;
      RECT -1.3 2.376 -1.295 2.748 ;
      RECT -1.305 2.368 -1.3 2.742 ;
      RECT -1.33 2.36 -1.305 2.722 ;
      RECT -1.35 2.349 -1.33 2.693 ;
      RECT -1.38 2.334 -1.35 2.664 ;
      RECT -1.4 2.32 -1.38 2.636 ;
      RECT -1.41 2.314 -1.4 2.615 ;
      RECT -1.415 2.311 -1.41 2.598 ;
      RECT -1.42 2.308 -1.415 2.583 ;
      RECT -1.435 2.303 -1.42 2.548 ;
      RECT -1.44 2.299 -1.435 2.515 ;
      RECT -1.46 2.294 -1.44 2.491 ;
      RECT -1.49 2.286 -1.46 2.456 ;
      RECT -1.505 2.28 -1.49 2.433 ;
      RECT -1.545 2.273 -1.505 2.418 ;
      RECT -1.57 2.265 -1.545 2.398 ;
      RECT -1.59 2.26 -1.57 2.388 ;
      RECT -1.625 2.254 -1.59 2.383 ;
      RECT -1.67 2.245 -1.625 2.382 ;
      RECT -1.7 2.241 -1.67 2.384 ;
      RECT -1.785 2.249 -1.7 2.388 ;
      RECT -1.855 2.26 -1.785 2.41 ;
      RECT -1.868 2.266 -1.855 2.433 ;
      RECT -1.954 2.273 -1.868 2.455 ;
      RECT -2.04 2.285 -1.954 2.492 ;
      RECT -2.04 2.662 -2.03 2.9 ;
      RECT -2.045 2.291 -2.04 2.515 ;
      RECT -2.05 2.547 -2.04 2.9 ;
      RECT -2.05 2.292 -2.045 2.52 ;
      RECT -2.055 2.293 -2.05 2.9 ;
      RECT -2.079 2.295 -2.055 2.901 ;
      RECT -2.165 2.303 -2.079 2.903 ;
      RECT -2.185 2.317 -2.165 2.906 ;
      RECT -2.19 2.345 -2.185 2.907 ;
      RECT -2.195 2.357 -2.19 2.908 ;
      RECT -2.2 2.372 -2.195 2.909 ;
      RECT -2.21 2.402 -2.2 2.91 ;
      RECT -2.215 2.44 -2.21 2.908 ;
      RECT -2.22 2.46 -2.215 2.903 ;
      RECT -2.235 2.495 -2.22 2.888 ;
      RECT -2.245 2.547 -2.235 2.868 ;
      RECT -2.25 2.577 -2.245 2.856 ;
      RECT -2.265 2.59 -2.25 2.839 ;
      RECT -2.29 2.594 -2.265 2.806 ;
      RECT -2.305 2.592 -2.29 2.783 ;
      RECT -2.32 2.591 -2.305 2.78 ;
      RECT -2.38 2.589 -2.32 2.778 ;
      RECT -2.39 2.587 -2.38 2.773 ;
      RECT -2.43 2.586 -2.39 2.77 ;
      RECT -2.5 2.583 -2.43 2.768 ;
      RECT -2.555 2.581 -2.5 2.763 ;
      RECT -2.625 2.575 -2.555 2.758 ;
      RECT -2.634 2.575 -2.625 2.755 ;
      RECT -2.72 2.575 -2.634 2.75 ;
      RECT -2.725 2.575 -2.72 2.745 ;
      RECT -1.42 1.81 -1.245 2.16 ;
      RECT -1.42 1.825 -1.235 2.158 ;
      RECT -1.445 1.775 -1.3 2.155 ;
      RECT -1.465 1.776 -1.3 2.148 ;
      RECT -1.475 1.777 -1.29 2.143 ;
      RECT -1.505 1.778 -1.29 2.13 ;
      RECT -1.555 1.779 -1.29 2.106 ;
      RECT -1.56 1.781 -1.29 2.091 ;
      RECT -1.56 1.847 -1.23 2.085 ;
      RECT -1.58 1.788 -1.275 2.065 ;
      RECT -1.59 1.797 -1.265 1.92 ;
      RECT -1.58 1.792 -1.265 2.065 ;
      RECT -1.56 1.782 -1.275 2.091 ;
      RECT -1.975 3.107 -1.805 3.395 ;
      RECT -1.98 3.125 -1.795 3.39 ;
      RECT -2.015 3.133 -1.73 3.31 ;
      RECT -2.015 3.133 -1.644 3.3 ;
      RECT -2.015 3.133 -1.59 3.246 ;
      RECT -1.73 3.03 -1.56 3.214 ;
      RECT -2.015 3.185 -1.555 3.202 ;
      RECT -2.03 3.155 -1.56 3.198 ;
      RECT -1.77 3.037 -1.73 3.349 ;
      RECT -1.89 3.074 -1.56 3.214 ;
      RECT -1.795 3.049 -1.77 3.375 ;
      RECT -1.805 3.056 -1.56 3.214 ;
      RECT -1.674 2.52 -1.605 2.779 ;
      RECT -1.674 2.575 -1.6 2.778 ;
      RECT -1.76 2.575 -1.6 2.777 ;
      RECT -1.765 2.575 -1.595 2.77 ;
      RECT -1.775 2.52 -1.605 2.765 ;
      RECT -2.395 1.819 -2.22 2.12 ;
      RECT -2.41 1.807 -2.395 2.105 ;
      RECT -2.44 1.806 -2.41 2.058 ;
      RECT -2.44 1.824 -2.215 2.053 ;
      RECT -2.455 1.808 -2.395 2.018 ;
      RECT -2.46 1.83 -2.205 1.918 ;
      RECT -2.46 1.813 -2.309 1.918 ;
      RECT -2.46 1.815 -2.305 1.918 ;
      RECT -2.455 1.811 -2.309 2.018 ;
      RECT -2.35 3.047 -2.345 3.395 ;
      RECT -2.36 3.037 -2.35 3.401 ;
      RECT -2.395 3.027 -2.36 3.403 ;
      RECT -2.433 3.022 -2.395 3.407 ;
      RECT -2.519 3.015 -2.433 3.414 ;
      RECT -2.605 3.005 -2.519 3.424 ;
      RECT -2.65 3 -2.605 3.432 ;
      RECT -2.654 3 -2.65 3.436 ;
      RECT -2.74 3 -2.654 3.443 ;
      RECT -2.755 3 -2.74 3.443 ;
      RECT -2.765 2.998 -2.755 3.415 ;
      RECT -2.775 2.994 -2.765 3.358 ;
      RECT -2.795 2.988 -2.775 3.29 ;
      RECT -2.8 2.984 -2.795 3.238 ;
      RECT -2.81 2.983 -2.8 3.205 ;
      RECT -2.86 2.981 -2.81 3.19 ;
      RECT -2.885 2.979 -2.86 3.185 ;
      RECT -2.928 2.977 -2.885 3.181 ;
      RECT -3.014 2.973 -2.928 3.169 ;
      RECT -3.1 2.968 -3.014 3.153 ;
      RECT -3.13 2.965 -3.1 3.14 ;
      RECT -3.155 2.964 -3.13 3.128 ;
      RECT -3.16 2.964 -3.155 3.118 ;
      RECT -3.2 2.963 -3.16 3.11 ;
      RECT -3.215 2.962 -3.2 3.103 ;
      RECT -3.265 2.961 -3.215 3.095 ;
      RECT -3.267 2.96 -3.265 3.09 ;
      RECT -3.353 2.958 -3.267 3.09 ;
      RECT -3.439 2.953 -3.353 3.09 ;
      RECT -3.525 2.949 -3.439 3.09 ;
      RECT -3.574 2.945 -3.525 3.088 ;
      RECT -3.66 2.942 -3.574 3.083 ;
      RECT -3.683 2.939 -3.66 3.079 ;
      RECT -3.769 2.936 -3.683 3.074 ;
      RECT -3.855 2.932 -3.769 3.065 ;
      RECT -3.88 2.925 -3.855 3.06 ;
      RECT -3.94 2.89 -3.88 3.057 ;
      RECT -3.96 2.815 -3.94 3.054 ;
      RECT -3.965 2.757 -3.96 3.053 ;
      RECT -3.99 2.697 -3.965 3.052 ;
      RECT -4.065 2.575 -3.99 3.048 ;
      RECT -4.075 2.575 -4.065 3.04 ;
      RECT -4.09 2.575 -4.075 3.03 ;
      RECT -4.105 2.575 -4.09 3 ;
      RECT -4.12 2.575 -4.105 2.945 ;
      RECT -4.135 2.575 -4.12 2.883 ;
      RECT -4.16 2.575 -4.135 2.808 ;
      RECT -4.165 2.575 -4.16 2.758 ;
      RECT -2.82 2.12 -2.8 2.429 ;
      RECT -2.834 2.122 -2.785 2.426 ;
      RECT -2.834 2.127 -2.765 2.417 ;
      RECT -2.92 2.125 -2.785 2.411 ;
      RECT -2.92 2.133 -2.73 2.394 ;
      RECT -2.955 2.135 -2.73 2.393 ;
      RECT -2.985 2.143 -2.73 2.384 ;
      RECT -2.995 2.148 -2.71 2.37 ;
      RECT -2.955 2.138 -2.71 2.37 ;
      RECT -2.955 2.141 -2.7 2.358 ;
      RECT -2.985 2.143 -2.69 2.345 ;
      RECT -2.985 2.147 -2.68 2.288 ;
      RECT -2.995 2.152 -2.675 2.203 ;
      RECT -2.834 2.12 -2.8 2.426 ;
      RECT -3.395 2.223 -3.39 2.435 ;
      RECT -3.52 2.22 -3.505 2.435 ;
      RECT -4.055 2.25 -3.985 2.435 ;
      RECT -4.17 2.25 -4.135 2.43 ;
      RECT -3.049 2.552 -3.03 2.746 ;
      RECT -3.135 2.507 -3.049 2.747 ;
      RECT -3.145 2.46 -3.135 2.749 ;
      RECT -3.15 2.44 -3.145 2.75 ;
      RECT -3.17 2.405 -3.15 2.751 ;
      RECT -3.185 2.355 -3.17 2.752 ;
      RECT -3.205 2.292 -3.185 2.753 ;
      RECT -3.215 2.255 -3.205 2.754 ;
      RECT -3.23 2.244 -3.215 2.755 ;
      RECT -3.235 2.236 -3.23 2.753 ;
      RECT -3.245 2.235 -3.235 2.745 ;
      RECT -3.275 2.232 -3.245 2.724 ;
      RECT -3.35 2.227 -3.275 2.669 ;
      RECT -3.365 2.223 -3.35 2.615 ;
      RECT -3.375 2.223 -3.365 2.51 ;
      RECT -3.39 2.223 -3.375 2.443 ;
      RECT -3.405 2.223 -3.395 2.433 ;
      RECT -3.46 2.222 -3.405 2.43 ;
      RECT -3.505 2.22 -3.46 2.433 ;
      RECT -3.533 2.22 -3.52 2.436 ;
      RECT -3.619 2.224 -3.533 2.438 ;
      RECT -3.705 2.23 -3.619 2.443 ;
      RECT -3.725 2.234 -3.705 2.445 ;
      RECT -3.727 2.235 -3.725 2.444 ;
      RECT -3.813 2.237 -3.727 2.443 ;
      RECT -3.899 2.242 -3.813 2.44 ;
      RECT -3.985 2.247 -3.899 2.437 ;
      RECT -4.135 2.25 -4.055 2.433 ;
      RECT -3.359 3.225 -3.31 3.559 ;
      RECT -3.359 3.225 -3.305 3.558 ;
      RECT -3.445 3.225 -3.305 3.557 ;
      RECT -3.67 3.333 -3.3 3.555 ;
      RECT -3.445 3.225 -3.275 3.548 ;
      RECT -3.475 3.237 -3.27 3.539 ;
      RECT -3.49 3.255 -3.265 3.536 ;
      RECT -3.675 3.339 -3.265 3.463 ;
      RECT -3.68 3.346 -3.265 3.423 ;
      RECT -3.665 3.312 -3.265 3.536 ;
      RECT -3.504 3.258 -3.3 3.555 ;
      RECT -3.59 3.278 -3.265 3.536 ;
      RECT -3.49 3.252 -3.27 3.539 ;
      RECT -3.72 2.576 -3.53 2.77 ;
      RECT -3.725 2.578 -3.53 2.769 ;
      RECT -3.73 2.582 -3.515 2.766 ;
      RECT -3.715 2.575 -3.515 2.766 ;
      RECT -3.73 2.685 -3.51 2.761 ;
      RECT -4.435 3.185 -4.344 3.483 ;
      RECT -4.44 3.187 -4.265 3.478 ;
      RECT -4.435 3.185 -4.265 3.478 ;
      RECT -4.44 3.191 -4.245 3.476 ;
      RECT -4.44 3.246 -4.205 3.475 ;
      RECT -4.44 3.281 -4.19 3.469 ;
      RECT -4.44 3.315 -4.18 3.459 ;
      RECT -4.45 3.195 -4.245 3.31 ;
      RECT -4.45 3.215 -4.23 3.31 ;
      RECT -4.45 3.198 -4.24 3.31 ;
      RECT -4.225 1.966 -4.22 2.028 ;
      RECT -4.23 1.888 -4.225 2.051 ;
      RECT -4.235 1.845 -4.23 2.062 ;
      RECT -4.24 1.835 -4.235 2.074 ;
      RECT -4.245 1.835 -4.24 2.083 ;
      RECT -4.27 1.835 -4.245 2.115 ;
      RECT -4.275 1.835 -4.27 2.148 ;
      RECT -4.29 1.835 -4.275 2.173 ;
      RECT -4.3 1.835 -4.29 2.2 ;
      RECT -4.305 1.835 -4.3 2.213 ;
      RECT -4.31 1.835 -4.305 2.228 ;
      RECT -4.32 1.835 -4.31 2.243 ;
      RECT -4.325 1.835 -4.32 2.263 ;
      RECT -4.35 1.835 -4.325 2.298 ;
      RECT -4.395 1.835 -4.35 2.343 ;
      RECT -4.405 1.835 -4.395 2.356 ;
      RECT -4.49 1.92 -4.405 2.363 ;
      RECT -4.525 2.042 -4.49 2.372 ;
      RECT -4.53 2.082 -4.525 2.376 ;
      RECT -4.55 2.105 -4.53 2.378 ;
      RECT -4.555 2.135 -4.55 2.381 ;
      RECT -4.565 2.147 -4.555 2.382 ;
      RECT -4.61 2.17 -4.565 2.387 ;
      RECT -4.65 2.2 -4.61 2.395 ;
      RECT -4.685 2.212 -4.65 2.401 ;
      RECT -4.69 2.217 -4.685 2.405 ;
      RECT -4.76 2.227 -4.69 2.412 ;
      RECT -4.8 2.237 -4.76 2.422 ;
      RECT -4.82 2.242 -4.8 2.428 ;
      RECT -4.83 2.246 -4.82 2.433 ;
      RECT -4.835 2.249 -4.83 2.436 ;
      RECT -4.845 2.25 -4.835 2.437 ;
      RECT -4.87 2.252 -4.845 2.441 ;
      RECT -4.88 2.257 -4.87 2.444 ;
      RECT -4.925 2.265 -4.88 2.445 ;
      RECT -5.05 2.27 -4.925 2.445 ;
      RECT -4.495 2.567 -4.475 2.749 ;
      RECT -4.544 2.552 -4.495 2.748 ;
      RECT -4.63 2.567 -4.475 2.746 ;
      RECT -4.645 2.567 -4.475 2.745 ;
      RECT -4.68 2.545 -4.51 2.73 ;
      RECT -4.61 3.565 -4.595 3.774 ;
      RECT -4.61 3.573 -4.59 3.773 ;
      RECT -4.665 3.573 -4.59 3.772 ;
      RECT -4.685 3.577 -4.585 3.77 ;
      RECT -4.705 3.527 -4.665 3.769 ;
      RECT -4.76 3.585 -4.58 3.767 ;
      RECT -4.795 3.542 -4.665 3.765 ;
      RECT -4.799 3.545 -4.61 3.764 ;
      RECT -4.885 3.553 -4.61 3.762 ;
      RECT -4.885 3.597 -4.575 3.755 ;
      RECT -4.895 3.69 -4.575 3.753 ;
      RECT -4.885 3.609 -4.57 3.738 ;
      RECT -4.885 3.63 -4.555 3.708 ;
      RECT -4.885 3.657 -4.55 3.678 ;
      RECT -4.76 3.535 -4.665 3.767 ;
      RECT -5.13 2.58 -5.125 3.118 ;
      RECT -5.325 2.91 -5.32 3.105 ;
      RECT -7.025 2.575 -7.01 2.955 ;
      RECT -4.96 2.575 -4.955 2.745 ;
      RECT -4.965 2.575 -4.96 2.755 ;
      RECT -4.97 2.575 -4.965 2.768 ;
      RECT -4.995 2.575 -4.97 2.81 ;
      RECT -5.02 2.575 -4.995 2.883 ;
      RECT -5.035 2.575 -5.02 2.935 ;
      RECT -5.04 2.575 -5.035 2.965 ;
      RECT -5.065 2.575 -5.04 3.005 ;
      RECT -5.08 2.575 -5.065 3.06 ;
      RECT -5.085 2.575 -5.08 3.093 ;
      RECT -5.11 2.575 -5.085 3.113 ;
      RECT -5.125 2.575 -5.11 3.119 ;
      RECT -5.195 2.61 -5.13 3.115 ;
      RECT -5.245 2.665 -5.195 3.11 ;
      RECT -5.255 2.697 -5.245 3.108 ;
      RECT -5.26 2.722 -5.255 3.108 ;
      RECT -5.28 2.795 -5.26 3.108 ;
      RECT -5.29 2.875 -5.28 3.107 ;
      RECT -5.305 2.905 -5.29 3.107 ;
      RECT -5.32 2.91 -5.305 3.106 ;
      RECT -5.38 2.912 -5.325 3.103 ;
      RECT -5.41 2.917 -5.38 3.099 ;
      RECT -5.412 2.92 -5.41 3.098 ;
      RECT -5.498 2.922 -5.412 3.095 ;
      RECT -5.584 2.928 -5.498 3.089 ;
      RECT -5.67 2.933 -5.584 3.083 ;
      RECT -5.743 2.938 -5.67 3.084 ;
      RECT -5.829 2.944 -5.743 3.092 ;
      RECT -5.915 2.95 -5.829 3.101 ;
      RECT -5.935 2.954 -5.915 3.106 ;
      RECT -5.982 2.956 -5.935 3.109 ;
      RECT -6.068 2.961 -5.982 3.115 ;
      RECT -6.154 2.966 -6.068 3.124 ;
      RECT -6.24 2.972 -6.154 3.132 ;
      RECT -6.325 2.97 -6.24 3.141 ;
      RECT -6.329 2.965 -6.325 3.145 ;
      RECT -6.415 2.96 -6.329 3.137 ;
      RECT -6.479 2.951 -6.415 3.125 ;
      RECT -6.565 2.942 -6.479 3.112 ;
      RECT -6.589 2.935 -6.565 3.103 ;
      RECT -6.675 2.929 -6.589 3.09 ;
      RECT -6.715 2.922 -6.675 3.076 ;
      RECT -6.72 2.912 -6.715 3.072 ;
      RECT -6.73 2.9 -6.72 3.071 ;
      RECT -6.75 2.87 -6.73 3.068 ;
      RECT -6.805 2.79 -6.75 3.062 ;
      RECT -6.825 2.709 -6.805 3.057 ;
      RECT -6.845 2.667 -6.825 3.053 ;
      RECT -6.87 2.62 -6.845 3.047 ;
      RECT -6.875 2.595 -6.87 3.044 ;
      RECT -6.91 2.575 -6.875 3.039 ;
      RECT -6.919 2.575 -6.91 3.032 ;
      RECT -7.005 2.575 -6.919 3.002 ;
      RECT -7.01 2.575 -7.005 2.965 ;
      RECT -7.045 2.575 -7.025 2.887 ;
      RECT -7.05 2.617 -7.045 2.852 ;
      RECT -7.055 2.692 -7.05 2.808 ;
      RECT -5.605 2.497 -5.43 2.745 ;
      RECT -5.605 2.497 -5.425 2.743 ;
      RECT -5.61 2.529 -5.425 2.703 ;
      RECT -5.58 2.47 -5.41 2.69 ;
      RECT -5.615 2.547 -5.41 2.623 ;
      RECT -6.305 2.01 -6.135 2.185 ;
      RECT -6.305 2.01 -5.963 2.177 ;
      RECT -6.305 2.01 -5.88 2.171 ;
      RECT -6.305 2.01 -5.845 2.167 ;
      RECT -6.305 2.01 -5.825 2.166 ;
      RECT -6.305 2.01 -5.739 2.162 ;
      RECT -5.845 1.835 -5.675 2.157 ;
      RECT -6.27 1.942 -5.645 2.155 ;
      RECT -6.28 1.997 -5.64 2.153 ;
      RECT -6.305 2.033 -5.63 2.148 ;
      RECT -6.305 2.06 -5.625 2.078 ;
      RECT -6.24 1.885 -5.665 2.155 ;
      RECT -6.049 1.87 -5.665 2.155 ;
      RECT -6.215 1.873 -5.665 2.155 ;
      RECT -6.135 1.871 -6.049 2.182 ;
      RECT -6.049 1.868 -5.67 2.155 ;
      RECT -5.865 1.845 -5.67 2.155 ;
      RECT -5.963 1.866 -5.67 2.155 ;
      RECT -5.88 1.86 -5.865 2.168 ;
      RECT -5.73 3.225 -5.725 3.425 ;
      RECT -6.265 3.29 -6.22 3.425 ;
      RECT -5.695 3.225 -5.675 3.398 ;
      RECT -5.725 3.225 -5.695 3.413 ;
      RECT -5.79 3.225 -5.73 3.45 ;
      RECT -5.805 3.225 -5.79 3.48 ;
      RECT -5.82 3.225 -5.805 3.493 ;
      RECT -5.84 3.225 -5.82 3.508 ;
      RECT -5.845 3.225 -5.84 3.517 ;
      RECT -5.855 3.229 -5.845 3.522 ;
      RECT -5.87 3.239 -5.855 3.533 ;
      RECT -5.895 3.255 -5.87 3.543 ;
      RECT -5.905 3.269 -5.895 3.545 ;
      RECT -5.925 3.281 -5.905 3.542 ;
      RECT -5.955 3.302 -5.925 3.536 ;
      RECT -5.965 3.314 -5.955 3.531 ;
      RECT -5.975 3.312 -5.965 3.528 ;
      RECT -5.99 3.311 -5.975 3.523 ;
      RECT -5.995 3.31 -5.99 3.518 ;
      RECT -6.03 3.308 -5.995 3.508 ;
      RECT -6.05 3.305 -6.03 3.49 ;
      RECT -6.06 3.303 -6.05 3.485 ;
      RECT -6.07 3.302 -6.06 3.48 ;
      RECT -6.105 3.3 -6.07 3.468 ;
      RECT -6.16 3.296 -6.105 3.448 ;
      RECT -6.17 3.294 -6.16 3.433 ;
      RECT -6.175 3.294 -6.17 3.428 ;
      RECT -6.22 3.292 -6.175 3.425 ;
      RECT -6.315 3.29 -6.265 3.429 ;
      RECT -6.325 3.291 -6.315 3.434 ;
      RECT -6.385 3.298 -6.325 3.448 ;
      RECT -6.41 3.306 -6.385 3.468 ;
      RECT -6.42 3.31 -6.41 3.48 ;
      RECT -6.425 3.311 -6.42 3.485 ;
      RECT -6.44 3.313 -6.425 3.488 ;
      RECT -6.455 3.315 -6.44 3.493 ;
      RECT -6.46 3.315 -6.455 3.496 ;
      RECT -6.505 3.32 -6.46 3.507 ;
      RECT -6.51 3.324 -6.505 3.519 ;
      RECT -6.535 3.32 -6.51 3.523 ;
      RECT -6.545 3.316 -6.535 3.527 ;
      RECT -6.555 3.315 -6.545 3.531 ;
      RECT -6.57 3.305 -6.555 3.537 ;
      RECT -6.575 3.293 -6.57 3.541 ;
      RECT -6.58 3.29 -6.575 3.542 ;
      RECT -6.585 3.287 -6.58 3.544 ;
      RECT -6.6 3.275 -6.585 3.543 ;
      RECT -6.615 3.257 -6.6 3.54 ;
      RECT -6.635 3.236 -6.615 3.533 ;
      RECT -6.7 3.225 -6.635 3.505 ;
      RECT -6.704 3.225 -6.7 3.484 ;
      RECT -6.79 3.225 -6.704 3.454 ;
      RECT -6.805 3.225 -6.79 3.41 ;
      RECT -6.23 2.325 -6.225 2.56 ;
      RECT -7.1 2.241 -7.095 2.445 ;
      RECT -6.52 2.27 -6.515 2.425 ;
      RECT -6.6 2.25 -6.595 2.425 ;
      RECT -5.93 2.392 -5.915 2.745 ;
      RECT -6.004 2.377 -5.93 2.745 ;
      RECT -6.09 2.36 -6.004 2.745 ;
      RECT -6.1 2.35 -6.09 2.743 ;
      RECT -6.105 2.348 -6.1 2.738 ;
      RECT -6.12 2.346 -6.105 2.724 ;
      RECT -6.19 2.338 -6.12 2.664 ;
      RECT -6.21 2.329 -6.19 2.598 ;
      RECT -6.215 2.326 -6.21 2.578 ;
      RECT -6.225 2.325 -6.215 2.568 ;
      RECT -6.235 2.325 -6.23 2.552 ;
      RECT -6.245 2.324 -6.235 2.542 ;
      RECT -6.255 2.322 -6.245 2.53 ;
      RECT -6.27 2.319 -6.255 2.51 ;
      RECT -6.28 2.317 -6.27 2.495 ;
      RECT -6.3 2.314 -6.28 2.483 ;
      RECT -6.305 2.312 -6.3 2.473 ;
      RECT -6.33 2.31 -6.305 2.46 ;
      RECT -6.36 2.305 -6.33 2.445 ;
      RECT -6.44 2.296 -6.36 2.436 ;
      RECT -6.485 2.285 -6.44 2.429 ;
      RECT -6.505 2.276 -6.485 2.426 ;
      RECT -6.515 2.271 -6.505 2.425 ;
      RECT -6.56 2.265 -6.52 2.425 ;
      RECT -6.575 2.257 -6.56 2.425 ;
      RECT -6.595 2.252 -6.575 2.425 ;
      RECT -6.615 2.249 -6.6 2.425 ;
      RECT -6.698 2.248 -6.615 2.424 ;
      RECT -6.784 2.247 -6.698 2.42 ;
      RECT -6.87 2.245 -6.784 2.417 ;
      RECT -6.923 2.244 -6.87 2.419 ;
      RECT -7.009 2.243 -6.923 2.428 ;
      RECT -7.095 2.242 -7.009 2.44 ;
      RECT -7.115 2.241 -7.1 2.448 ;
      RECT -7.195 2.24 -7.115 2.46 ;
      RECT -7.22 2.24 -7.195 2.473 ;
      RECT -7.245 2.24 -7.22 2.488 ;
      RECT -7.25 2.24 -7.245 2.51 ;
      RECT -7.255 2.24 -7.25 2.528 ;
      RECT -7.26 2.24 -7.255 2.545 ;
      RECT -7.265 2.24 -7.26 2.558 ;
      RECT -7.27 2.24 -7.265 2.568 ;
      RECT -7.31 2.24 -7.27 2.653 ;
      RECT -7.325 2.24 -7.31 2.738 ;
      RECT -7.335 2.241 -7.325 2.75 ;
      RECT -7.37 2.246 -7.335 2.755 ;
      RECT -7.41 2.255 -7.37 2.755 ;
      RECT -7.425 2.265 -7.41 2.755 ;
      RECT -7.43 2.275 -7.425 2.755 ;
      RECT -7.45 2.302 -7.43 2.755 ;
      RECT -7.5 2.385 -7.45 2.755 ;
      RECT -7.505 2.447 -7.5 2.755 ;
      RECT -7.515 2.46 -7.505 2.755 ;
      RECT -7.525 2.482 -7.515 2.755 ;
      RECT -7.535 2.507 -7.525 2.75 ;
      RECT -7.54 2.545 -7.535 2.743 ;
      RECT -7.55 2.655 -7.54 2.738 ;
      RECT -6.155 3.576 -6.14 3.835 ;
      RECT -6.155 3.591 -6.135 3.834 ;
      RECT -6.239 3.591 -6.135 3.832 ;
      RECT -6.239 3.605 -6.13 3.831 ;
      RECT -6.325 3.647 -6.125 3.828 ;
      RECT -6.33 3.59 -6.14 3.823 ;
      RECT -6.33 3.661 -6.12 3.82 ;
      RECT -6.335 3.692 -6.12 3.818 ;
      RECT -6.33 3.689 -6.105 3.808 ;
      RECT -6.335 3.735 -6.09 3.793 ;
      RECT -6.335 3.763 -6.085 3.778 ;
      RECT -6.325 3.565 -6.155 3.828 ;
      RECT -6.565 2.575 -6.395 2.745 ;
      RECT -6.6 2.575 -6.395 2.74 ;
      RECT -6.61 2.575 -6.395 2.733 ;
      RECT -6.615 2.56 -6.445 2.73 ;
      RECT -7.785 3.097 -7.52 3.54 ;
      RECT -7.79 3.068 -7.575 3.538 ;
      RECT -7.795 3.222 -7.515 3.533 ;
      RECT -7.79 3.117 -7.515 3.533 ;
      RECT -7.79 3.128 -7.505 3.52 ;
      RECT -7.79 3.075 -7.545 3.538 ;
      RECT -7.785 3.062 -7.575 3.54 ;
      RECT -7.785 3.06 -7.625 3.54 ;
      RECT -7.684 3.052 -7.625 3.54 ;
      RECT -7.77 3.053 -7.625 3.54 ;
      RECT -7.684 3.051 -7.635 3.54 ;
      RECT -7.88 1.866 -7.705 2.165 ;
      RECT -7.83 1.828 -7.705 2.165 ;
      RECT -7.845 1.83 -7.619 2.157 ;
      RECT -7.845 1.833 -7.58 2.144 ;
      RECT -7.845 1.834 -7.57 2.13 ;
      RECT -7.89 1.885 -7.57 2.12 ;
      RECT -7.845 1.835 -7.565 2.115 ;
      RECT -7.89 2.045 -7.56 2.105 ;
      RECT -7.905 1.905 -7.565 2.045 ;
      RECT -7.91 1.921 -7.565 1.985 ;
      RECT -7.865 1.845 -7.565 2.115 ;
      RECT -7.83 1.826 -7.744 2.165 ;
      RECT 5.895 0.575 6.065 1.085 ;
      RECT 5.895 2.395 6.065 3.865 ;
      RECT 5.895 5.015 6.065 6.485 ;
      RECT 5.895 7.795 6.065 8.305 ;
      RECT 4.905 0.575 5.075 1.085 ;
      RECT 4.905 2.395 5.075 3.865 ;
      RECT 4.905 5.015 5.075 6.485 ;
      RECT 4.905 7.795 5.075 8.305 ;
      RECT 3.54 0.575 3.71 3.865 ;
      RECT 3.54 5.015 3.71 8.305 ;
      RECT 3.11 0.575 3.28 1.085 ;
      RECT 3.11 1.655 3.28 3.865 ;
      RECT 3.11 5.015 3.28 7.225 ;
      RECT 3.11 7.795 3.28 8.305 ;
      RECT 1.74 1.66 1.91 2.935 ;
      RECT 1.74 5.945 1.91 7.22 ;
  END
END sky130_osu_single_mpr2ya_8

END LIBRARY
