magic
tech sky130A
magscale 1 2
timestamp 1712684334
<< nwell >>
rect 3560 1748 3694 1749
rect 3009 1461 4277 1748
rect 6971 1745 7128 1749
rect 10418 1746 10456 1749
rect 13862 1748 14043 1749
rect 17305 1748 17466 1749
rect 7159 1636 7215 1692
rect 10603 1637 10659 1693
rect 14047 1636 14103 1692
rect 17491 1636 17547 1692
rect 3006 1405 4277 1461
rect 3000 1400 4294 1405
rect 3000 1283 4388 1400
rect 3000 955 4277 1283
rect 5807 1086 7716 1406
rect 9251 1086 11161 1406
rect 12695 1086 14605 1406
rect 16139 1086 18049 1406
rect 19583 1086 20780 1406
rect 6883 986 6941 1044
rect 10327 986 10385 1044
rect 13771 987 13829 1045
rect 17215 986 17273 1044
rect 20659 986 20717 1044
rect 2999 742 4277 955
rect 6970 743 7029 757
rect 13862 750 13906 751
rect 10417 743 10470 750
rect 13860 743 13906 750
rect 13860 742 13904 743
rect 17305 742 17335 745
<< ndiff >>
rect 6894 441 6929 475
rect 10338 441 10373 475
rect 13782 442 13817 476
rect 13786 441 13817 442
rect 17226 441 17261 475
rect 20670 441 20705 475
<< pdiff >>
rect 3045 1647 3079 1681
rect 3728 1646 3762 1680
rect 7172 1646 7206 1680
rect 10616 1646 10650 1680
rect 14060 1646 14094 1680
rect 17504 1646 17538 1680
<< locali >>
rect 9 2172 20783 2492
rect 3406 1405 3440 1470
rect 0 1400 4294 1405
rect 0 1283 4388 1400
rect 0 1085 3879 1283
rect 5807 1086 7716 1406
rect 9251 1086 11161 1406
rect 12695 1086 14605 1406
rect 16139 1086 18049 1406
rect 19583 1086 20780 1406
rect 6968 1085 7007 1086
rect 17301 1085 17347 1086
rect 9 0 20783 320
<< viali >>
rect 3045 1647 3079 1681
rect 6894 441 6929 475
rect 10338 441 10373 475
rect 13782 442 13817 476
rect 17226 441 17261 475
rect 20670 441 20705 475
<< metal1 >>
rect 9 2172 20783 2492
rect 20704 1982 20706 2013
rect 20665 1975 20730 1982
rect 20665 1923 20672 1975
rect 20724 1923 20730 1975
rect 3302 1862 3308 1918
rect 3364 1862 3370 1918
rect 20665 1917 20730 1923
rect 6896 1847 6961 1854
rect 4084 1826 4088 1829
rect 6896 1795 6903 1847
rect 6955 1795 6961 1847
rect 6896 1789 6961 1795
rect 10340 1847 10405 1854
rect 10340 1795 10347 1847
rect 10399 1795 10405 1847
rect 10340 1789 10405 1795
rect 13784 1848 13849 1855
rect 13784 1796 13791 1848
rect 13843 1796 13849 1848
rect 13784 1790 13849 1796
rect 17228 1847 17293 1854
rect 17228 1795 17235 1847
rect 17287 1795 17293 1847
rect 17228 1789 17293 1795
rect 3227 1714 3233 1770
rect 3289 1714 3295 1770
rect 3034 1681 3092 1686
rect 3034 1647 3045 1681
rect 3079 1647 3092 1681
rect 3034 1640 3092 1647
rect 0 1400 4294 1405
rect 0 1283 4388 1400
rect 0 1085 3879 1283
rect 5807 1086 7716 1406
rect 9251 1086 11161 1406
rect 12695 1086 14605 1406
rect 16139 1086 18049 1406
rect 19583 1086 20780 1406
rect 6968 1085 7007 1086
rect 17301 1085 17347 1086
rect 17228 640 17262 674
rect 13783 441 13817 442
rect 9 0 20783 320
<< via1 >>
rect 20672 1923 20724 1975
rect 3308 1862 3364 1918
rect 6903 1795 6955 1847
rect 10347 1795 10399 1847
rect 13791 1796 13843 1848
rect 17235 1795 17287 1847
rect 3233 1714 3289 1770
rect 3715 1636 3771 1692
rect 7159 1636 7215 1692
rect 10603 1637 10659 1693
rect 14047 1636 14103 1692
rect 17491 1636 17547 1692
rect 6883 986 6941 1044
rect 10327 986 10385 1044
rect 13771 987 13829 1045
rect 17215 986 17273 1044
rect 20659 986 20717 1044
<< metal2 >>
rect 3242 2011 20706 2045
rect 3242 1776 3276 2011
rect 20672 1982 20706 2011
rect 20665 1975 20730 1982
rect 3308 1918 3364 1924
rect 20665 1923 20672 1975
rect 20724 1923 20730 1975
rect 20665 1917 20730 1923
rect 3364 1869 3549 1903
rect 3308 1856 3364 1862
rect 3515 1828 3549 1869
rect 6896 1847 6961 1854
rect 3515 1794 4086 1828
rect 6896 1795 6903 1847
rect 6955 1829 6961 1847
rect 10340 1847 10405 1854
rect 6955 1828 7143 1829
rect 6955 1795 7522 1828
rect 6896 1789 6961 1795
rect 7143 1794 7522 1795
rect 10340 1795 10347 1847
rect 10399 1829 10405 1847
rect 13784 1848 13849 1855
rect 10399 1828 10577 1829
rect 10399 1795 11024 1828
rect 10340 1789 10405 1795
rect 10577 1794 11024 1795
rect 13784 1796 13791 1848
rect 13843 1830 13849 1848
rect 17228 1847 17293 1854
rect 13843 1829 13994 1830
rect 13843 1828 14009 1829
rect 13843 1796 14466 1828
rect 13784 1790 13849 1796
rect 13994 1795 14466 1796
rect 14009 1794 14466 1795
rect 17228 1795 17235 1847
rect 17287 1829 17293 1847
rect 17287 1828 17385 1829
rect 17287 1795 17910 1828
rect 17228 1789 17293 1795
rect 17385 1794 17910 1795
rect 3233 1770 3289 1776
rect 3233 1708 3289 1714
<< via2 >>
rect 3715 1636 3771 1692
rect 7159 1636 7215 1692
rect 10603 1637 10659 1693
rect 14047 1636 14103 1692
rect 17491 1636 17547 1692
rect 6883 986 6941 1044
rect 10327 986 10385 1044
rect 13771 987 13829 1045
rect 17215 986 17273 1044
rect 20659 986 20717 1044
<< metal3 >>
rect 3709 1692 3776 2477
rect 7153 1692 7220 2477
rect 10597 1693 10664 2478
rect 14041 1692 14108 2477
rect 17485 1692 17552 2477
rect 6874 0 6950 986
rect 10318 0 10394 986
rect 13762 1 13838 987
rect 17206 0 17282 986
rect 20650 0 20726 986
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1710278372
transform 1 0 3009 0 -1 2233
box -10 0 552 902
use sky130_osu_single_mpr2ct_8_b0r2  sky130_osu_single_mpr2ct_8_b0r2_0
timestamp 1712684334
transform 1 0 17334 0 1 0
box 0 0 3449 2492
use sky130_osu_single_mpr2ct_8_b0r2  sky130_osu_single_mpr2ct_8_b0r2_1
timestamp 1712684334
transform 1 0 3558 0 1 0
box 0 0 3449 2492
use sky130_osu_single_mpr2ct_8_b0r2  sky130_osu_single_mpr2ct_8_b0r2_2
timestamp 1712684334
transform 1 0 7002 0 1 0
box 0 0 3449 2492
use sky130_osu_single_mpr2ct_8_b0r2  sky130_osu_single_mpr2ct_8_b0r2_3
timestamp 1712684334
transform 1 0 10446 0 1 1
box 0 0 3449 2492
use sky130_osu_single_mpr2ct_8_b0r2  sky130_osu_single_mpr2ct_8_b0r2_4
timestamp 1712684334
transform 1 0 13890 0 1 0
box 0 0 3449 2492
<< labels >>
flabel metal1 s 3034 1640 3092 1686 0 FreeSans 100 0 0 0 start
port 15 nsew signal input
flabel metal1 s 6894 441 6929 475 0 FreeSans 100 0 0 0 X1_Y1
port 10 s signal output
flabel metal1 s 17225 441 17261 475 0 FreeSans 100 0 0 0 X4_Y1
port 19 nsew signal output
flabel metal1 s 20670 441 20705 475 0 FreeSans 100 0 0 0 X5_Y1
port 6 s signal output
flabel metal1 s 5807 1086 7716 1406 0 FreeSans 100 0 0 0 vccd1
port 17 nsew power bidirectional
flabel metal1 s 9251 1086 11161 1406 0 FreeSans 100 0 0 0 vccd1
port 17 nsew power bidirectional
flabel metal1 s 12695 1086 14605 1406 0 FreeSans 100 0 0 0 vccd1
port 17 nsew power bidirectional
flabel metal1 s 16139 1086 18049 1406 0 FreeSans 100 0 0 0 vccd1
port 17 nsew power bidirectional
flabel metal1 s 19583 1086 20780 1406 0 FreeSans 100 0 0 0 vccd1
port 17 nsew power bidirectional
flabel metal1 s 9 2172 20783 2492 0 FreeSans 100 0 0 0 vssd1
port 18 nsew ground bidirectional
flabel metal1 s 0 1085 3879 1405 0 FreeSans 100 0 0 0 vccd1
port 17 nsew power bidirectional
flabel metal1 s 9 0 20783 320 0 FreeSans 100 0 0 0 vssd1
port 18 nsew ground bidirectional
flabel metal1 s 3727 1647 3761 1681 0 FreeSans 100 0 0 0 s1
port 1 n signal input
flabel metal1 s 7171 1647 7205 1681 0 FreeSans 100 0 0 0 s2
port 2 n signal input
flabel metal1 s 10615 1647 10649 1681 0 FreeSans 100 0 0 0 s3
port 3 n signal input
flabel metal1 s 14059 1647 14093 1681 0 FreeSans 100 0 0 0 s4
port 14 n signal input
flabel metal1 s 17503 1647 17537 1681 0 FreeSans 100 0 0 0 s5
port 13 n signal input
flabel metal1 s 13782 442 13817 476 0 FreeSans 100 0 0 0 X3_Y1
port 8 s signal output
flabel metal1 s 10338 441 10373 475 0 FreeSans 100 0 0 0 X2_Y1
port 9 s signal output
<< end >>
