VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_osu_ring_oscillator_mpr2aa_8_b0r1
  CLASS CORE ;
  ORIGIN 4.14 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2aa_8_b0r1 -4.14 0 ;
  SIZE 142.495 BY 3.2 ;
  SYMMETRY X Y ;
  SITE b0r1_b0r2_HFix ;
  OBS
    LAYER met4 ;
      RECT 134.775 0.84 135.105 1.175 ;
      RECT -2.005 0.07 -1.675 0.945 ;
      RECT 134.775 0.07 135.1 1.175 ;
      RECT -2.005 0.07 135.1 0.39 ;
      RECT 126.83 1.65 132.075 1.98 ;
      RECT 113.8 1.645 114.14 1.98 ;
      RECT 113.8 1.655 132.075 1.975 ;
      RECT 130.765 0.695 131.22 1.18 ;
      RECT 130.76 0.695 131.22 1.125 ;
      RECT 126.215 0.69 126.755 1.1 ;
      RECT 112.955 0.71 113.285 1.04 ;
      RECT 112.955 0.715 113.48 1.035 ;
      RECT 112.955 0.715 131.22 1.015 ;
      RECT 113.67 0.695 131.22 1.015 ;
      RECT 126.045 0.69 127.085 1.015 ;
      RECT 99.235 1.65 104.48 1.98 ;
      RECT 86.205 1.645 86.545 1.98 ;
      RECT 86.205 1.655 104.48 1.975 ;
      RECT 103.17 0.695 103.625 1.18 ;
      RECT 103.165 0.695 103.625 1.125 ;
      RECT 98.62 0.69 99.16 1.1 ;
      RECT 85.36 0.71 85.69 1.04 ;
      RECT 85.36 0.715 85.885 1.035 ;
      RECT 85.36 0.715 103.625 1.015 ;
      RECT 86.075 0.695 103.625 1.015 ;
      RECT 98.45 0.69 99.49 1.015 ;
      RECT 71.64 1.65 76.885 1.98 ;
      RECT 58.61 1.645 58.95 1.98 ;
      RECT 58.61 1.655 76.885 1.975 ;
      RECT 75.575 0.695 76.03 1.18 ;
      RECT 75.57 0.695 76.03 1.125 ;
      RECT 71.025 0.69 71.565 1.1 ;
      RECT 57.765 0.71 58.095 1.04 ;
      RECT 57.765 0.715 58.29 1.035 ;
      RECT 57.765 0.715 76.03 1.015 ;
      RECT 58.48 0.695 76.03 1.015 ;
      RECT 70.855 0.69 71.895 1.015 ;
      RECT 44.045 1.65 49.29 1.98 ;
      RECT 31.015 1.645 31.355 1.98 ;
      RECT 31.015 1.655 49.29 1.975 ;
      RECT 47.98 0.695 48.435 1.18 ;
      RECT 47.975 0.695 48.435 1.125 ;
      RECT 43.43 0.69 43.97 1.1 ;
      RECT 30.17 0.71 30.5 1.04 ;
      RECT 30.17 0.715 30.695 1.035 ;
      RECT 30.17 0.715 48.435 1.015 ;
      RECT 30.885 0.695 48.435 1.015 ;
      RECT 43.26 0.69 44.3 1.015 ;
      RECT 16.45 1.65 21.695 1.98 ;
      RECT 3.42 1.645 3.76 1.98 ;
      RECT 3.42 1.655 21.695 1.975 ;
      RECT 20.385 0.695 20.84 1.18 ;
      RECT 20.38 0.695 20.84 1.125 ;
      RECT 15.835 0.69 16.375 1.1 ;
      RECT 2.575 0.71 2.905 1.04 ;
      RECT 2.575 0.715 3.1 1.035 ;
      RECT 2.575 0.715 20.84 1.015 ;
      RECT 3.29 0.695 20.84 1.015 ;
      RECT 15.665 0.69 16.705 1.015 ;
      RECT 116.4 2.38 126.245 2.715 ;
      RECT 88.805 2.38 98.65 2.715 ;
      RECT 61.21 2.38 71.055 2.715 ;
      RECT 33.615 2.38 43.46 2.715 ;
      RECT 6.02 2.38 15.865 2.715 ;
    LAYER via3 ;
      RECT 134.84 0.905 135.04 1.105 ;
      RECT 131.81 1.715 132.01 1.915 ;
      RECT 130.955 0.845 131.155 1.045 ;
      RECT 127.675 1.715 127.875 1.915 ;
      RECT 126.415 0.785 126.615 0.985 ;
      RECT 125.97 2.445 126.17 2.645 ;
      RECT 116.465 2.445 116.665 2.645 ;
      RECT 113.875 1.715 114.075 1.915 ;
      RECT 113.02 0.775 113.22 0.975 ;
      RECT 104.215 1.715 104.415 1.915 ;
      RECT 103.36 0.845 103.56 1.045 ;
      RECT 100.08 1.715 100.28 1.915 ;
      RECT 98.82 0.785 99.02 0.985 ;
      RECT 98.375 2.445 98.575 2.645 ;
      RECT 88.87 2.445 89.07 2.645 ;
      RECT 86.28 1.715 86.48 1.915 ;
      RECT 85.425 0.775 85.625 0.975 ;
      RECT 76.62 1.715 76.82 1.915 ;
      RECT 75.765 0.845 75.965 1.045 ;
      RECT 72.485 1.715 72.685 1.915 ;
      RECT 71.225 0.785 71.425 0.985 ;
      RECT 70.78 2.445 70.98 2.645 ;
      RECT 61.275 2.445 61.475 2.645 ;
      RECT 58.685 1.715 58.885 1.915 ;
      RECT 57.83 0.775 58.03 0.975 ;
      RECT 49.025 1.715 49.225 1.915 ;
      RECT 48.17 0.845 48.37 1.045 ;
      RECT 44.89 1.715 45.09 1.915 ;
      RECT 43.63 0.785 43.83 0.985 ;
      RECT 43.185 2.445 43.385 2.645 ;
      RECT 33.68 2.445 33.88 2.645 ;
      RECT 31.09 1.715 31.29 1.915 ;
      RECT 30.235 0.775 30.435 0.975 ;
      RECT 21.43 1.715 21.63 1.915 ;
      RECT 20.575 0.845 20.775 1.045 ;
      RECT 17.295 1.715 17.495 1.915 ;
      RECT 16.035 0.785 16.235 0.985 ;
      RECT 15.59 2.445 15.79 2.645 ;
      RECT 6.085 2.445 6.285 2.645 ;
      RECT 3.495 1.715 3.695 1.915 ;
      RECT 2.64 0.775 2.84 0.975 ;
      RECT -1.94 0.68 -1.74 0.88 ;
    LAYER met3 ;
      RECT 125.89 2.38 126.23 2.735 ;
      RECT 129.91 0.59 130.28 2.71 ;
      RECT 125.895 2.34 130.28 2.71 ;
      RECT 125.895 1.4 126.245 2.71 ;
      RECT 125.895 1.4 126.265 1.77 ;
      RECT 123.6 1.715 123.93 2.445 ;
      RECT 123.6 1.715 124.56 2.045 ;
      RECT 124.23 0.06 124.56 2.045 ;
      RECT 124.21 0.06 124.58 0.43 ;
      RECT 110.53 1.71 110.995 2.08 ;
      RECT 110.66 0.07 110.995 2.08 ;
      RECT 119.96 0.755 120.29 1.485 ;
      RECT 119.08 0.07 119.41 1.485 ;
      RECT 123.12 0.59 123.45 1.32 ;
      RECT 123.08 0.475 123.26 1.125 ;
      RECT 119.08 0.755 123.45 1.09 ;
      RECT 119.08 0.15 119.415 1.09 ;
      RECT 119.075 0.15 119.415 0.485 ;
      RECT 110.66 0.07 111.165 0.485 ;
      RECT 110.66 0.07 119.41 0.37 ;
      RECT 119.58 2.275 119.91 2.605 ;
      RECT 118.375 2.29 119.91 2.59 ;
      RECT 118.375 1.17 118.675 2.59 ;
      RECT 118.12 1.155 118.45 1.485 ;
      RECT 116.405 0.595 116.725 2.735 ;
      RECT 116.4 0.595 116.73 2.72 ;
      RECT 98.295 2.38 98.635 2.735 ;
      RECT 102.315 0.59 102.685 2.71 ;
      RECT 98.3 2.34 102.685 2.71 ;
      RECT 98.3 1.4 98.65 2.71 ;
      RECT 98.3 1.4 98.67 1.77 ;
      RECT 96.005 1.715 96.335 2.445 ;
      RECT 96.005 1.715 96.965 2.045 ;
      RECT 96.635 0.06 96.965 2.045 ;
      RECT 96.615 0.06 96.985 0.43 ;
      RECT 82.935 1.71 83.4 2.08 ;
      RECT 83.065 0.07 83.4 2.08 ;
      RECT 92.365 0.755 92.695 1.485 ;
      RECT 91.485 0.07 91.815 1.485 ;
      RECT 95.525 0.59 95.855 1.32 ;
      RECT 95.485 0.475 95.665 1.125 ;
      RECT 91.485 0.755 95.855 1.09 ;
      RECT 91.485 0.15 91.82 1.09 ;
      RECT 91.48 0.15 91.82 0.485 ;
      RECT 83.065 0.07 83.57 0.485 ;
      RECT 83.065 0.07 91.815 0.37 ;
      RECT 91.985 2.275 92.315 2.605 ;
      RECT 90.78 2.29 92.315 2.59 ;
      RECT 90.78 1.17 91.08 2.59 ;
      RECT 90.525 1.155 90.855 1.485 ;
      RECT 88.81 0.595 89.13 2.735 ;
      RECT 88.805 0.595 89.135 2.72 ;
      RECT 70.7 2.38 71.04 2.735 ;
      RECT 74.72 0.59 75.09 2.71 ;
      RECT 70.705 2.34 75.09 2.71 ;
      RECT 70.705 1.4 71.055 2.71 ;
      RECT 70.705 1.4 71.075 1.77 ;
      RECT 68.41 1.715 68.74 2.445 ;
      RECT 68.41 1.715 69.37 2.045 ;
      RECT 69.04 0.06 69.37 2.045 ;
      RECT 69.02 0.06 69.39 0.43 ;
      RECT 55.34 1.71 55.805 2.08 ;
      RECT 55.47 0.07 55.805 2.08 ;
      RECT 64.77 0.755 65.1 1.485 ;
      RECT 63.89 0.07 64.22 1.485 ;
      RECT 67.93 0.59 68.26 1.32 ;
      RECT 67.89 0.475 68.07 1.125 ;
      RECT 63.89 0.755 68.26 1.09 ;
      RECT 63.89 0.15 64.225 1.09 ;
      RECT 63.885 0.15 64.225 0.485 ;
      RECT 55.47 0.07 55.975 0.485 ;
      RECT 55.47 0.07 64.22 0.37 ;
      RECT 64.39 2.275 64.72 2.605 ;
      RECT 63.185 2.29 64.72 2.59 ;
      RECT 63.185 1.17 63.485 2.59 ;
      RECT 62.93 1.155 63.26 1.485 ;
      RECT 61.215 0.595 61.535 2.735 ;
      RECT 61.21 0.595 61.54 2.72 ;
      RECT 43.105 2.38 43.445 2.735 ;
      RECT 47.125 0.59 47.495 2.71 ;
      RECT 43.11 2.34 47.495 2.71 ;
      RECT 43.11 1.4 43.46 2.71 ;
      RECT 43.11 1.4 43.48 1.77 ;
      RECT 40.815 1.715 41.145 2.445 ;
      RECT 40.815 1.715 41.775 2.045 ;
      RECT 41.445 0.06 41.775 2.045 ;
      RECT 41.425 0.06 41.795 0.43 ;
      RECT 27.745 1.71 28.21 2.08 ;
      RECT 27.875 0.07 28.21 2.08 ;
      RECT 37.175 0.755 37.505 1.485 ;
      RECT 36.295 0.07 36.625 1.485 ;
      RECT 40.335 0.59 40.665 1.32 ;
      RECT 40.295 0.475 40.475 1.125 ;
      RECT 36.295 0.755 40.665 1.09 ;
      RECT 36.295 0.15 36.63 1.09 ;
      RECT 36.29 0.15 36.63 0.485 ;
      RECT 27.875 0.07 28.38 0.485 ;
      RECT 27.875 0.07 36.625 0.37 ;
      RECT 36.795 2.275 37.125 2.605 ;
      RECT 35.59 2.29 37.125 2.59 ;
      RECT 35.59 1.17 35.89 2.59 ;
      RECT 35.335 1.155 35.665 1.485 ;
      RECT 33.62 0.595 33.94 2.735 ;
      RECT 33.615 0.595 33.945 2.72 ;
      RECT 15.51 2.38 15.85 2.735 ;
      RECT 19.53 0.59 19.9 2.71 ;
      RECT 15.515 2.34 19.9 2.71 ;
      RECT 15.515 1.4 15.865 2.71 ;
      RECT 15.515 1.4 15.885 1.77 ;
      RECT 13.22 1.715 13.55 2.445 ;
      RECT 13.22 1.715 14.18 2.045 ;
      RECT 13.85 0.06 14.18 2.045 ;
      RECT 13.83 0.06 14.2 0.43 ;
      RECT 0.15 1.71 0.615 2.08 ;
      RECT 0.28 0.07 0.615 2.08 ;
      RECT 9.58 0.755 9.91 1.485 ;
      RECT 8.7 0.07 9.03 1.485 ;
      RECT 12.74 0.59 13.07 1.32 ;
      RECT 12.7 0.475 12.88 1.125 ;
      RECT 8.7 0.755 13.07 1.09 ;
      RECT 8.7 0.15 9.035 1.09 ;
      RECT 8.695 0.15 9.035 0.485 ;
      RECT 0.28 0.07 0.785 0.485 ;
      RECT 0.28 0.07 9.03 0.37 ;
      RECT 9.2 2.275 9.53 2.605 ;
      RECT 7.995 2.29 9.53 2.59 ;
      RECT 7.995 1.17 8.295 2.59 ;
      RECT 7.74 1.155 8.07 1.485 ;
      RECT 6.025 0.595 6.345 2.735 ;
      RECT 6.02 0.595 6.35 2.72 ;
      RECT 134.735 0.8 135.105 1.515 ;
      RECT 131.61 1.575 132.15 2.045 ;
      RECT 130.765 0.695 131.305 1.16 ;
      RECT 127.475 1.575 128.015 2.04 ;
      RECT 126.215 0.635 126.755 1.1 ;
      RECT 121.52 1.315 121.85 2.045 ;
      RECT 117.4 1.155 117.73 1.885 ;
      RECT 114.96 1.315 115.29 2.045 ;
      RECT 113.615 1.57 114.155 2.035 ;
      RECT 112.47 0.69 113.67 1.095 ;
      RECT 104.015 1.575 104.555 2.045 ;
      RECT 103.17 0.695 103.71 1.16 ;
      RECT 99.88 1.575 100.42 2.04 ;
      RECT 98.62 0.635 99.16 1.1 ;
      RECT 93.925 1.315 94.255 2.045 ;
      RECT 89.805 1.155 90.135 1.885 ;
      RECT 87.365 1.315 87.695 2.045 ;
      RECT 86.02 1.57 86.56 2.035 ;
      RECT 84.875 0.69 86.075 1.095 ;
      RECT 76.42 1.575 76.96 2.045 ;
      RECT 75.575 0.695 76.115 1.16 ;
      RECT 72.285 1.575 72.825 2.04 ;
      RECT 71.025 0.635 71.565 1.1 ;
      RECT 66.33 1.315 66.66 2.045 ;
      RECT 62.21 1.155 62.54 1.885 ;
      RECT 59.77 1.315 60.1 2.045 ;
      RECT 58.425 1.57 58.965 2.035 ;
      RECT 57.28 0.69 58.48 1.095 ;
      RECT 48.825 1.575 49.365 2.045 ;
      RECT 47.98 0.695 48.52 1.16 ;
      RECT 44.69 1.575 45.23 2.04 ;
      RECT 43.43 0.635 43.97 1.1 ;
      RECT 38.735 1.315 39.065 2.045 ;
      RECT 34.615 1.155 34.945 1.885 ;
      RECT 32.175 1.315 32.505 2.045 ;
      RECT 30.83 1.57 31.37 2.035 ;
      RECT 29.685 0.69 30.885 1.095 ;
      RECT 21.23 1.575 21.77 2.045 ;
      RECT 20.385 0.695 20.925 1.16 ;
      RECT 17.095 1.575 17.635 2.04 ;
      RECT 15.835 0.635 16.375 1.1 ;
      RECT 11.14 1.315 11.47 2.045 ;
      RECT 7.02 1.155 7.35 1.885 ;
      RECT 4.58 1.315 4.91 2.045 ;
      RECT 3.235 1.57 3.775 2.035 ;
      RECT 2.09 0.69 3.29 1.095 ;
      RECT -2.075 0.53 -1.59 1.04 ;
    LAYER via2 ;
      RECT 134.82 0.885 135.02 1.085 ;
      RECT 131.79 1.695 131.99 1.895 ;
      RECT 130.935 0.825 131.135 1.025 ;
      RECT 129.995 0.675 130.195 0.875 ;
      RECT 127.655 1.695 127.855 1.895 ;
      RECT 126.395 0.765 126.595 0.965 ;
      RECT 125.98 1.485 126.18 1.685 ;
      RECT 124.295 0.145 124.495 0.345 ;
      RECT 123.665 1.78 123.865 1.98 ;
      RECT 123.185 1.055 123.385 1.255 ;
      RECT 121.585 1.78 121.785 1.98 ;
      RECT 120.025 1.22 120.225 1.42 ;
      RECT 119.645 2.34 119.845 2.54 ;
      RECT 119.145 1.22 119.345 1.42 ;
      RECT 118.185 1.22 118.385 1.42 ;
      RECT 117.465 1.22 117.665 1.42 ;
      RECT 116.465 0.66 116.665 0.86 ;
      RECT 115.025 1.78 115.225 1.98 ;
      RECT 113.855 1.695 114.055 1.895 ;
      RECT 113 0.755 113.2 0.955 ;
      RECT 110.615 1.795 110.815 1.995 ;
      RECT 104.195 1.695 104.395 1.895 ;
      RECT 103.34 0.825 103.54 1.025 ;
      RECT 102.4 0.675 102.6 0.875 ;
      RECT 100.06 1.695 100.26 1.895 ;
      RECT 98.8 0.765 99 0.965 ;
      RECT 98.385 1.485 98.585 1.685 ;
      RECT 96.7 0.145 96.9 0.345 ;
      RECT 96.07 1.78 96.27 1.98 ;
      RECT 95.59 1.055 95.79 1.255 ;
      RECT 93.99 1.78 94.19 1.98 ;
      RECT 92.43 1.22 92.63 1.42 ;
      RECT 92.05 2.34 92.25 2.54 ;
      RECT 91.55 1.22 91.75 1.42 ;
      RECT 90.59 1.22 90.79 1.42 ;
      RECT 89.87 1.22 90.07 1.42 ;
      RECT 88.87 0.66 89.07 0.86 ;
      RECT 87.43 1.78 87.63 1.98 ;
      RECT 86.26 1.695 86.46 1.895 ;
      RECT 85.405 0.755 85.605 0.955 ;
      RECT 83.02 1.795 83.22 1.995 ;
      RECT 76.6 1.695 76.8 1.895 ;
      RECT 75.745 0.825 75.945 1.025 ;
      RECT 74.805 0.675 75.005 0.875 ;
      RECT 72.465 1.695 72.665 1.895 ;
      RECT 71.205 0.765 71.405 0.965 ;
      RECT 70.79 1.485 70.99 1.685 ;
      RECT 69.105 0.145 69.305 0.345 ;
      RECT 68.475 1.78 68.675 1.98 ;
      RECT 67.995 1.055 68.195 1.255 ;
      RECT 66.395 1.78 66.595 1.98 ;
      RECT 64.835 1.22 65.035 1.42 ;
      RECT 64.455 2.34 64.655 2.54 ;
      RECT 63.955 1.22 64.155 1.42 ;
      RECT 62.995 1.22 63.195 1.42 ;
      RECT 62.275 1.22 62.475 1.42 ;
      RECT 61.275 0.66 61.475 0.86 ;
      RECT 59.835 1.78 60.035 1.98 ;
      RECT 58.665 1.695 58.865 1.895 ;
      RECT 57.81 0.755 58.01 0.955 ;
      RECT 55.425 1.795 55.625 1.995 ;
      RECT 49.005 1.695 49.205 1.895 ;
      RECT 48.15 0.825 48.35 1.025 ;
      RECT 47.21 0.675 47.41 0.875 ;
      RECT 44.87 1.695 45.07 1.895 ;
      RECT 43.61 0.765 43.81 0.965 ;
      RECT 43.195 1.485 43.395 1.685 ;
      RECT 41.51 0.145 41.71 0.345 ;
      RECT 40.88 1.78 41.08 1.98 ;
      RECT 40.4 1.055 40.6 1.255 ;
      RECT 38.8 1.78 39 1.98 ;
      RECT 37.24 1.22 37.44 1.42 ;
      RECT 36.86 2.34 37.06 2.54 ;
      RECT 36.36 1.22 36.56 1.42 ;
      RECT 35.4 1.22 35.6 1.42 ;
      RECT 34.68 1.22 34.88 1.42 ;
      RECT 33.68 0.66 33.88 0.86 ;
      RECT 32.24 1.78 32.44 1.98 ;
      RECT 31.07 1.695 31.27 1.895 ;
      RECT 30.215 0.755 30.415 0.955 ;
      RECT 27.83 1.795 28.03 1.995 ;
      RECT 21.41 1.695 21.61 1.895 ;
      RECT 20.555 0.825 20.755 1.025 ;
      RECT 19.615 0.675 19.815 0.875 ;
      RECT 17.275 1.695 17.475 1.895 ;
      RECT 16.015 0.765 16.215 0.965 ;
      RECT 15.6 1.485 15.8 1.685 ;
      RECT 13.915 0.145 14.115 0.345 ;
      RECT 13.285 1.78 13.485 1.98 ;
      RECT 12.805 1.055 13.005 1.255 ;
      RECT 11.205 1.78 11.405 1.98 ;
      RECT 9.645 1.22 9.845 1.42 ;
      RECT 9.265 2.34 9.465 2.54 ;
      RECT 8.765 1.22 8.965 1.42 ;
      RECT 7.805 1.22 8.005 1.42 ;
      RECT 7.085 1.22 7.285 1.42 ;
      RECT 6.085 0.66 6.285 0.86 ;
      RECT 4.645 1.78 4.845 1.98 ;
      RECT 3.475 1.695 3.675 1.895 ;
      RECT 2.62 0.755 2.82 0.955 ;
      RECT 0.235 1.795 0.435 1.995 ;
      RECT -1.94 0.68 -1.74 0.88 ;
    LAYER met2 ;
      RECT 129.91 0.59 130.28 0.96 ;
      RECT 130.425 0.605 130.685 0.93 ;
      RECT 129.91 0.635 130.685 0.895 ;
      RECT 120.695 1.195 120.93 1.455 ;
      RECT 123.84 0.975 124.005 1.235 ;
      RECT 123.745 0.965 123.76 1.235 ;
      RECT 122.345 0.535 122.385 0.675 ;
      RECT 123.76 0.97 123.84 1.235 ;
      RECT 123.705 0.965 123.745 1.201 ;
      RECT 123.691 0.965 123.705 1.201 ;
      RECT 123.605 0.97 123.691 1.203 ;
      RECT 123.56 0.977 123.605 1.205 ;
      RECT 123.53 0.977 123.56 1.207 ;
      RECT 123.505 0.972 123.53 1.209 ;
      RECT 123.475 0.968 123.505 1.218 ;
      RECT 123.465 0.965 123.475 1.23 ;
      RECT 123.46 0.965 123.465 1.238 ;
      RECT 123.455 0.965 123.46 1.243 ;
      RECT 123.445 0.964 123.455 1.253 ;
      RECT 123.44 0.963 123.445 1.263 ;
      RECT 123.425 0.962 123.44 1.268 ;
      RECT 123.397 0.959 123.425 1.295 ;
      RECT 123.311 0.951 123.397 1.295 ;
      RECT 123.225 0.94 123.311 1.295 ;
      RECT 123.185 0.925 123.225 1.295 ;
      RECT 123.145 0.899 123.185 1.295 ;
      RECT 123.14 0.881 123.145 1.107 ;
      RECT 123.13 0.877 123.14 1.097 ;
      RECT 123.115 0.867 123.13 1.084 ;
      RECT 123.095 0.851 123.115 1.069 ;
      RECT 123.08 0.836 123.095 1.054 ;
      RECT 123.07 0.825 123.08 1.044 ;
      RECT 123.045 0.809 123.07 1.033 ;
      RECT 123.04 0.796 123.045 1.023 ;
      RECT 123.035 0.792 123.04 1.018 ;
      RECT 122.98 0.778 123.035 0.996 ;
      RECT 122.941 0.759 122.98 0.96 ;
      RECT 122.855 0.733 122.941 0.913 ;
      RECT 122.851 0.715 122.855 0.879 ;
      RECT 122.765 0.696 122.851 0.857 ;
      RECT 122.76 0.678 122.765 0.835 ;
      RECT 122.755 0.676 122.76 0.833 ;
      RECT 122.745 0.675 122.755 0.828 ;
      RECT 122.685 0.662 122.745 0.814 ;
      RECT 122.64 0.64 122.685 0.793 ;
      RECT 122.58 0.617 122.64 0.772 ;
      RECT 122.516 0.592 122.58 0.747 ;
      RECT 122.43 0.562 122.516 0.716 ;
      RECT 122.415 0.542 122.43 0.695 ;
      RECT 122.385 0.537 122.415 0.686 ;
      RECT 122.332 0.535 122.345 0.675 ;
      RECT 122.246 0.535 122.332 0.677 ;
      RECT 122.16 0.535 122.246 0.679 ;
      RECT 122.14 0.535 122.16 0.683 ;
      RECT 122.095 0.537 122.14 0.694 ;
      RECT 122.055 0.547 122.095 0.71 ;
      RECT 122.051 0.556 122.055 0.718 ;
      RECT 121.965 0.576 122.051 0.734 ;
      RECT 121.955 0.595 121.965 0.752 ;
      RECT 121.95 0.597 121.955 0.755 ;
      RECT 121.94 0.601 121.95 0.758 ;
      RECT 121.92 0.606 121.94 0.768 ;
      RECT 121.89 0.616 121.92 0.788 ;
      RECT 121.885 0.623 121.89 0.802 ;
      RECT 121.875 0.627 121.885 0.809 ;
      RECT 121.86 0.635 121.875 0.82 ;
      RECT 121.85 0.645 121.86 0.831 ;
      RECT 121.84 0.652 121.85 0.839 ;
      RECT 121.815 0.665 121.84 0.854 ;
      RECT 121.751 0.701 121.815 0.893 ;
      RECT 121.665 0.764 121.751 0.957 ;
      RECT 121.63 0.815 121.665 1.01 ;
      RECT 121.625 0.832 121.63 1.027 ;
      RECT 121.61 0.841 121.625 1.034 ;
      RECT 121.59 0.856 121.61 1.048 ;
      RECT 121.585 0.867 121.59 1.058 ;
      RECT 121.565 0.88 121.585 1.068 ;
      RECT 121.56 0.89 121.565 1.078 ;
      RECT 121.545 0.895 121.56 1.087 ;
      RECT 121.535 0.905 121.545 1.098 ;
      RECT 121.505 0.922 121.535 1.115 ;
      RECT 121.495 0.94 121.505 1.133 ;
      RECT 121.48 0.951 121.495 1.144 ;
      RECT 121.44 0.975 121.48 1.16 ;
      RECT 121.405 1.009 121.44 1.177 ;
      RECT 121.375 1.032 121.405 1.189 ;
      RECT 121.36 1.042 121.375 1.198 ;
      RECT 121.32 1.052 121.36 1.209 ;
      RECT 121.3 1.063 121.32 1.221 ;
      RECT 121.295 1.067 121.3 1.228 ;
      RECT 121.28 1.071 121.295 1.233 ;
      RECT 121.27 1.076 121.28 1.238 ;
      RECT 121.265 1.079 121.27 1.241 ;
      RECT 121.235 1.085 121.265 1.248 ;
      RECT 121.2 1.095 121.235 1.262 ;
      RECT 121.14 1.11 121.2 1.282 ;
      RECT 121.085 1.13 121.14 1.306 ;
      RECT 121.056 1.145 121.085 1.324 ;
      RECT 120.97 1.165 121.056 1.349 ;
      RECT 120.965 1.18 120.97 1.369 ;
      RECT 120.955 1.183 120.965 1.37 ;
      RECT 120.93 1.19 120.955 1.455 ;
      RECT 123.625 1.683 123.905 2.02 ;
      RECT 123.625 1.693 123.91 1.978 ;
      RECT 123.625 1.702 123.915 1.875 ;
      RECT 123.625 1.717 123.92 1.743 ;
      RECT 123.625 1.545 123.885 2.02 ;
      RECT 121.345 2.425 121.355 2.615 ;
      RECT 119.605 2.3 119.885 2.58 ;
      RECT 122.65 1.24 122.655 1.725 ;
      RECT 122.545 1.24 122.605 1.5 ;
      RECT 122.87 2.21 122.875 2.285 ;
      RECT 122.86 2.077 122.87 2.32 ;
      RECT 122.85 1.912 122.86 2.341 ;
      RECT 122.845 1.782 122.85 2.357 ;
      RECT 122.835 1.672 122.845 2.373 ;
      RECT 122.83 1.571 122.835 2.39 ;
      RECT 122.825 1.553 122.83 2.4 ;
      RECT 122.82 1.535 122.825 2.41 ;
      RECT 122.81 1.51 122.82 2.425 ;
      RECT 122.805 1.49 122.81 2.44 ;
      RECT 122.785 1.24 122.805 2.465 ;
      RECT 122.77 1.24 122.785 2.498 ;
      RECT 122.74 1.24 122.77 2.52 ;
      RECT 122.72 1.24 122.74 2.534 ;
      RECT 122.7 1.24 122.72 2.05 ;
      RECT 122.715 2.117 122.72 2.539 ;
      RECT 122.71 2.147 122.715 2.541 ;
      RECT 122.705 2.16 122.71 2.544 ;
      RECT 122.7 2.17 122.705 2.548 ;
      RECT 122.695 1.24 122.7 1.968 ;
      RECT 122.695 2.18 122.7 2.55 ;
      RECT 122.69 1.24 122.695 1.945 ;
      RECT 122.68 2.202 122.695 2.55 ;
      RECT 122.675 1.24 122.69 1.89 ;
      RECT 122.67 2.227 122.68 2.55 ;
      RECT 122.67 1.24 122.675 1.835 ;
      RECT 122.66 1.24 122.67 1.783 ;
      RECT 122.665 2.24 122.67 2.551 ;
      RECT 122.66 2.252 122.665 2.552 ;
      RECT 122.655 1.24 122.66 1.743 ;
      RECT 122.655 2.265 122.66 2.553 ;
      RECT 122.64 2.28 122.655 2.554 ;
      RECT 122.645 1.24 122.65 1.705 ;
      RECT 122.64 1.24 122.645 1.67 ;
      RECT 122.635 1.24 122.64 1.645 ;
      RECT 122.63 2.307 122.64 2.556 ;
      RECT 122.625 1.24 122.635 1.603 ;
      RECT 122.625 2.325 122.63 2.557 ;
      RECT 122.62 1.24 122.625 1.563 ;
      RECT 122.62 2.332 122.625 2.558 ;
      RECT 122.615 1.24 122.62 1.535 ;
      RECT 122.61 2.35 122.62 2.559 ;
      RECT 122.605 1.24 122.615 1.515 ;
      RECT 122.6 2.37 122.61 2.561 ;
      RECT 122.59 2.387 122.6 2.562 ;
      RECT 122.555 2.41 122.59 2.565 ;
      RECT 122.5 2.428 122.555 2.571 ;
      RECT 122.414 2.436 122.5 2.58 ;
      RECT 122.328 2.447 122.414 2.591 ;
      RECT 122.242 2.457 122.328 2.602 ;
      RECT 122.156 2.467 122.242 2.614 ;
      RECT 122.07 2.477 122.156 2.625 ;
      RECT 122.05 2.483 122.07 2.631 ;
      RECT 121.97 2.485 122.05 2.635 ;
      RECT 121.965 2.484 121.97 2.64 ;
      RECT 121.957 2.483 121.965 2.64 ;
      RECT 121.871 2.479 121.957 2.638 ;
      RECT 121.785 2.471 121.871 2.635 ;
      RECT 121.699 2.462 121.785 2.631 ;
      RECT 121.613 2.454 121.699 2.628 ;
      RECT 121.527 2.446 121.613 2.624 ;
      RECT 121.441 2.437 121.527 2.621 ;
      RECT 121.355 2.429 121.441 2.617 ;
      RECT 121.3 2.422 121.345 2.615 ;
      RECT 121.215 2.415 121.3 2.613 ;
      RECT 121.141 2.407 121.215 2.609 ;
      RECT 121.055 2.399 121.141 2.606 ;
      RECT 121.052 2.395 121.055 2.604 ;
      RECT 120.966 2.391 121.052 2.603 ;
      RECT 120.88 2.383 120.966 2.6 ;
      RECT 120.795 2.378 120.88 2.597 ;
      RECT 120.709 2.375 120.795 2.594 ;
      RECT 120.623 2.373 120.709 2.591 ;
      RECT 120.537 2.37 120.623 2.588 ;
      RECT 120.451 2.367 120.537 2.585 ;
      RECT 120.365 2.364 120.451 2.582 ;
      RECT 120.289 2.362 120.365 2.579 ;
      RECT 120.203 2.359 120.289 2.576 ;
      RECT 120.117 2.356 120.203 2.574 ;
      RECT 120.031 2.354 120.117 2.571 ;
      RECT 119.945 2.351 120.031 2.568 ;
      RECT 119.885 2.342 119.945 2.566 ;
      RECT 122.395 1.96 122.47 2.22 ;
      RECT 122.375 1.94 122.38 2.22 ;
      RECT 121.695 1.725 121.8 2.02 ;
      RECT 116.14 1.7 116.21 1.96 ;
      RECT 122.035 1.575 122.04 1.946 ;
      RECT 122.025 1.63 122.03 1.946 ;
      RECT 122.33 0.8 122.39 1.06 ;
      RECT 122.385 1.955 122.395 2.22 ;
      RECT 122.38 1.945 122.385 2.22 ;
      RECT 122.3 1.892 122.375 2.22 ;
      RECT 122.325 0.8 122.33 1.08 ;
      RECT 122.315 0.8 122.325 1.1 ;
      RECT 122.3 0.8 122.315 1.13 ;
      RECT 122.285 0.8 122.3 1.173 ;
      RECT 122.28 1.835 122.3 2.22 ;
      RECT 122.27 0.8 122.285 1.21 ;
      RECT 122.265 1.815 122.28 2.22 ;
      RECT 122.265 0.8 122.27 1.233 ;
      RECT 122.255 0.8 122.265 1.258 ;
      RECT 122.225 1.782 122.265 2.22 ;
      RECT 122.23 0.8 122.255 1.308 ;
      RECT 122.225 0.8 122.23 1.363 ;
      RECT 122.22 0.8 122.225 1.405 ;
      RECT 122.21 1.745 122.225 2.22 ;
      RECT 122.215 0.8 122.22 1.448 ;
      RECT 122.21 0.8 122.215 1.513 ;
      RECT 122.205 0.8 122.21 1.535 ;
      RECT 122.205 1.733 122.21 2.085 ;
      RECT 122.2 0.8 122.205 1.603 ;
      RECT 122.2 1.725 122.205 2.068 ;
      RECT 122.195 0.8 122.2 1.648 ;
      RECT 122.19 1.707 122.2 2.045 ;
      RECT 122.19 0.8 122.195 1.685 ;
      RECT 122.18 0.8 122.19 2.025 ;
      RECT 122.175 0.8 122.18 2.008 ;
      RECT 122.17 0.8 122.175 1.993 ;
      RECT 122.165 0.8 122.17 1.978 ;
      RECT 122.145 0.8 122.165 1.968 ;
      RECT 122.14 0.8 122.145 1.958 ;
      RECT 122.13 0.8 122.14 1.954 ;
      RECT 122.125 1.077 122.13 1.953 ;
      RECT 122.12 1.1 122.125 1.952 ;
      RECT 122.115 1.13 122.12 1.951 ;
      RECT 122.11 1.157 122.115 1.95 ;
      RECT 122.105 1.185 122.11 1.95 ;
      RECT 122.1 1.212 122.105 1.95 ;
      RECT 122.095 1.232 122.1 1.95 ;
      RECT 122.09 1.26 122.095 1.95 ;
      RECT 122.08 1.302 122.09 1.95 ;
      RECT 122.07 1.347 122.08 1.949 ;
      RECT 122.065 1.4 122.07 1.948 ;
      RECT 122.06 1.432 122.065 1.947 ;
      RECT 122.055 1.452 122.06 1.946 ;
      RECT 122.05 1.49 122.055 1.946 ;
      RECT 122.045 1.512 122.05 1.946 ;
      RECT 122.04 1.537 122.045 1.946 ;
      RECT 122.03 1.602 122.035 1.946 ;
      RECT 122.015 1.662 122.025 1.946 ;
      RECT 122 1.672 122.015 1.946 ;
      RECT 121.98 1.682 122 1.946 ;
      RECT 121.95 1.687 121.98 1.943 ;
      RECT 121.89 1.697 121.95 1.94 ;
      RECT 121.87 1.706 121.89 1.945 ;
      RECT 121.845 1.712 121.87 1.958 ;
      RECT 121.825 1.717 121.845 1.973 ;
      RECT 121.8 1.722 121.825 2.02 ;
      RECT 121.671 1.724 121.695 2.02 ;
      RECT 121.585 1.719 121.671 2.02 ;
      RECT 121.545 1.716 121.585 2.02 ;
      RECT 121.495 1.718 121.545 2 ;
      RECT 121.465 1.722 121.495 2 ;
      RECT 121.386 1.732 121.465 2 ;
      RECT 121.3 1.747 121.386 2.001 ;
      RECT 121.25 1.757 121.3 2.002 ;
      RECT 121.242 1.76 121.25 2.002 ;
      RECT 121.156 1.762 121.242 2.003 ;
      RECT 121.07 1.766 121.156 2.003 ;
      RECT 120.984 1.77 121.07 2.004 ;
      RECT 120.898 1.773 120.984 2.005 ;
      RECT 120.812 1.777 120.898 2.005 ;
      RECT 120.726 1.781 120.812 2.006 ;
      RECT 120.64 1.784 120.726 2.007 ;
      RECT 120.554 1.788 120.64 2.007 ;
      RECT 120.468 1.792 120.554 2.008 ;
      RECT 120.382 1.796 120.468 2.009 ;
      RECT 120.296 1.799 120.382 2.009 ;
      RECT 120.21 1.803 120.296 2.01 ;
      RECT 120.18 1.805 120.21 2.01 ;
      RECT 120.094 1.808 120.18 2.011 ;
      RECT 120.008 1.812 120.094 2.012 ;
      RECT 119.922 1.816 120.008 2.013 ;
      RECT 119.836 1.819 119.922 2.013 ;
      RECT 119.75 1.823 119.836 2.014 ;
      RECT 119.715 1.828 119.75 2.015 ;
      RECT 119.66 1.838 119.715 2.022 ;
      RECT 119.635 1.85 119.66 2.032 ;
      RECT 119.6 1.863 119.635 2.04 ;
      RECT 119.56 1.88 119.6 2.063 ;
      RECT 119.54 1.893 119.56 2.09 ;
      RECT 119.51 1.905 119.54 2.118 ;
      RECT 119.505 1.913 119.51 2.138 ;
      RECT 119.5 1.916 119.505 2.148 ;
      RECT 119.45 1.928 119.5 2.182 ;
      RECT 119.44 1.943 119.45 2.215 ;
      RECT 119.43 1.949 119.44 2.228 ;
      RECT 119.42 1.956 119.43 2.24 ;
      RECT 119.395 1.969 119.42 2.258 ;
      RECT 119.38 1.984 119.395 2.28 ;
      RECT 119.37 1.992 119.38 2.296 ;
      RECT 119.355 2.001 119.37 2.311 ;
      RECT 119.345 2.011 119.355 2.325 ;
      RECT 119.326 2.024 119.345 2.342 ;
      RECT 119.24 2.069 119.326 2.407 ;
      RECT 119.225 2.114 119.24 2.465 ;
      RECT 119.22 2.123 119.225 2.478 ;
      RECT 119.21 2.13 119.22 2.483 ;
      RECT 119.205 2.135 119.21 2.487 ;
      RECT 119.185 2.145 119.205 2.494 ;
      RECT 119.16 2.165 119.185 2.508 ;
      RECT 119.125 2.19 119.16 2.528 ;
      RECT 119.11 2.213 119.125 2.543 ;
      RECT 119.1 2.223 119.11 2.548 ;
      RECT 119.09 2.231 119.1 2.555 ;
      RECT 119.08 2.24 119.09 2.561 ;
      RECT 119.06 2.252 119.08 2.563 ;
      RECT 119.05 2.265 119.06 2.565 ;
      RECT 119.025 2.28 119.05 2.568 ;
      RECT 119.005 2.297 119.025 2.572 ;
      RECT 118.965 2.325 119.005 2.578 ;
      RECT 118.9 2.372 118.965 2.587 ;
      RECT 118.885 2.405 118.9 2.595 ;
      RECT 118.88 2.412 118.885 2.597 ;
      RECT 118.83 2.437 118.88 2.602 ;
      RECT 118.815 2.461 118.83 2.609 ;
      RECT 118.765 2.466 118.815 2.61 ;
      RECT 118.679 2.47 118.765 2.61 ;
      RECT 118.593 2.47 118.679 2.61 ;
      RECT 118.507 2.47 118.593 2.611 ;
      RECT 118.421 2.47 118.507 2.611 ;
      RECT 118.335 2.47 118.421 2.611 ;
      RECT 118.269 2.47 118.335 2.611 ;
      RECT 118.183 2.47 118.269 2.612 ;
      RECT 118.097 2.47 118.183 2.612 ;
      RECT 118.011 2.471 118.097 2.613 ;
      RECT 117.925 2.471 118.011 2.613 ;
      RECT 117.839 2.471 117.925 2.613 ;
      RECT 117.753 2.471 117.839 2.614 ;
      RECT 117.667 2.471 117.753 2.614 ;
      RECT 117.581 2.472 117.667 2.615 ;
      RECT 117.495 2.472 117.581 2.615 ;
      RECT 117.475 2.472 117.495 2.615 ;
      RECT 117.389 2.472 117.475 2.615 ;
      RECT 117.303 2.472 117.389 2.615 ;
      RECT 117.217 2.473 117.303 2.615 ;
      RECT 117.131 2.473 117.217 2.615 ;
      RECT 117.045 2.473 117.131 2.615 ;
      RECT 116.959 2.474 117.045 2.615 ;
      RECT 116.873 2.474 116.959 2.615 ;
      RECT 116.787 2.474 116.873 2.615 ;
      RECT 116.701 2.474 116.787 2.615 ;
      RECT 116.615 2.475 116.701 2.615 ;
      RECT 116.565 2.472 116.615 2.615 ;
      RECT 116.555 2.47 116.565 2.614 ;
      RECT 116.551 2.47 116.555 2.613 ;
      RECT 116.465 2.465 116.551 2.608 ;
      RECT 116.443 2.458 116.465 2.602 ;
      RECT 116.357 2.449 116.443 2.596 ;
      RECT 116.271 2.436 116.357 2.587 ;
      RECT 116.185 2.422 116.271 2.577 ;
      RECT 116.14 2.412 116.185 2.57 ;
      RECT 116.12 1.7 116.14 1.978 ;
      RECT 116.12 2.405 116.14 2.566 ;
      RECT 116.09 1.7 116.12 2 ;
      RECT 116.08 2.372 116.12 2.563 ;
      RECT 116.075 1.7 116.09 2.02 ;
      RECT 116.075 2.337 116.08 2.561 ;
      RECT 116.07 1.7 116.075 2.145 ;
      RECT 116.07 2.297 116.075 2.561 ;
      RECT 116.06 1.7 116.07 2.561 ;
      RECT 115.985 1.7 116.06 2.555 ;
      RECT 115.955 1.7 115.985 2.545 ;
      RECT 115.95 1.7 115.955 2.537 ;
      RECT 115.945 1.742 115.95 2.53 ;
      RECT 115.935 1.811 115.945 2.521 ;
      RECT 115.93 1.881 115.935 2.473 ;
      RECT 115.925 1.945 115.93 2.37 ;
      RECT 115.92 1.98 115.925 2.325 ;
      RECT 115.918 2.017 115.92 2.217 ;
      RECT 115.915 2.025 115.918 2.21 ;
      RECT 115.91 2.09 115.915 2.153 ;
      RECT 119.985 1.18 120.265 1.46 ;
      RECT 119.975 1.18 120.265 1.323 ;
      RECT 119.93 1.045 120.19 1.305 ;
      RECT 119.93 1.16 120.245 1.305 ;
      RECT 119.93 1.13 120.24 1.305 ;
      RECT 119.93 1.117 120.23 1.305 ;
      RECT 119.93 1.107 120.225 1.305 ;
      RECT 115.905 1.09 116.165 1.35 ;
      RECT 119.675 0.64 119.935 0.9 ;
      RECT 119.665 0.665 119.935 0.86 ;
      RECT 119.66 0.665 119.665 0.859 ;
      RECT 119.59 0.66 119.66 0.851 ;
      RECT 119.505 0.647 119.59 0.834 ;
      RECT 119.501 0.639 119.505 0.824 ;
      RECT 119.415 0.632 119.501 0.814 ;
      RECT 119.406 0.624 119.415 0.804 ;
      RECT 119.32 0.617 119.406 0.792 ;
      RECT 119.3 0.608 119.32 0.778 ;
      RECT 119.245 0.603 119.3 0.77 ;
      RECT 119.235 0.597 119.245 0.764 ;
      RECT 119.215 0.595 119.235 0.76 ;
      RECT 119.207 0.594 119.215 0.756 ;
      RECT 119.121 0.586 119.207 0.745 ;
      RECT 119.035 0.572 119.121 0.725 ;
      RECT 118.975 0.56 119.035 0.71 ;
      RECT 118.965 0.555 118.975 0.705 ;
      RECT 118.915 0.555 118.965 0.707 ;
      RECT 118.868 0.557 118.915 0.711 ;
      RECT 118.782 0.564 118.868 0.716 ;
      RECT 118.696 0.572 118.782 0.722 ;
      RECT 118.61 0.581 118.696 0.728 ;
      RECT 118.551 0.587 118.61 0.733 ;
      RECT 118.465 0.592 118.551 0.739 ;
      RECT 118.39 0.597 118.465 0.745 ;
      RECT 118.351 0.599 118.39 0.75 ;
      RECT 118.265 0.596 118.351 0.755 ;
      RECT 118.18 0.594 118.265 0.762 ;
      RECT 118.148 0.593 118.18 0.765 ;
      RECT 118.062 0.592 118.148 0.766 ;
      RECT 117.976 0.591 118.062 0.767 ;
      RECT 117.89 0.59 117.976 0.767 ;
      RECT 117.804 0.589 117.89 0.768 ;
      RECT 117.718 0.588 117.804 0.769 ;
      RECT 117.632 0.587 117.718 0.77 ;
      RECT 117.546 0.586 117.632 0.77 ;
      RECT 117.46 0.585 117.546 0.771 ;
      RECT 117.41 0.585 117.46 0.772 ;
      RECT 117.396 0.586 117.41 0.772 ;
      RECT 117.31 0.593 117.396 0.773 ;
      RECT 117.236 0.604 117.31 0.774 ;
      RECT 117.15 0.613 117.236 0.775 ;
      RECT 117.115 0.62 117.15 0.79 ;
      RECT 117.09 0.623 117.115 0.82 ;
      RECT 117.065 0.632 117.09 0.849 ;
      RECT 117.055 0.643 117.065 0.869 ;
      RECT 117.045 0.651 117.055 0.883 ;
      RECT 117.04 0.657 117.045 0.893 ;
      RECT 117.015 0.674 117.04 0.91 ;
      RECT 117 0.696 117.015 0.938 ;
      RECT 116.97 0.722 117 0.968 ;
      RECT 116.95 0.751 116.97 0.998 ;
      RECT 116.945 0.766 116.95 1.015 ;
      RECT 116.925 0.781 116.945 1.03 ;
      RECT 116.915 0.799 116.925 1.048 ;
      RECT 116.905 0.81 116.915 1.063 ;
      RECT 116.855 0.842 116.905 1.089 ;
      RECT 116.85 0.872 116.855 1.109 ;
      RECT 116.84 0.885 116.85 1.115 ;
      RECT 116.831 0.895 116.84 1.123 ;
      RECT 116.82 0.906 116.831 1.131 ;
      RECT 116.815 0.916 116.82 1.137 ;
      RECT 116.8 0.937 116.815 1.144 ;
      RECT 116.785 0.967 116.8 1.152 ;
      RECT 116.75 0.997 116.785 1.158 ;
      RECT 116.725 1.015 116.75 1.165 ;
      RECT 116.675 1.023 116.725 1.174 ;
      RECT 116.65 1.028 116.675 1.183 ;
      RECT 116.595 1.034 116.65 1.193 ;
      RECT 116.59 1.039 116.595 1.201 ;
      RECT 116.576 1.042 116.59 1.203 ;
      RECT 116.49 1.054 116.576 1.215 ;
      RECT 116.48 1.066 116.49 1.228 ;
      RECT 116.395 1.079 116.48 1.24 ;
      RECT 116.351 1.096 116.395 1.254 ;
      RECT 116.265 1.113 116.351 1.27 ;
      RECT 116.235 1.127 116.265 1.284 ;
      RECT 116.225 1.132 116.235 1.289 ;
      RECT 116.165 1.135 116.225 1.298 ;
      RECT 119.055 1.405 119.315 1.665 ;
      RECT 119.055 1.405 119.335 1.518 ;
      RECT 119.055 1.405 119.36 1.485 ;
      RECT 119.055 1.405 119.365 1.465 ;
      RECT 119.105 1.18 119.385 1.46 ;
      RECT 118.66 1.915 118.92 2.175 ;
      RECT 118.65 1.772 118.845 2.113 ;
      RECT 118.645 1.88 118.86 2.105 ;
      RECT 118.64 1.93 118.92 2.095 ;
      RECT 118.63 2.007 118.92 2.08 ;
      RECT 118.65 1.855 118.86 2.113 ;
      RECT 118.66 1.73 118.845 2.175 ;
      RECT 118.66 1.625 118.825 2.175 ;
      RECT 118.67 1.612 118.825 2.175 ;
      RECT 118.67 1.57 118.815 2.175 ;
      RECT 118.675 1.495 118.815 2.175 ;
      RECT 118.705 1.145 118.815 2.175 ;
      RECT 118.71 0.875 118.835 1.498 ;
      RECT 118.68 1.45 118.835 1.498 ;
      RECT 118.695 1.252 118.815 2.175 ;
      RECT 118.685 1.362 118.835 1.498 ;
      RECT 118.71 0.875 118.85 1.355 ;
      RECT 118.71 0.875 118.87 1.23 ;
      RECT 118.675 0.875 118.935 1.135 ;
      RECT 118.145 1.18 118.425 1.46 ;
      RECT 118.13 1.18 118.425 1.44 ;
      RECT 116.185 2.045 116.445 2.305 ;
      RECT 117.97 1.9 118.23 2.16 ;
      RECT 117.95 1.92 118.23 2.135 ;
      RECT 117.907 1.92 117.95 2.134 ;
      RECT 117.821 1.921 117.907 2.131 ;
      RECT 117.735 1.922 117.821 2.127 ;
      RECT 117.66 1.924 117.735 2.124 ;
      RECT 117.637 1.925 117.66 2.122 ;
      RECT 117.551 1.926 117.637 2.12 ;
      RECT 117.465 1.927 117.551 2.117 ;
      RECT 117.441 1.928 117.465 2.115 ;
      RECT 117.355 1.93 117.441 2.112 ;
      RECT 117.27 1.932 117.355 2.113 ;
      RECT 117.213 1.933 117.27 2.119 ;
      RECT 117.127 1.935 117.213 2.129 ;
      RECT 117.041 1.938 117.127 2.142 ;
      RECT 116.955 1.94 117.041 2.154 ;
      RECT 116.941 1.941 116.955 2.161 ;
      RECT 116.855 1.942 116.941 2.169 ;
      RECT 116.815 1.944 116.855 2.178 ;
      RECT 116.806 1.945 116.815 2.181 ;
      RECT 116.72 1.953 116.806 2.187 ;
      RECT 116.7 1.962 116.72 2.195 ;
      RECT 116.615 1.977 116.7 2.203 ;
      RECT 116.555 2 116.615 2.214 ;
      RECT 116.545 2.012 116.555 2.219 ;
      RECT 116.505 2.022 116.545 2.223 ;
      RECT 116.45 2.039 116.505 2.231 ;
      RECT 116.445 2.049 116.45 2.235 ;
      RECT 117.511 1.18 117.57 1.577 ;
      RECT 117.425 1.18 117.63 1.568 ;
      RECT 117.42 1.21 117.63 1.563 ;
      RECT 117.386 1.21 117.63 1.561 ;
      RECT 117.3 1.21 117.63 1.555 ;
      RECT 117.255 1.21 117.65 1.533 ;
      RECT 117.255 1.21 117.67 1.488 ;
      RECT 117.215 1.21 117.67 1.478 ;
      RECT 117.425 1.18 117.705 1.46 ;
      RECT 117.16 1.18 117.42 1.44 ;
      RECT 116.345 0.66 116.605 0.92 ;
      RECT 116.425 0.62 116.705 0.9 ;
      RECT 114.985 1.74 115.265 2.02 ;
      RECT 114.955 1.702 115.21 2.005 ;
      RECT 114.95 1.703 115.21 2.003 ;
      RECT 114.945 1.704 115.21 1.997 ;
      RECT 114.94 1.707 115.21 1.99 ;
      RECT 114.935 1.74 115.265 1.983 ;
      RECT 114.905 1.71 115.21 1.97 ;
      RECT 114.905 1.737 115.23 1.97 ;
      RECT 114.905 1.727 115.225 1.97 ;
      RECT 114.905 1.712 115.22 1.97 ;
      RECT 114.985 1.699 115.2 2.02 ;
      RECT 115.071 1.697 115.2 2.02 ;
      RECT 115.157 1.695 115.185 2.02 ;
      RECT 102.315 0.59 102.685 0.96 ;
      RECT 102.83 0.605 103.09 0.93 ;
      RECT 102.315 0.635 103.09 0.895 ;
      RECT 93.1 1.195 93.335 1.455 ;
      RECT 96.245 0.975 96.41 1.235 ;
      RECT 96.15 0.965 96.165 1.235 ;
      RECT 94.75 0.535 94.79 0.675 ;
      RECT 96.165 0.97 96.245 1.235 ;
      RECT 96.11 0.965 96.15 1.201 ;
      RECT 96.096 0.965 96.11 1.201 ;
      RECT 96.01 0.97 96.096 1.203 ;
      RECT 95.965 0.977 96.01 1.205 ;
      RECT 95.935 0.977 95.965 1.207 ;
      RECT 95.91 0.972 95.935 1.209 ;
      RECT 95.88 0.968 95.91 1.218 ;
      RECT 95.87 0.965 95.88 1.23 ;
      RECT 95.865 0.965 95.87 1.238 ;
      RECT 95.86 0.965 95.865 1.243 ;
      RECT 95.85 0.964 95.86 1.253 ;
      RECT 95.845 0.963 95.85 1.263 ;
      RECT 95.83 0.962 95.845 1.268 ;
      RECT 95.802 0.959 95.83 1.295 ;
      RECT 95.716 0.951 95.802 1.295 ;
      RECT 95.63 0.94 95.716 1.295 ;
      RECT 95.59 0.925 95.63 1.295 ;
      RECT 95.55 0.899 95.59 1.295 ;
      RECT 95.545 0.881 95.55 1.107 ;
      RECT 95.535 0.877 95.545 1.097 ;
      RECT 95.52 0.867 95.535 1.084 ;
      RECT 95.5 0.851 95.52 1.069 ;
      RECT 95.485 0.836 95.5 1.054 ;
      RECT 95.475 0.825 95.485 1.044 ;
      RECT 95.45 0.809 95.475 1.033 ;
      RECT 95.445 0.796 95.45 1.023 ;
      RECT 95.44 0.792 95.445 1.018 ;
      RECT 95.385 0.778 95.44 0.996 ;
      RECT 95.346 0.759 95.385 0.96 ;
      RECT 95.26 0.733 95.346 0.913 ;
      RECT 95.256 0.715 95.26 0.879 ;
      RECT 95.17 0.696 95.256 0.857 ;
      RECT 95.165 0.678 95.17 0.835 ;
      RECT 95.16 0.676 95.165 0.833 ;
      RECT 95.15 0.675 95.16 0.828 ;
      RECT 95.09 0.662 95.15 0.814 ;
      RECT 95.045 0.64 95.09 0.793 ;
      RECT 94.985 0.617 95.045 0.772 ;
      RECT 94.921 0.592 94.985 0.747 ;
      RECT 94.835 0.562 94.921 0.716 ;
      RECT 94.82 0.542 94.835 0.695 ;
      RECT 94.79 0.537 94.82 0.686 ;
      RECT 94.737 0.535 94.75 0.675 ;
      RECT 94.651 0.535 94.737 0.677 ;
      RECT 94.565 0.535 94.651 0.679 ;
      RECT 94.545 0.535 94.565 0.683 ;
      RECT 94.5 0.537 94.545 0.694 ;
      RECT 94.46 0.547 94.5 0.71 ;
      RECT 94.456 0.556 94.46 0.718 ;
      RECT 94.37 0.576 94.456 0.734 ;
      RECT 94.36 0.595 94.37 0.752 ;
      RECT 94.355 0.597 94.36 0.755 ;
      RECT 94.345 0.601 94.355 0.758 ;
      RECT 94.325 0.606 94.345 0.768 ;
      RECT 94.295 0.616 94.325 0.788 ;
      RECT 94.29 0.623 94.295 0.802 ;
      RECT 94.28 0.627 94.29 0.809 ;
      RECT 94.265 0.635 94.28 0.82 ;
      RECT 94.255 0.645 94.265 0.831 ;
      RECT 94.245 0.652 94.255 0.839 ;
      RECT 94.22 0.665 94.245 0.854 ;
      RECT 94.156 0.701 94.22 0.893 ;
      RECT 94.07 0.764 94.156 0.957 ;
      RECT 94.035 0.815 94.07 1.01 ;
      RECT 94.03 0.832 94.035 1.027 ;
      RECT 94.015 0.841 94.03 1.034 ;
      RECT 93.995 0.856 94.015 1.048 ;
      RECT 93.99 0.867 93.995 1.058 ;
      RECT 93.97 0.88 93.99 1.068 ;
      RECT 93.965 0.89 93.97 1.078 ;
      RECT 93.95 0.895 93.965 1.087 ;
      RECT 93.94 0.905 93.95 1.098 ;
      RECT 93.91 0.922 93.94 1.115 ;
      RECT 93.9 0.94 93.91 1.133 ;
      RECT 93.885 0.951 93.9 1.144 ;
      RECT 93.845 0.975 93.885 1.16 ;
      RECT 93.81 1.009 93.845 1.177 ;
      RECT 93.78 1.032 93.81 1.189 ;
      RECT 93.765 1.042 93.78 1.198 ;
      RECT 93.725 1.052 93.765 1.209 ;
      RECT 93.705 1.063 93.725 1.221 ;
      RECT 93.7 1.067 93.705 1.228 ;
      RECT 93.685 1.071 93.7 1.233 ;
      RECT 93.675 1.076 93.685 1.238 ;
      RECT 93.67 1.079 93.675 1.241 ;
      RECT 93.64 1.085 93.67 1.248 ;
      RECT 93.605 1.095 93.64 1.262 ;
      RECT 93.545 1.11 93.605 1.282 ;
      RECT 93.49 1.13 93.545 1.306 ;
      RECT 93.461 1.145 93.49 1.324 ;
      RECT 93.375 1.165 93.461 1.349 ;
      RECT 93.37 1.18 93.375 1.369 ;
      RECT 93.36 1.183 93.37 1.37 ;
      RECT 93.335 1.19 93.36 1.455 ;
      RECT 96.03 1.683 96.31 2.02 ;
      RECT 96.03 1.693 96.315 1.978 ;
      RECT 96.03 1.702 96.32 1.875 ;
      RECT 96.03 1.717 96.325 1.743 ;
      RECT 96.03 1.545 96.29 2.02 ;
      RECT 93.75 2.425 93.76 2.615 ;
      RECT 92.01 2.3 92.29 2.58 ;
      RECT 95.055 1.24 95.06 1.725 ;
      RECT 94.95 1.24 95.01 1.5 ;
      RECT 95.275 2.21 95.28 2.285 ;
      RECT 95.265 2.077 95.275 2.32 ;
      RECT 95.255 1.912 95.265 2.341 ;
      RECT 95.25 1.782 95.255 2.357 ;
      RECT 95.24 1.672 95.25 2.373 ;
      RECT 95.235 1.571 95.24 2.39 ;
      RECT 95.23 1.553 95.235 2.4 ;
      RECT 95.225 1.535 95.23 2.41 ;
      RECT 95.215 1.51 95.225 2.425 ;
      RECT 95.21 1.49 95.215 2.44 ;
      RECT 95.19 1.24 95.21 2.465 ;
      RECT 95.175 1.24 95.19 2.498 ;
      RECT 95.145 1.24 95.175 2.52 ;
      RECT 95.125 1.24 95.145 2.534 ;
      RECT 95.105 1.24 95.125 2.05 ;
      RECT 95.12 2.117 95.125 2.539 ;
      RECT 95.115 2.147 95.12 2.541 ;
      RECT 95.11 2.16 95.115 2.544 ;
      RECT 95.105 2.17 95.11 2.548 ;
      RECT 95.1 1.24 95.105 1.968 ;
      RECT 95.1 2.18 95.105 2.55 ;
      RECT 95.095 1.24 95.1 1.945 ;
      RECT 95.085 2.202 95.1 2.55 ;
      RECT 95.08 1.24 95.095 1.89 ;
      RECT 95.075 2.227 95.085 2.55 ;
      RECT 95.075 1.24 95.08 1.835 ;
      RECT 95.065 1.24 95.075 1.783 ;
      RECT 95.07 2.24 95.075 2.551 ;
      RECT 95.065 2.252 95.07 2.552 ;
      RECT 95.06 1.24 95.065 1.743 ;
      RECT 95.06 2.265 95.065 2.553 ;
      RECT 95.045 2.28 95.06 2.554 ;
      RECT 95.05 1.24 95.055 1.705 ;
      RECT 95.045 1.24 95.05 1.67 ;
      RECT 95.04 1.24 95.045 1.645 ;
      RECT 95.035 2.307 95.045 2.556 ;
      RECT 95.03 1.24 95.04 1.603 ;
      RECT 95.03 2.325 95.035 2.557 ;
      RECT 95.025 1.24 95.03 1.563 ;
      RECT 95.025 2.332 95.03 2.558 ;
      RECT 95.02 1.24 95.025 1.535 ;
      RECT 95.015 2.35 95.025 2.559 ;
      RECT 95.01 1.24 95.02 1.515 ;
      RECT 95.005 2.37 95.015 2.561 ;
      RECT 94.995 2.387 95.005 2.562 ;
      RECT 94.96 2.41 94.995 2.565 ;
      RECT 94.905 2.428 94.96 2.571 ;
      RECT 94.819 2.436 94.905 2.58 ;
      RECT 94.733 2.447 94.819 2.591 ;
      RECT 94.647 2.457 94.733 2.602 ;
      RECT 94.561 2.467 94.647 2.614 ;
      RECT 94.475 2.477 94.561 2.625 ;
      RECT 94.455 2.483 94.475 2.631 ;
      RECT 94.375 2.485 94.455 2.635 ;
      RECT 94.37 2.484 94.375 2.64 ;
      RECT 94.362 2.483 94.37 2.64 ;
      RECT 94.276 2.479 94.362 2.638 ;
      RECT 94.19 2.471 94.276 2.635 ;
      RECT 94.104 2.462 94.19 2.631 ;
      RECT 94.018 2.454 94.104 2.628 ;
      RECT 93.932 2.446 94.018 2.624 ;
      RECT 93.846 2.437 93.932 2.621 ;
      RECT 93.76 2.429 93.846 2.617 ;
      RECT 93.705 2.422 93.75 2.615 ;
      RECT 93.62 2.415 93.705 2.613 ;
      RECT 93.546 2.407 93.62 2.609 ;
      RECT 93.46 2.399 93.546 2.606 ;
      RECT 93.457 2.395 93.46 2.604 ;
      RECT 93.371 2.391 93.457 2.603 ;
      RECT 93.285 2.383 93.371 2.6 ;
      RECT 93.2 2.378 93.285 2.597 ;
      RECT 93.114 2.375 93.2 2.594 ;
      RECT 93.028 2.373 93.114 2.591 ;
      RECT 92.942 2.37 93.028 2.588 ;
      RECT 92.856 2.367 92.942 2.585 ;
      RECT 92.77 2.364 92.856 2.582 ;
      RECT 92.694 2.362 92.77 2.579 ;
      RECT 92.608 2.359 92.694 2.576 ;
      RECT 92.522 2.356 92.608 2.574 ;
      RECT 92.436 2.354 92.522 2.571 ;
      RECT 92.35 2.351 92.436 2.568 ;
      RECT 92.29 2.342 92.35 2.566 ;
      RECT 94.8 1.96 94.875 2.22 ;
      RECT 94.78 1.94 94.785 2.22 ;
      RECT 94.1 1.725 94.205 2.02 ;
      RECT 88.545 1.7 88.615 1.96 ;
      RECT 94.44 1.575 94.445 1.946 ;
      RECT 94.43 1.63 94.435 1.946 ;
      RECT 94.735 0.8 94.795 1.06 ;
      RECT 94.79 1.955 94.8 2.22 ;
      RECT 94.785 1.945 94.79 2.22 ;
      RECT 94.705 1.892 94.78 2.22 ;
      RECT 94.73 0.8 94.735 1.08 ;
      RECT 94.72 0.8 94.73 1.1 ;
      RECT 94.705 0.8 94.72 1.13 ;
      RECT 94.69 0.8 94.705 1.173 ;
      RECT 94.685 1.835 94.705 2.22 ;
      RECT 94.675 0.8 94.69 1.21 ;
      RECT 94.67 1.815 94.685 2.22 ;
      RECT 94.67 0.8 94.675 1.233 ;
      RECT 94.66 0.8 94.67 1.258 ;
      RECT 94.63 1.782 94.67 2.22 ;
      RECT 94.635 0.8 94.66 1.308 ;
      RECT 94.63 0.8 94.635 1.363 ;
      RECT 94.625 0.8 94.63 1.405 ;
      RECT 94.615 1.745 94.63 2.22 ;
      RECT 94.62 0.8 94.625 1.448 ;
      RECT 94.615 0.8 94.62 1.513 ;
      RECT 94.61 0.8 94.615 1.535 ;
      RECT 94.61 1.733 94.615 2.085 ;
      RECT 94.605 0.8 94.61 1.603 ;
      RECT 94.605 1.725 94.61 2.068 ;
      RECT 94.6 0.8 94.605 1.648 ;
      RECT 94.595 1.707 94.605 2.045 ;
      RECT 94.595 0.8 94.6 1.685 ;
      RECT 94.585 0.8 94.595 2.025 ;
      RECT 94.58 0.8 94.585 2.008 ;
      RECT 94.575 0.8 94.58 1.993 ;
      RECT 94.57 0.8 94.575 1.978 ;
      RECT 94.55 0.8 94.57 1.968 ;
      RECT 94.545 0.8 94.55 1.958 ;
      RECT 94.535 0.8 94.545 1.954 ;
      RECT 94.53 1.077 94.535 1.953 ;
      RECT 94.525 1.1 94.53 1.952 ;
      RECT 94.52 1.13 94.525 1.951 ;
      RECT 94.515 1.157 94.52 1.95 ;
      RECT 94.51 1.185 94.515 1.95 ;
      RECT 94.505 1.212 94.51 1.95 ;
      RECT 94.5 1.232 94.505 1.95 ;
      RECT 94.495 1.26 94.5 1.95 ;
      RECT 94.485 1.302 94.495 1.95 ;
      RECT 94.475 1.347 94.485 1.949 ;
      RECT 94.47 1.4 94.475 1.948 ;
      RECT 94.465 1.432 94.47 1.947 ;
      RECT 94.46 1.452 94.465 1.946 ;
      RECT 94.455 1.49 94.46 1.946 ;
      RECT 94.45 1.512 94.455 1.946 ;
      RECT 94.445 1.537 94.45 1.946 ;
      RECT 94.435 1.602 94.44 1.946 ;
      RECT 94.42 1.662 94.43 1.946 ;
      RECT 94.405 1.672 94.42 1.946 ;
      RECT 94.385 1.682 94.405 1.946 ;
      RECT 94.355 1.687 94.385 1.943 ;
      RECT 94.295 1.697 94.355 1.94 ;
      RECT 94.275 1.706 94.295 1.945 ;
      RECT 94.25 1.712 94.275 1.958 ;
      RECT 94.23 1.717 94.25 1.973 ;
      RECT 94.205 1.722 94.23 2.02 ;
      RECT 94.076 1.724 94.1 2.02 ;
      RECT 93.99 1.719 94.076 2.02 ;
      RECT 93.95 1.716 93.99 2.02 ;
      RECT 93.9 1.718 93.95 2 ;
      RECT 93.87 1.722 93.9 2 ;
      RECT 93.791 1.732 93.87 2 ;
      RECT 93.705 1.747 93.791 2.001 ;
      RECT 93.655 1.757 93.705 2.002 ;
      RECT 93.647 1.76 93.655 2.002 ;
      RECT 93.561 1.762 93.647 2.003 ;
      RECT 93.475 1.766 93.561 2.003 ;
      RECT 93.389 1.77 93.475 2.004 ;
      RECT 93.303 1.773 93.389 2.005 ;
      RECT 93.217 1.777 93.303 2.005 ;
      RECT 93.131 1.781 93.217 2.006 ;
      RECT 93.045 1.784 93.131 2.007 ;
      RECT 92.959 1.788 93.045 2.007 ;
      RECT 92.873 1.792 92.959 2.008 ;
      RECT 92.787 1.796 92.873 2.009 ;
      RECT 92.701 1.799 92.787 2.009 ;
      RECT 92.615 1.803 92.701 2.01 ;
      RECT 92.585 1.805 92.615 2.01 ;
      RECT 92.499 1.808 92.585 2.011 ;
      RECT 92.413 1.812 92.499 2.012 ;
      RECT 92.327 1.816 92.413 2.013 ;
      RECT 92.241 1.819 92.327 2.013 ;
      RECT 92.155 1.823 92.241 2.014 ;
      RECT 92.12 1.828 92.155 2.015 ;
      RECT 92.065 1.838 92.12 2.022 ;
      RECT 92.04 1.85 92.065 2.032 ;
      RECT 92.005 1.863 92.04 2.04 ;
      RECT 91.965 1.88 92.005 2.063 ;
      RECT 91.945 1.893 91.965 2.09 ;
      RECT 91.915 1.905 91.945 2.118 ;
      RECT 91.91 1.913 91.915 2.138 ;
      RECT 91.905 1.916 91.91 2.148 ;
      RECT 91.855 1.928 91.905 2.182 ;
      RECT 91.845 1.943 91.855 2.215 ;
      RECT 91.835 1.949 91.845 2.228 ;
      RECT 91.825 1.956 91.835 2.24 ;
      RECT 91.8 1.969 91.825 2.258 ;
      RECT 91.785 1.984 91.8 2.28 ;
      RECT 91.775 1.992 91.785 2.296 ;
      RECT 91.76 2.001 91.775 2.311 ;
      RECT 91.75 2.011 91.76 2.325 ;
      RECT 91.731 2.024 91.75 2.342 ;
      RECT 91.645 2.069 91.731 2.407 ;
      RECT 91.63 2.114 91.645 2.465 ;
      RECT 91.625 2.123 91.63 2.478 ;
      RECT 91.615 2.13 91.625 2.483 ;
      RECT 91.61 2.135 91.615 2.487 ;
      RECT 91.59 2.145 91.61 2.494 ;
      RECT 91.565 2.165 91.59 2.508 ;
      RECT 91.53 2.19 91.565 2.528 ;
      RECT 91.515 2.213 91.53 2.543 ;
      RECT 91.505 2.223 91.515 2.548 ;
      RECT 91.495 2.231 91.505 2.555 ;
      RECT 91.485 2.24 91.495 2.561 ;
      RECT 91.465 2.252 91.485 2.563 ;
      RECT 91.455 2.265 91.465 2.565 ;
      RECT 91.43 2.28 91.455 2.568 ;
      RECT 91.41 2.297 91.43 2.572 ;
      RECT 91.37 2.325 91.41 2.578 ;
      RECT 91.305 2.372 91.37 2.587 ;
      RECT 91.29 2.405 91.305 2.595 ;
      RECT 91.285 2.412 91.29 2.597 ;
      RECT 91.235 2.437 91.285 2.602 ;
      RECT 91.22 2.461 91.235 2.609 ;
      RECT 91.17 2.466 91.22 2.61 ;
      RECT 91.084 2.47 91.17 2.61 ;
      RECT 90.998 2.47 91.084 2.61 ;
      RECT 90.912 2.47 90.998 2.611 ;
      RECT 90.826 2.47 90.912 2.611 ;
      RECT 90.74 2.47 90.826 2.611 ;
      RECT 90.674 2.47 90.74 2.611 ;
      RECT 90.588 2.47 90.674 2.612 ;
      RECT 90.502 2.47 90.588 2.612 ;
      RECT 90.416 2.471 90.502 2.613 ;
      RECT 90.33 2.471 90.416 2.613 ;
      RECT 90.244 2.471 90.33 2.613 ;
      RECT 90.158 2.471 90.244 2.614 ;
      RECT 90.072 2.471 90.158 2.614 ;
      RECT 89.986 2.472 90.072 2.615 ;
      RECT 89.9 2.472 89.986 2.615 ;
      RECT 89.88 2.472 89.9 2.615 ;
      RECT 89.794 2.472 89.88 2.615 ;
      RECT 89.708 2.472 89.794 2.615 ;
      RECT 89.622 2.473 89.708 2.615 ;
      RECT 89.536 2.473 89.622 2.615 ;
      RECT 89.45 2.473 89.536 2.615 ;
      RECT 89.364 2.474 89.45 2.615 ;
      RECT 89.278 2.474 89.364 2.615 ;
      RECT 89.192 2.474 89.278 2.615 ;
      RECT 89.106 2.474 89.192 2.615 ;
      RECT 89.02 2.475 89.106 2.615 ;
      RECT 88.97 2.472 89.02 2.615 ;
      RECT 88.96 2.47 88.97 2.614 ;
      RECT 88.956 2.47 88.96 2.613 ;
      RECT 88.87 2.465 88.956 2.608 ;
      RECT 88.848 2.458 88.87 2.602 ;
      RECT 88.762 2.449 88.848 2.596 ;
      RECT 88.676 2.436 88.762 2.587 ;
      RECT 88.59 2.422 88.676 2.577 ;
      RECT 88.545 2.412 88.59 2.57 ;
      RECT 88.525 1.7 88.545 1.978 ;
      RECT 88.525 2.405 88.545 2.566 ;
      RECT 88.495 1.7 88.525 2 ;
      RECT 88.485 2.372 88.525 2.563 ;
      RECT 88.48 1.7 88.495 2.02 ;
      RECT 88.48 2.337 88.485 2.561 ;
      RECT 88.475 1.7 88.48 2.145 ;
      RECT 88.475 2.297 88.48 2.561 ;
      RECT 88.465 1.7 88.475 2.561 ;
      RECT 88.39 1.7 88.465 2.555 ;
      RECT 88.36 1.7 88.39 2.545 ;
      RECT 88.355 1.7 88.36 2.537 ;
      RECT 88.35 1.742 88.355 2.53 ;
      RECT 88.34 1.811 88.35 2.521 ;
      RECT 88.335 1.881 88.34 2.473 ;
      RECT 88.33 1.945 88.335 2.37 ;
      RECT 88.325 1.98 88.33 2.325 ;
      RECT 88.323 2.017 88.325 2.217 ;
      RECT 88.32 2.025 88.323 2.21 ;
      RECT 88.315 2.09 88.32 2.153 ;
      RECT 92.39 1.18 92.67 1.46 ;
      RECT 92.38 1.18 92.67 1.323 ;
      RECT 92.335 1.045 92.595 1.305 ;
      RECT 92.335 1.16 92.65 1.305 ;
      RECT 92.335 1.13 92.645 1.305 ;
      RECT 92.335 1.117 92.635 1.305 ;
      RECT 92.335 1.107 92.63 1.305 ;
      RECT 88.31 1.09 88.57 1.35 ;
      RECT 92.08 0.64 92.34 0.9 ;
      RECT 92.07 0.665 92.34 0.86 ;
      RECT 92.065 0.665 92.07 0.859 ;
      RECT 91.995 0.66 92.065 0.851 ;
      RECT 91.91 0.647 91.995 0.834 ;
      RECT 91.906 0.639 91.91 0.824 ;
      RECT 91.82 0.632 91.906 0.814 ;
      RECT 91.811 0.624 91.82 0.804 ;
      RECT 91.725 0.617 91.811 0.792 ;
      RECT 91.705 0.608 91.725 0.778 ;
      RECT 91.65 0.603 91.705 0.77 ;
      RECT 91.64 0.597 91.65 0.764 ;
      RECT 91.62 0.595 91.64 0.76 ;
      RECT 91.612 0.594 91.62 0.756 ;
      RECT 91.526 0.586 91.612 0.745 ;
      RECT 91.44 0.572 91.526 0.725 ;
      RECT 91.38 0.56 91.44 0.71 ;
      RECT 91.37 0.555 91.38 0.705 ;
      RECT 91.32 0.555 91.37 0.707 ;
      RECT 91.273 0.557 91.32 0.711 ;
      RECT 91.187 0.564 91.273 0.716 ;
      RECT 91.101 0.572 91.187 0.722 ;
      RECT 91.015 0.581 91.101 0.728 ;
      RECT 90.956 0.587 91.015 0.733 ;
      RECT 90.87 0.592 90.956 0.739 ;
      RECT 90.795 0.597 90.87 0.745 ;
      RECT 90.756 0.599 90.795 0.75 ;
      RECT 90.67 0.596 90.756 0.755 ;
      RECT 90.585 0.594 90.67 0.762 ;
      RECT 90.553 0.593 90.585 0.765 ;
      RECT 90.467 0.592 90.553 0.766 ;
      RECT 90.381 0.591 90.467 0.767 ;
      RECT 90.295 0.59 90.381 0.767 ;
      RECT 90.209 0.589 90.295 0.768 ;
      RECT 90.123 0.588 90.209 0.769 ;
      RECT 90.037 0.587 90.123 0.77 ;
      RECT 89.951 0.586 90.037 0.77 ;
      RECT 89.865 0.585 89.951 0.771 ;
      RECT 89.815 0.585 89.865 0.772 ;
      RECT 89.801 0.586 89.815 0.772 ;
      RECT 89.715 0.593 89.801 0.773 ;
      RECT 89.641 0.604 89.715 0.774 ;
      RECT 89.555 0.613 89.641 0.775 ;
      RECT 89.52 0.62 89.555 0.79 ;
      RECT 89.495 0.623 89.52 0.82 ;
      RECT 89.47 0.632 89.495 0.849 ;
      RECT 89.46 0.643 89.47 0.869 ;
      RECT 89.45 0.651 89.46 0.883 ;
      RECT 89.445 0.657 89.45 0.893 ;
      RECT 89.42 0.674 89.445 0.91 ;
      RECT 89.405 0.696 89.42 0.938 ;
      RECT 89.375 0.722 89.405 0.968 ;
      RECT 89.355 0.751 89.375 0.998 ;
      RECT 89.35 0.766 89.355 1.015 ;
      RECT 89.33 0.781 89.35 1.03 ;
      RECT 89.32 0.799 89.33 1.048 ;
      RECT 89.31 0.81 89.32 1.063 ;
      RECT 89.26 0.842 89.31 1.089 ;
      RECT 89.255 0.872 89.26 1.109 ;
      RECT 89.245 0.885 89.255 1.115 ;
      RECT 89.236 0.895 89.245 1.123 ;
      RECT 89.225 0.906 89.236 1.131 ;
      RECT 89.22 0.916 89.225 1.137 ;
      RECT 89.205 0.937 89.22 1.144 ;
      RECT 89.19 0.967 89.205 1.152 ;
      RECT 89.155 0.997 89.19 1.158 ;
      RECT 89.13 1.015 89.155 1.165 ;
      RECT 89.08 1.023 89.13 1.174 ;
      RECT 89.055 1.028 89.08 1.183 ;
      RECT 89 1.034 89.055 1.193 ;
      RECT 88.995 1.039 89 1.201 ;
      RECT 88.981 1.042 88.995 1.203 ;
      RECT 88.895 1.054 88.981 1.215 ;
      RECT 88.885 1.066 88.895 1.228 ;
      RECT 88.8 1.079 88.885 1.24 ;
      RECT 88.756 1.096 88.8 1.254 ;
      RECT 88.67 1.113 88.756 1.27 ;
      RECT 88.64 1.127 88.67 1.284 ;
      RECT 88.63 1.132 88.64 1.289 ;
      RECT 88.57 1.135 88.63 1.298 ;
      RECT 91.46 1.405 91.72 1.665 ;
      RECT 91.46 1.405 91.74 1.518 ;
      RECT 91.46 1.405 91.765 1.485 ;
      RECT 91.46 1.405 91.77 1.465 ;
      RECT 91.51 1.18 91.79 1.46 ;
      RECT 91.065 1.915 91.325 2.175 ;
      RECT 91.055 1.772 91.25 2.113 ;
      RECT 91.05 1.88 91.265 2.105 ;
      RECT 91.045 1.93 91.325 2.095 ;
      RECT 91.035 2.007 91.325 2.08 ;
      RECT 91.055 1.855 91.265 2.113 ;
      RECT 91.065 1.73 91.25 2.175 ;
      RECT 91.065 1.625 91.23 2.175 ;
      RECT 91.075 1.612 91.23 2.175 ;
      RECT 91.075 1.57 91.22 2.175 ;
      RECT 91.08 1.495 91.22 2.175 ;
      RECT 91.11 1.145 91.22 2.175 ;
      RECT 91.115 0.875 91.24 1.498 ;
      RECT 91.085 1.45 91.24 1.498 ;
      RECT 91.1 1.252 91.22 2.175 ;
      RECT 91.09 1.362 91.24 1.498 ;
      RECT 91.115 0.875 91.255 1.355 ;
      RECT 91.115 0.875 91.275 1.23 ;
      RECT 91.08 0.875 91.34 1.135 ;
      RECT 90.55 1.18 90.83 1.46 ;
      RECT 90.535 1.18 90.83 1.44 ;
      RECT 88.59 2.045 88.85 2.305 ;
      RECT 90.375 1.9 90.635 2.16 ;
      RECT 90.355 1.92 90.635 2.135 ;
      RECT 90.312 1.92 90.355 2.134 ;
      RECT 90.226 1.921 90.312 2.131 ;
      RECT 90.14 1.922 90.226 2.127 ;
      RECT 90.065 1.924 90.14 2.124 ;
      RECT 90.042 1.925 90.065 2.122 ;
      RECT 89.956 1.926 90.042 2.12 ;
      RECT 89.87 1.927 89.956 2.117 ;
      RECT 89.846 1.928 89.87 2.115 ;
      RECT 89.76 1.93 89.846 2.112 ;
      RECT 89.675 1.932 89.76 2.113 ;
      RECT 89.618 1.933 89.675 2.119 ;
      RECT 89.532 1.935 89.618 2.129 ;
      RECT 89.446 1.938 89.532 2.142 ;
      RECT 89.36 1.94 89.446 2.154 ;
      RECT 89.346 1.941 89.36 2.161 ;
      RECT 89.26 1.942 89.346 2.169 ;
      RECT 89.22 1.944 89.26 2.178 ;
      RECT 89.211 1.945 89.22 2.181 ;
      RECT 89.125 1.953 89.211 2.187 ;
      RECT 89.105 1.962 89.125 2.195 ;
      RECT 89.02 1.977 89.105 2.203 ;
      RECT 88.96 2 89.02 2.214 ;
      RECT 88.95 2.012 88.96 2.219 ;
      RECT 88.91 2.022 88.95 2.223 ;
      RECT 88.855 2.039 88.91 2.231 ;
      RECT 88.85 2.049 88.855 2.235 ;
      RECT 89.916 1.18 89.975 1.577 ;
      RECT 89.83 1.18 90.035 1.568 ;
      RECT 89.825 1.21 90.035 1.563 ;
      RECT 89.791 1.21 90.035 1.561 ;
      RECT 89.705 1.21 90.035 1.555 ;
      RECT 89.66 1.21 90.055 1.533 ;
      RECT 89.66 1.21 90.075 1.488 ;
      RECT 89.62 1.21 90.075 1.478 ;
      RECT 89.83 1.18 90.11 1.46 ;
      RECT 89.565 1.18 89.825 1.44 ;
      RECT 88.75 0.66 89.01 0.92 ;
      RECT 88.83 0.62 89.11 0.9 ;
      RECT 87.39 1.74 87.67 2.02 ;
      RECT 87.36 1.702 87.615 2.005 ;
      RECT 87.355 1.703 87.615 2.003 ;
      RECT 87.35 1.704 87.615 1.997 ;
      RECT 87.345 1.707 87.615 1.99 ;
      RECT 87.34 1.74 87.67 1.983 ;
      RECT 87.31 1.71 87.615 1.97 ;
      RECT 87.31 1.737 87.635 1.97 ;
      RECT 87.31 1.727 87.63 1.97 ;
      RECT 87.31 1.712 87.625 1.97 ;
      RECT 87.39 1.699 87.605 2.02 ;
      RECT 87.476 1.697 87.605 2.02 ;
      RECT 87.562 1.695 87.59 2.02 ;
      RECT 74.72 0.59 75.09 0.96 ;
      RECT 75.235 0.605 75.495 0.93 ;
      RECT 74.72 0.635 75.495 0.895 ;
      RECT 65.505 1.195 65.74 1.455 ;
      RECT 68.65 0.975 68.815 1.235 ;
      RECT 68.555 0.965 68.57 1.235 ;
      RECT 67.155 0.535 67.195 0.675 ;
      RECT 68.57 0.97 68.65 1.235 ;
      RECT 68.515 0.965 68.555 1.201 ;
      RECT 68.501 0.965 68.515 1.201 ;
      RECT 68.415 0.97 68.501 1.203 ;
      RECT 68.37 0.977 68.415 1.205 ;
      RECT 68.34 0.977 68.37 1.207 ;
      RECT 68.315 0.972 68.34 1.209 ;
      RECT 68.285 0.968 68.315 1.218 ;
      RECT 68.275 0.965 68.285 1.23 ;
      RECT 68.27 0.965 68.275 1.238 ;
      RECT 68.265 0.965 68.27 1.243 ;
      RECT 68.255 0.964 68.265 1.253 ;
      RECT 68.25 0.963 68.255 1.263 ;
      RECT 68.235 0.962 68.25 1.268 ;
      RECT 68.207 0.959 68.235 1.295 ;
      RECT 68.121 0.951 68.207 1.295 ;
      RECT 68.035 0.94 68.121 1.295 ;
      RECT 67.995 0.925 68.035 1.295 ;
      RECT 67.955 0.899 67.995 1.295 ;
      RECT 67.95 0.881 67.955 1.107 ;
      RECT 67.94 0.877 67.95 1.097 ;
      RECT 67.925 0.867 67.94 1.084 ;
      RECT 67.905 0.851 67.925 1.069 ;
      RECT 67.89 0.836 67.905 1.054 ;
      RECT 67.88 0.825 67.89 1.044 ;
      RECT 67.855 0.809 67.88 1.033 ;
      RECT 67.85 0.796 67.855 1.023 ;
      RECT 67.845 0.792 67.85 1.018 ;
      RECT 67.79 0.778 67.845 0.996 ;
      RECT 67.751 0.759 67.79 0.96 ;
      RECT 67.665 0.733 67.751 0.913 ;
      RECT 67.661 0.715 67.665 0.879 ;
      RECT 67.575 0.696 67.661 0.857 ;
      RECT 67.57 0.678 67.575 0.835 ;
      RECT 67.565 0.676 67.57 0.833 ;
      RECT 67.555 0.675 67.565 0.828 ;
      RECT 67.495 0.662 67.555 0.814 ;
      RECT 67.45 0.64 67.495 0.793 ;
      RECT 67.39 0.617 67.45 0.772 ;
      RECT 67.326 0.592 67.39 0.747 ;
      RECT 67.24 0.562 67.326 0.716 ;
      RECT 67.225 0.542 67.24 0.695 ;
      RECT 67.195 0.537 67.225 0.686 ;
      RECT 67.142 0.535 67.155 0.675 ;
      RECT 67.056 0.535 67.142 0.677 ;
      RECT 66.97 0.535 67.056 0.679 ;
      RECT 66.95 0.535 66.97 0.683 ;
      RECT 66.905 0.537 66.95 0.694 ;
      RECT 66.865 0.547 66.905 0.71 ;
      RECT 66.861 0.556 66.865 0.718 ;
      RECT 66.775 0.576 66.861 0.734 ;
      RECT 66.765 0.595 66.775 0.752 ;
      RECT 66.76 0.597 66.765 0.755 ;
      RECT 66.75 0.601 66.76 0.758 ;
      RECT 66.73 0.606 66.75 0.768 ;
      RECT 66.7 0.616 66.73 0.788 ;
      RECT 66.695 0.623 66.7 0.802 ;
      RECT 66.685 0.627 66.695 0.809 ;
      RECT 66.67 0.635 66.685 0.82 ;
      RECT 66.66 0.645 66.67 0.831 ;
      RECT 66.65 0.652 66.66 0.839 ;
      RECT 66.625 0.665 66.65 0.854 ;
      RECT 66.561 0.701 66.625 0.893 ;
      RECT 66.475 0.764 66.561 0.957 ;
      RECT 66.44 0.815 66.475 1.01 ;
      RECT 66.435 0.832 66.44 1.027 ;
      RECT 66.42 0.841 66.435 1.034 ;
      RECT 66.4 0.856 66.42 1.048 ;
      RECT 66.395 0.867 66.4 1.058 ;
      RECT 66.375 0.88 66.395 1.068 ;
      RECT 66.37 0.89 66.375 1.078 ;
      RECT 66.355 0.895 66.37 1.087 ;
      RECT 66.345 0.905 66.355 1.098 ;
      RECT 66.315 0.922 66.345 1.115 ;
      RECT 66.305 0.94 66.315 1.133 ;
      RECT 66.29 0.951 66.305 1.144 ;
      RECT 66.25 0.975 66.29 1.16 ;
      RECT 66.215 1.009 66.25 1.177 ;
      RECT 66.185 1.032 66.215 1.189 ;
      RECT 66.17 1.042 66.185 1.198 ;
      RECT 66.13 1.052 66.17 1.209 ;
      RECT 66.11 1.063 66.13 1.221 ;
      RECT 66.105 1.067 66.11 1.228 ;
      RECT 66.09 1.071 66.105 1.233 ;
      RECT 66.08 1.076 66.09 1.238 ;
      RECT 66.075 1.079 66.08 1.241 ;
      RECT 66.045 1.085 66.075 1.248 ;
      RECT 66.01 1.095 66.045 1.262 ;
      RECT 65.95 1.11 66.01 1.282 ;
      RECT 65.895 1.13 65.95 1.306 ;
      RECT 65.866 1.145 65.895 1.324 ;
      RECT 65.78 1.165 65.866 1.349 ;
      RECT 65.775 1.18 65.78 1.369 ;
      RECT 65.765 1.183 65.775 1.37 ;
      RECT 65.74 1.19 65.765 1.455 ;
      RECT 68.435 1.683 68.715 2.02 ;
      RECT 68.435 1.693 68.72 1.978 ;
      RECT 68.435 1.702 68.725 1.875 ;
      RECT 68.435 1.717 68.73 1.743 ;
      RECT 68.435 1.545 68.695 2.02 ;
      RECT 66.155 2.425 66.165 2.615 ;
      RECT 64.415 2.3 64.695 2.58 ;
      RECT 67.46 1.24 67.465 1.725 ;
      RECT 67.355 1.24 67.415 1.5 ;
      RECT 67.68 2.21 67.685 2.285 ;
      RECT 67.67 2.077 67.68 2.32 ;
      RECT 67.66 1.912 67.67 2.341 ;
      RECT 67.655 1.782 67.66 2.357 ;
      RECT 67.645 1.672 67.655 2.373 ;
      RECT 67.64 1.571 67.645 2.39 ;
      RECT 67.635 1.553 67.64 2.4 ;
      RECT 67.63 1.535 67.635 2.41 ;
      RECT 67.62 1.51 67.63 2.425 ;
      RECT 67.615 1.49 67.62 2.44 ;
      RECT 67.595 1.24 67.615 2.465 ;
      RECT 67.58 1.24 67.595 2.498 ;
      RECT 67.55 1.24 67.58 2.52 ;
      RECT 67.53 1.24 67.55 2.534 ;
      RECT 67.51 1.24 67.53 2.05 ;
      RECT 67.525 2.117 67.53 2.539 ;
      RECT 67.52 2.147 67.525 2.541 ;
      RECT 67.515 2.16 67.52 2.544 ;
      RECT 67.51 2.17 67.515 2.548 ;
      RECT 67.505 1.24 67.51 1.968 ;
      RECT 67.505 2.18 67.51 2.55 ;
      RECT 67.5 1.24 67.505 1.945 ;
      RECT 67.49 2.202 67.505 2.55 ;
      RECT 67.485 1.24 67.5 1.89 ;
      RECT 67.48 2.227 67.49 2.55 ;
      RECT 67.48 1.24 67.485 1.835 ;
      RECT 67.47 1.24 67.48 1.783 ;
      RECT 67.475 2.24 67.48 2.551 ;
      RECT 67.47 2.252 67.475 2.552 ;
      RECT 67.465 1.24 67.47 1.743 ;
      RECT 67.465 2.265 67.47 2.553 ;
      RECT 67.45 2.28 67.465 2.554 ;
      RECT 67.455 1.24 67.46 1.705 ;
      RECT 67.45 1.24 67.455 1.67 ;
      RECT 67.445 1.24 67.45 1.645 ;
      RECT 67.44 2.307 67.45 2.556 ;
      RECT 67.435 1.24 67.445 1.603 ;
      RECT 67.435 2.325 67.44 2.557 ;
      RECT 67.43 1.24 67.435 1.563 ;
      RECT 67.43 2.332 67.435 2.558 ;
      RECT 67.425 1.24 67.43 1.535 ;
      RECT 67.42 2.35 67.43 2.559 ;
      RECT 67.415 1.24 67.425 1.515 ;
      RECT 67.41 2.37 67.42 2.561 ;
      RECT 67.4 2.387 67.41 2.562 ;
      RECT 67.365 2.41 67.4 2.565 ;
      RECT 67.31 2.428 67.365 2.571 ;
      RECT 67.224 2.436 67.31 2.58 ;
      RECT 67.138 2.447 67.224 2.591 ;
      RECT 67.052 2.457 67.138 2.602 ;
      RECT 66.966 2.467 67.052 2.614 ;
      RECT 66.88 2.477 66.966 2.625 ;
      RECT 66.86 2.483 66.88 2.631 ;
      RECT 66.78 2.485 66.86 2.635 ;
      RECT 66.775 2.484 66.78 2.64 ;
      RECT 66.767 2.483 66.775 2.64 ;
      RECT 66.681 2.479 66.767 2.638 ;
      RECT 66.595 2.471 66.681 2.635 ;
      RECT 66.509 2.462 66.595 2.631 ;
      RECT 66.423 2.454 66.509 2.628 ;
      RECT 66.337 2.446 66.423 2.624 ;
      RECT 66.251 2.437 66.337 2.621 ;
      RECT 66.165 2.429 66.251 2.617 ;
      RECT 66.11 2.422 66.155 2.615 ;
      RECT 66.025 2.415 66.11 2.613 ;
      RECT 65.951 2.407 66.025 2.609 ;
      RECT 65.865 2.399 65.951 2.606 ;
      RECT 65.862 2.395 65.865 2.604 ;
      RECT 65.776 2.391 65.862 2.603 ;
      RECT 65.69 2.383 65.776 2.6 ;
      RECT 65.605 2.378 65.69 2.597 ;
      RECT 65.519 2.375 65.605 2.594 ;
      RECT 65.433 2.373 65.519 2.591 ;
      RECT 65.347 2.37 65.433 2.588 ;
      RECT 65.261 2.367 65.347 2.585 ;
      RECT 65.175 2.364 65.261 2.582 ;
      RECT 65.099 2.362 65.175 2.579 ;
      RECT 65.013 2.359 65.099 2.576 ;
      RECT 64.927 2.356 65.013 2.574 ;
      RECT 64.841 2.354 64.927 2.571 ;
      RECT 64.755 2.351 64.841 2.568 ;
      RECT 64.695 2.342 64.755 2.566 ;
      RECT 67.205 1.96 67.28 2.22 ;
      RECT 67.185 1.94 67.19 2.22 ;
      RECT 66.505 1.725 66.61 2.02 ;
      RECT 60.95 1.7 61.02 1.96 ;
      RECT 66.845 1.575 66.85 1.946 ;
      RECT 66.835 1.63 66.84 1.946 ;
      RECT 67.14 0.8 67.2 1.06 ;
      RECT 67.195 1.955 67.205 2.22 ;
      RECT 67.19 1.945 67.195 2.22 ;
      RECT 67.11 1.892 67.185 2.22 ;
      RECT 67.135 0.8 67.14 1.08 ;
      RECT 67.125 0.8 67.135 1.1 ;
      RECT 67.11 0.8 67.125 1.13 ;
      RECT 67.095 0.8 67.11 1.173 ;
      RECT 67.09 1.835 67.11 2.22 ;
      RECT 67.08 0.8 67.095 1.21 ;
      RECT 67.075 1.815 67.09 2.22 ;
      RECT 67.075 0.8 67.08 1.233 ;
      RECT 67.065 0.8 67.075 1.258 ;
      RECT 67.035 1.782 67.075 2.22 ;
      RECT 67.04 0.8 67.065 1.308 ;
      RECT 67.035 0.8 67.04 1.363 ;
      RECT 67.03 0.8 67.035 1.405 ;
      RECT 67.02 1.745 67.035 2.22 ;
      RECT 67.025 0.8 67.03 1.448 ;
      RECT 67.02 0.8 67.025 1.513 ;
      RECT 67.015 0.8 67.02 1.535 ;
      RECT 67.015 1.733 67.02 2.085 ;
      RECT 67.01 0.8 67.015 1.603 ;
      RECT 67.01 1.725 67.015 2.068 ;
      RECT 67.005 0.8 67.01 1.648 ;
      RECT 67 1.707 67.01 2.045 ;
      RECT 67 0.8 67.005 1.685 ;
      RECT 66.99 0.8 67 2.025 ;
      RECT 66.985 0.8 66.99 2.008 ;
      RECT 66.98 0.8 66.985 1.993 ;
      RECT 66.975 0.8 66.98 1.978 ;
      RECT 66.955 0.8 66.975 1.968 ;
      RECT 66.95 0.8 66.955 1.958 ;
      RECT 66.94 0.8 66.95 1.954 ;
      RECT 66.935 1.077 66.94 1.953 ;
      RECT 66.93 1.1 66.935 1.952 ;
      RECT 66.925 1.13 66.93 1.951 ;
      RECT 66.92 1.157 66.925 1.95 ;
      RECT 66.915 1.185 66.92 1.95 ;
      RECT 66.91 1.212 66.915 1.95 ;
      RECT 66.905 1.232 66.91 1.95 ;
      RECT 66.9 1.26 66.905 1.95 ;
      RECT 66.89 1.302 66.9 1.95 ;
      RECT 66.88 1.347 66.89 1.949 ;
      RECT 66.875 1.4 66.88 1.948 ;
      RECT 66.87 1.432 66.875 1.947 ;
      RECT 66.865 1.452 66.87 1.946 ;
      RECT 66.86 1.49 66.865 1.946 ;
      RECT 66.855 1.512 66.86 1.946 ;
      RECT 66.85 1.537 66.855 1.946 ;
      RECT 66.84 1.602 66.845 1.946 ;
      RECT 66.825 1.662 66.835 1.946 ;
      RECT 66.81 1.672 66.825 1.946 ;
      RECT 66.79 1.682 66.81 1.946 ;
      RECT 66.76 1.687 66.79 1.943 ;
      RECT 66.7 1.697 66.76 1.94 ;
      RECT 66.68 1.706 66.7 1.945 ;
      RECT 66.655 1.712 66.68 1.958 ;
      RECT 66.635 1.717 66.655 1.973 ;
      RECT 66.61 1.722 66.635 2.02 ;
      RECT 66.481 1.724 66.505 2.02 ;
      RECT 66.395 1.719 66.481 2.02 ;
      RECT 66.355 1.716 66.395 2.02 ;
      RECT 66.305 1.718 66.355 2 ;
      RECT 66.275 1.722 66.305 2 ;
      RECT 66.196 1.732 66.275 2 ;
      RECT 66.11 1.747 66.196 2.001 ;
      RECT 66.06 1.757 66.11 2.002 ;
      RECT 66.052 1.76 66.06 2.002 ;
      RECT 65.966 1.762 66.052 2.003 ;
      RECT 65.88 1.766 65.966 2.003 ;
      RECT 65.794 1.77 65.88 2.004 ;
      RECT 65.708 1.773 65.794 2.005 ;
      RECT 65.622 1.777 65.708 2.005 ;
      RECT 65.536 1.781 65.622 2.006 ;
      RECT 65.45 1.784 65.536 2.007 ;
      RECT 65.364 1.788 65.45 2.007 ;
      RECT 65.278 1.792 65.364 2.008 ;
      RECT 65.192 1.796 65.278 2.009 ;
      RECT 65.106 1.799 65.192 2.009 ;
      RECT 65.02 1.803 65.106 2.01 ;
      RECT 64.99 1.805 65.02 2.01 ;
      RECT 64.904 1.808 64.99 2.011 ;
      RECT 64.818 1.812 64.904 2.012 ;
      RECT 64.732 1.816 64.818 2.013 ;
      RECT 64.646 1.819 64.732 2.013 ;
      RECT 64.56 1.823 64.646 2.014 ;
      RECT 64.525 1.828 64.56 2.015 ;
      RECT 64.47 1.838 64.525 2.022 ;
      RECT 64.445 1.85 64.47 2.032 ;
      RECT 64.41 1.863 64.445 2.04 ;
      RECT 64.37 1.88 64.41 2.063 ;
      RECT 64.35 1.893 64.37 2.09 ;
      RECT 64.32 1.905 64.35 2.118 ;
      RECT 64.315 1.913 64.32 2.138 ;
      RECT 64.31 1.916 64.315 2.148 ;
      RECT 64.26 1.928 64.31 2.182 ;
      RECT 64.25 1.943 64.26 2.215 ;
      RECT 64.24 1.949 64.25 2.228 ;
      RECT 64.23 1.956 64.24 2.24 ;
      RECT 64.205 1.969 64.23 2.258 ;
      RECT 64.19 1.984 64.205 2.28 ;
      RECT 64.18 1.992 64.19 2.296 ;
      RECT 64.165 2.001 64.18 2.311 ;
      RECT 64.155 2.011 64.165 2.325 ;
      RECT 64.136 2.024 64.155 2.342 ;
      RECT 64.05 2.069 64.136 2.407 ;
      RECT 64.035 2.114 64.05 2.465 ;
      RECT 64.03 2.123 64.035 2.478 ;
      RECT 64.02 2.13 64.03 2.483 ;
      RECT 64.015 2.135 64.02 2.487 ;
      RECT 63.995 2.145 64.015 2.494 ;
      RECT 63.97 2.165 63.995 2.508 ;
      RECT 63.935 2.19 63.97 2.528 ;
      RECT 63.92 2.213 63.935 2.543 ;
      RECT 63.91 2.223 63.92 2.548 ;
      RECT 63.9 2.231 63.91 2.555 ;
      RECT 63.89 2.24 63.9 2.561 ;
      RECT 63.87 2.252 63.89 2.563 ;
      RECT 63.86 2.265 63.87 2.565 ;
      RECT 63.835 2.28 63.86 2.568 ;
      RECT 63.815 2.297 63.835 2.572 ;
      RECT 63.775 2.325 63.815 2.578 ;
      RECT 63.71 2.372 63.775 2.587 ;
      RECT 63.695 2.405 63.71 2.595 ;
      RECT 63.69 2.412 63.695 2.597 ;
      RECT 63.64 2.437 63.69 2.602 ;
      RECT 63.625 2.461 63.64 2.609 ;
      RECT 63.575 2.466 63.625 2.61 ;
      RECT 63.489 2.47 63.575 2.61 ;
      RECT 63.403 2.47 63.489 2.61 ;
      RECT 63.317 2.47 63.403 2.611 ;
      RECT 63.231 2.47 63.317 2.611 ;
      RECT 63.145 2.47 63.231 2.611 ;
      RECT 63.079 2.47 63.145 2.611 ;
      RECT 62.993 2.47 63.079 2.612 ;
      RECT 62.907 2.47 62.993 2.612 ;
      RECT 62.821 2.471 62.907 2.613 ;
      RECT 62.735 2.471 62.821 2.613 ;
      RECT 62.649 2.471 62.735 2.613 ;
      RECT 62.563 2.471 62.649 2.614 ;
      RECT 62.477 2.471 62.563 2.614 ;
      RECT 62.391 2.472 62.477 2.615 ;
      RECT 62.305 2.472 62.391 2.615 ;
      RECT 62.285 2.472 62.305 2.615 ;
      RECT 62.199 2.472 62.285 2.615 ;
      RECT 62.113 2.472 62.199 2.615 ;
      RECT 62.027 2.473 62.113 2.615 ;
      RECT 61.941 2.473 62.027 2.615 ;
      RECT 61.855 2.473 61.941 2.615 ;
      RECT 61.769 2.474 61.855 2.615 ;
      RECT 61.683 2.474 61.769 2.615 ;
      RECT 61.597 2.474 61.683 2.615 ;
      RECT 61.511 2.474 61.597 2.615 ;
      RECT 61.425 2.475 61.511 2.615 ;
      RECT 61.375 2.472 61.425 2.615 ;
      RECT 61.365 2.47 61.375 2.614 ;
      RECT 61.361 2.47 61.365 2.613 ;
      RECT 61.275 2.465 61.361 2.608 ;
      RECT 61.253 2.458 61.275 2.602 ;
      RECT 61.167 2.449 61.253 2.596 ;
      RECT 61.081 2.436 61.167 2.587 ;
      RECT 60.995 2.422 61.081 2.577 ;
      RECT 60.95 2.412 60.995 2.57 ;
      RECT 60.93 1.7 60.95 1.978 ;
      RECT 60.93 2.405 60.95 2.566 ;
      RECT 60.9 1.7 60.93 2 ;
      RECT 60.89 2.372 60.93 2.563 ;
      RECT 60.885 1.7 60.9 2.02 ;
      RECT 60.885 2.337 60.89 2.561 ;
      RECT 60.88 1.7 60.885 2.145 ;
      RECT 60.88 2.297 60.885 2.561 ;
      RECT 60.87 1.7 60.88 2.561 ;
      RECT 60.795 1.7 60.87 2.555 ;
      RECT 60.765 1.7 60.795 2.545 ;
      RECT 60.76 1.7 60.765 2.537 ;
      RECT 60.755 1.742 60.76 2.53 ;
      RECT 60.745 1.811 60.755 2.521 ;
      RECT 60.74 1.881 60.745 2.473 ;
      RECT 60.735 1.945 60.74 2.37 ;
      RECT 60.73 1.98 60.735 2.325 ;
      RECT 60.728 2.017 60.73 2.217 ;
      RECT 60.725 2.025 60.728 2.21 ;
      RECT 60.72 2.09 60.725 2.153 ;
      RECT 64.795 1.18 65.075 1.46 ;
      RECT 64.785 1.18 65.075 1.323 ;
      RECT 64.74 1.045 65 1.305 ;
      RECT 64.74 1.16 65.055 1.305 ;
      RECT 64.74 1.13 65.05 1.305 ;
      RECT 64.74 1.117 65.04 1.305 ;
      RECT 64.74 1.107 65.035 1.305 ;
      RECT 60.715 1.09 60.975 1.35 ;
      RECT 64.485 0.64 64.745 0.9 ;
      RECT 64.475 0.665 64.745 0.86 ;
      RECT 64.47 0.665 64.475 0.859 ;
      RECT 64.4 0.66 64.47 0.851 ;
      RECT 64.315 0.647 64.4 0.834 ;
      RECT 64.311 0.639 64.315 0.824 ;
      RECT 64.225 0.632 64.311 0.814 ;
      RECT 64.216 0.624 64.225 0.804 ;
      RECT 64.13 0.617 64.216 0.792 ;
      RECT 64.11 0.608 64.13 0.778 ;
      RECT 64.055 0.603 64.11 0.77 ;
      RECT 64.045 0.597 64.055 0.764 ;
      RECT 64.025 0.595 64.045 0.76 ;
      RECT 64.017 0.594 64.025 0.756 ;
      RECT 63.931 0.586 64.017 0.745 ;
      RECT 63.845 0.572 63.931 0.725 ;
      RECT 63.785 0.56 63.845 0.71 ;
      RECT 63.775 0.555 63.785 0.705 ;
      RECT 63.725 0.555 63.775 0.707 ;
      RECT 63.678 0.557 63.725 0.711 ;
      RECT 63.592 0.564 63.678 0.716 ;
      RECT 63.506 0.572 63.592 0.722 ;
      RECT 63.42 0.581 63.506 0.728 ;
      RECT 63.361 0.587 63.42 0.733 ;
      RECT 63.275 0.592 63.361 0.739 ;
      RECT 63.2 0.597 63.275 0.745 ;
      RECT 63.161 0.599 63.2 0.75 ;
      RECT 63.075 0.596 63.161 0.755 ;
      RECT 62.99 0.594 63.075 0.762 ;
      RECT 62.958 0.593 62.99 0.765 ;
      RECT 62.872 0.592 62.958 0.766 ;
      RECT 62.786 0.591 62.872 0.767 ;
      RECT 62.7 0.59 62.786 0.767 ;
      RECT 62.614 0.589 62.7 0.768 ;
      RECT 62.528 0.588 62.614 0.769 ;
      RECT 62.442 0.587 62.528 0.77 ;
      RECT 62.356 0.586 62.442 0.77 ;
      RECT 62.27 0.585 62.356 0.771 ;
      RECT 62.22 0.585 62.27 0.772 ;
      RECT 62.206 0.586 62.22 0.772 ;
      RECT 62.12 0.593 62.206 0.773 ;
      RECT 62.046 0.604 62.12 0.774 ;
      RECT 61.96 0.613 62.046 0.775 ;
      RECT 61.925 0.62 61.96 0.79 ;
      RECT 61.9 0.623 61.925 0.82 ;
      RECT 61.875 0.632 61.9 0.849 ;
      RECT 61.865 0.643 61.875 0.869 ;
      RECT 61.855 0.651 61.865 0.883 ;
      RECT 61.85 0.657 61.855 0.893 ;
      RECT 61.825 0.674 61.85 0.91 ;
      RECT 61.81 0.696 61.825 0.938 ;
      RECT 61.78 0.722 61.81 0.968 ;
      RECT 61.76 0.751 61.78 0.998 ;
      RECT 61.755 0.766 61.76 1.015 ;
      RECT 61.735 0.781 61.755 1.03 ;
      RECT 61.725 0.799 61.735 1.048 ;
      RECT 61.715 0.81 61.725 1.063 ;
      RECT 61.665 0.842 61.715 1.089 ;
      RECT 61.66 0.872 61.665 1.109 ;
      RECT 61.65 0.885 61.66 1.115 ;
      RECT 61.641 0.895 61.65 1.123 ;
      RECT 61.63 0.906 61.641 1.131 ;
      RECT 61.625 0.916 61.63 1.137 ;
      RECT 61.61 0.937 61.625 1.144 ;
      RECT 61.595 0.967 61.61 1.152 ;
      RECT 61.56 0.997 61.595 1.158 ;
      RECT 61.535 1.015 61.56 1.165 ;
      RECT 61.485 1.023 61.535 1.174 ;
      RECT 61.46 1.028 61.485 1.183 ;
      RECT 61.405 1.034 61.46 1.193 ;
      RECT 61.4 1.039 61.405 1.201 ;
      RECT 61.386 1.042 61.4 1.203 ;
      RECT 61.3 1.054 61.386 1.215 ;
      RECT 61.29 1.066 61.3 1.228 ;
      RECT 61.205 1.079 61.29 1.24 ;
      RECT 61.161 1.096 61.205 1.254 ;
      RECT 61.075 1.113 61.161 1.27 ;
      RECT 61.045 1.127 61.075 1.284 ;
      RECT 61.035 1.132 61.045 1.289 ;
      RECT 60.975 1.135 61.035 1.298 ;
      RECT 63.865 1.405 64.125 1.665 ;
      RECT 63.865 1.405 64.145 1.518 ;
      RECT 63.865 1.405 64.17 1.485 ;
      RECT 63.865 1.405 64.175 1.465 ;
      RECT 63.915 1.18 64.195 1.46 ;
      RECT 63.47 1.915 63.73 2.175 ;
      RECT 63.46 1.772 63.655 2.113 ;
      RECT 63.455 1.88 63.67 2.105 ;
      RECT 63.45 1.93 63.73 2.095 ;
      RECT 63.44 2.007 63.73 2.08 ;
      RECT 63.46 1.855 63.67 2.113 ;
      RECT 63.47 1.73 63.655 2.175 ;
      RECT 63.47 1.625 63.635 2.175 ;
      RECT 63.48 1.612 63.635 2.175 ;
      RECT 63.48 1.57 63.625 2.175 ;
      RECT 63.485 1.495 63.625 2.175 ;
      RECT 63.515 1.145 63.625 2.175 ;
      RECT 63.52 0.875 63.645 1.498 ;
      RECT 63.49 1.45 63.645 1.498 ;
      RECT 63.505 1.252 63.625 2.175 ;
      RECT 63.495 1.362 63.645 1.498 ;
      RECT 63.52 0.875 63.66 1.355 ;
      RECT 63.52 0.875 63.68 1.23 ;
      RECT 63.485 0.875 63.745 1.135 ;
      RECT 62.955 1.18 63.235 1.46 ;
      RECT 62.94 1.18 63.235 1.44 ;
      RECT 60.995 2.045 61.255 2.305 ;
      RECT 62.78 1.9 63.04 2.16 ;
      RECT 62.76 1.92 63.04 2.135 ;
      RECT 62.717 1.92 62.76 2.134 ;
      RECT 62.631 1.921 62.717 2.131 ;
      RECT 62.545 1.922 62.631 2.127 ;
      RECT 62.47 1.924 62.545 2.124 ;
      RECT 62.447 1.925 62.47 2.122 ;
      RECT 62.361 1.926 62.447 2.12 ;
      RECT 62.275 1.927 62.361 2.117 ;
      RECT 62.251 1.928 62.275 2.115 ;
      RECT 62.165 1.93 62.251 2.112 ;
      RECT 62.08 1.932 62.165 2.113 ;
      RECT 62.023 1.933 62.08 2.119 ;
      RECT 61.937 1.935 62.023 2.129 ;
      RECT 61.851 1.938 61.937 2.142 ;
      RECT 61.765 1.94 61.851 2.154 ;
      RECT 61.751 1.941 61.765 2.161 ;
      RECT 61.665 1.942 61.751 2.169 ;
      RECT 61.625 1.944 61.665 2.178 ;
      RECT 61.616 1.945 61.625 2.181 ;
      RECT 61.53 1.953 61.616 2.187 ;
      RECT 61.51 1.962 61.53 2.195 ;
      RECT 61.425 1.977 61.51 2.203 ;
      RECT 61.365 2 61.425 2.214 ;
      RECT 61.355 2.012 61.365 2.219 ;
      RECT 61.315 2.022 61.355 2.223 ;
      RECT 61.26 2.039 61.315 2.231 ;
      RECT 61.255 2.049 61.26 2.235 ;
      RECT 62.321 1.18 62.38 1.577 ;
      RECT 62.235 1.18 62.44 1.568 ;
      RECT 62.23 1.21 62.44 1.563 ;
      RECT 62.196 1.21 62.44 1.561 ;
      RECT 62.11 1.21 62.44 1.555 ;
      RECT 62.065 1.21 62.46 1.533 ;
      RECT 62.065 1.21 62.48 1.488 ;
      RECT 62.025 1.21 62.48 1.478 ;
      RECT 62.235 1.18 62.515 1.46 ;
      RECT 61.97 1.18 62.23 1.44 ;
      RECT 61.155 0.66 61.415 0.92 ;
      RECT 61.235 0.62 61.515 0.9 ;
      RECT 59.795 1.74 60.075 2.02 ;
      RECT 59.765 1.702 60.02 2.005 ;
      RECT 59.76 1.703 60.02 2.003 ;
      RECT 59.755 1.704 60.02 1.997 ;
      RECT 59.75 1.707 60.02 1.99 ;
      RECT 59.745 1.74 60.075 1.983 ;
      RECT 59.715 1.71 60.02 1.97 ;
      RECT 59.715 1.737 60.04 1.97 ;
      RECT 59.715 1.727 60.035 1.97 ;
      RECT 59.715 1.712 60.03 1.97 ;
      RECT 59.795 1.699 60.01 2.02 ;
      RECT 59.881 1.697 60.01 2.02 ;
      RECT 59.967 1.695 59.995 2.02 ;
      RECT 47.125 0.59 47.495 0.96 ;
      RECT 47.64 0.605 47.9 0.93 ;
      RECT 47.125 0.635 47.9 0.895 ;
      RECT 37.91 1.195 38.145 1.455 ;
      RECT 41.055 0.975 41.22 1.235 ;
      RECT 40.96 0.965 40.975 1.235 ;
      RECT 39.56 0.535 39.6 0.675 ;
      RECT 40.975 0.97 41.055 1.235 ;
      RECT 40.92 0.965 40.96 1.201 ;
      RECT 40.906 0.965 40.92 1.201 ;
      RECT 40.82 0.97 40.906 1.203 ;
      RECT 40.775 0.977 40.82 1.205 ;
      RECT 40.745 0.977 40.775 1.207 ;
      RECT 40.72 0.972 40.745 1.209 ;
      RECT 40.69 0.968 40.72 1.218 ;
      RECT 40.68 0.965 40.69 1.23 ;
      RECT 40.675 0.965 40.68 1.238 ;
      RECT 40.67 0.965 40.675 1.243 ;
      RECT 40.66 0.964 40.67 1.253 ;
      RECT 40.655 0.963 40.66 1.263 ;
      RECT 40.64 0.962 40.655 1.268 ;
      RECT 40.612 0.959 40.64 1.295 ;
      RECT 40.526 0.951 40.612 1.295 ;
      RECT 40.44 0.94 40.526 1.295 ;
      RECT 40.4 0.925 40.44 1.295 ;
      RECT 40.36 0.899 40.4 1.295 ;
      RECT 40.355 0.881 40.36 1.107 ;
      RECT 40.345 0.877 40.355 1.097 ;
      RECT 40.33 0.867 40.345 1.084 ;
      RECT 40.31 0.851 40.33 1.069 ;
      RECT 40.295 0.836 40.31 1.054 ;
      RECT 40.285 0.825 40.295 1.044 ;
      RECT 40.26 0.809 40.285 1.033 ;
      RECT 40.255 0.796 40.26 1.023 ;
      RECT 40.25 0.792 40.255 1.018 ;
      RECT 40.195 0.778 40.25 0.996 ;
      RECT 40.156 0.759 40.195 0.96 ;
      RECT 40.07 0.733 40.156 0.913 ;
      RECT 40.066 0.715 40.07 0.879 ;
      RECT 39.98 0.696 40.066 0.857 ;
      RECT 39.975 0.678 39.98 0.835 ;
      RECT 39.97 0.676 39.975 0.833 ;
      RECT 39.96 0.675 39.97 0.828 ;
      RECT 39.9 0.662 39.96 0.814 ;
      RECT 39.855 0.64 39.9 0.793 ;
      RECT 39.795 0.617 39.855 0.772 ;
      RECT 39.731 0.592 39.795 0.747 ;
      RECT 39.645 0.562 39.731 0.716 ;
      RECT 39.63 0.542 39.645 0.695 ;
      RECT 39.6 0.537 39.63 0.686 ;
      RECT 39.547 0.535 39.56 0.675 ;
      RECT 39.461 0.535 39.547 0.677 ;
      RECT 39.375 0.535 39.461 0.679 ;
      RECT 39.355 0.535 39.375 0.683 ;
      RECT 39.31 0.537 39.355 0.694 ;
      RECT 39.27 0.547 39.31 0.71 ;
      RECT 39.266 0.556 39.27 0.718 ;
      RECT 39.18 0.576 39.266 0.734 ;
      RECT 39.17 0.595 39.18 0.752 ;
      RECT 39.165 0.597 39.17 0.755 ;
      RECT 39.155 0.601 39.165 0.758 ;
      RECT 39.135 0.606 39.155 0.768 ;
      RECT 39.105 0.616 39.135 0.788 ;
      RECT 39.1 0.623 39.105 0.802 ;
      RECT 39.09 0.627 39.1 0.809 ;
      RECT 39.075 0.635 39.09 0.82 ;
      RECT 39.065 0.645 39.075 0.831 ;
      RECT 39.055 0.652 39.065 0.839 ;
      RECT 39.03 0.665 39.055 0.854 ;
      RECT 38.966 0.701 39.03 0.893 ;
      RECT 38.88 0.764 38.966 0.957 ;
      RECT 38.845 0.815 38.88 1.01 ;
      RECT 38.84 0.832 38.845 1.027 ;
      RECT 38.825 0.841 38.84 1.034 ;
      RECT 38.805 0.856 38.825 1.048 ;
      RECT 38.8 0.867 38.805 1.058 ;
      RECT 38.78 0.88 38.8 1.068 ;
      RECT 38.775 0.89 38.78 1.078 ;
      RECT 38.76 0.895 38.775 1.087 ;
      RECT 38.75 0.905 38.76 1.098 ;
      RECT 38.72 0.922 38.75 1.115 ;
      RECT 38.71 0.94 38.72 1.133 ;
      RECT 38.695 0.951 38.71 1.144 ;
      RECT 38.655 0.975 38.695 1.16 ;
      RECT 38.62 1.009 38.655 1.177 ;
      RECT 38.59 1.032 38.62 1.189 ;
      RECT 38.575 1.042 38.59 1.198 ;
      RECT 38.535 1.052 38.575 1.209 ;
      RECT 38.515 1.063 38.535 1.221 ;
      RECT 38.51 1.067 38.515 1.228 ;
      RECT 38.495 1.071 38.51 1.233 ;
      RECT 38.485 1.076 38.495 1.238 ;
      RECT 38.48 1.079 38.485 1.241 ;
      RECT 38.45 1.085 38.48 1.248 ;
      RECT 38.415 1.095 38.45 1.262 ;
      RECT 38.355 1.11 38.415 1.282 ;
      RECT 38.3 1.13 38.355 1.306 ;
      RECT 38.271 1.145 38.3 1.324 ;
      RECT 38.185 1.165 38.271 1.349 ;
      RECT 38.18 1.18 38.185 1.369 ;
      RECT 38.17 1.183 38.18 1.37 ;
      RECT 38.145 1.19 38.17 1.455 ;
      RECT 40.84 1.683 41.12 2.02 ;
      RECT 40.84 1.693 41.125 1.978 ;
      RECT 40.84 1.702 41.13 1.875 ;
      RECT 40.84 1.717 41.135 1.743 ;
      RECT 40.84 1.545 41.1 2.02 ;
      RECT 38.56 2.425 38.57 2.615 ;
      RECT 36.82 2.3 37.1 2.58 ;
      RECT 39.865 1.24 39.87 1.725 ;
      RECT 39.76 1.24 39.82 1.5 ;
      RECT 40.085 2.21 40.09 2.285 ;
      RECT 40.075 2.077 40.085 2.32 ;
      RECT 40.065 1.912 40.075 2.341 ;
      RECT 40.06 1.782 40.065 2.357 ;
      RECT 40.05 1.672 40.06 2.373 ;
      RECT 40.045 1.571 40.05 2.39 ;
      RECT 40.04 1.553 40.045 2.4 ;
      RECT 40.035 1.535 40.04 2.41 ;
      RECT 40.025 1.51 40.035 2.425 ;
      RECT 40.02 1.49 40.025 2.44 ;
      RECT 40 1.24 40.02 2.465 ;
      RECT 39.985 1.24 40 2.498 ;
      RECT 39.955 1.24 39.985 2.52 ;
      RECT 39.935 1.24 39.955 2.534 ;
      RECT 39.915 1.24 39.935 2.05 ;
      RECT 39.93 2.117 39.935 2.539 ;
      RECT 39.925 2.147 39.93 2.541 ;
      RECT 39.92 2.16 39.925 2.544 ;
      RECT 39.915 2.17 39.92 2.548 ;
      RECT 39.91 1.24 39.915 1.968 ;
      RECT 39.91 2.18 39.915 2.55 ;
      RECT 39.905 1.24 39.91 1.945 ;
      RECT 39.895 2.202 39.91 2.55 ;
      RECT 39.89 1.24 39.905 1.89 ;
      RECT 39.885 2.227 39.895 2.55 ;
      RECT 39.885 1.24 39.89 1.835 ;
      RECT 39.875 1.24 39.885 1.783 ;
      RECT 39.88 2.24 39.885 2.551 ;
      RECT 39.875 2.252 39.88 2.552 ;
      RECT 39.87 1.24 39.875 1.743 ;
      RECT 39.87 2.265 39.875 2.553 ;
      RECT 39.855 2.28 39.87 2.554 ;
      RECT 39.86 1.24 39.865 1.705 ;
      RECT 39.855 1.24 39.86 1.67 ;
      RECT 39.85 1.24 39.855 1.645 ;
      RECT 39.845 2.307 39.855 2.556 ;
      RECT 39.84 1.24 39.85 1.603 ;
      RECT 39.84 2.325 39.845 2.557 ;
      RECT 39.835 1.24 39.84 1.563 ;
      RECT 39.835 2.332 39.84 2.558 ;
      RECT 39.83 1.24 39.835 1.535 ;
      RECT 39.825 2.35 39.835 2.559 ;
      RECT 39.82 1.24 39.83 1.515 ;
      RECT 39.815 2.37 39.825 2.561 ;
      RECT 39.805 2.387 39.815 2.562 ;
      RECT 39.77 2.41 39.805 2.565 ;
      RECT 39.715 2.428 39.77 2.571 ;
      RECT 39.629 2.436 39.715 2.58 ;
      RECT 39.543 2.447 39.629 2.591 ;
      RECT 39.457 2.457 39.543 2.602 ;
      RECT 39.371 2.467 39.457 2.614 ;
      RECT 39.285 2.477 39.371 2.625 ;
      RECT 39.265 2.483 39.285 2.631 ;
      RECT 39.185 2.485 39.265 2.635 ;
      RECT 39.18 2.484 39.185 2.64 ;
      RECT 39.172 2.483 39.18 2.64 ;
      RECT 39.086 2.479 39.172 2.638 ;
      RECT 39 2.471 39.086 2.635 ;
      RECT 38.914 2.462 39 2.631 ;
      RECT 38.828 2.454 38.914 2.628 ;
      RECT 38.742 2.446 38.828 2.624 ;
      RECT 38.656 2.437 38.742 2.621 ;
      RECT 38.57 2.429 38.656 2.617 ;
      RECT 38.515 2.422 38.56 2.615 ;
      RECT 38.43 2.415 38.515 2.613 ;
      RECT 38.356 2.407 38.43 2.609 ;
      RECT 38.27 2.399 38.356 2.606 ;
      RECT 38.267 2.395 38.27 2.604 ;
      RECT 38.181 2.391 38.267 2.603 ;
      RECT 38.095 2.383 38.181 2.6 ;
      RECT 38.01 2.378 38.095 2.597 ;
      RECT 37.924 2.375 38.01 2.594 ;
      RECT 37.838 2.373 37.924 2.591 ;
      RECT 37.752 2.37 37.838 2.588 ;
      RECT 37.666 2.367 37.752 2.585 ;
      RECT 37.58 2.364 37.666 2.582 ;
      RECT 37.504 2.362 37.58 2.579 ;
      RECT 37.418 2.359 37.504 2.576 ;
      RECT 37.332 2.356 37.418 2.574 ;
      RECT 37.246 2.354 37.332 2.571 ;
      RECT 37.16 2.351 37.246 2.568 ;
      RECT 37.1 2.342 37.16 2.566 ;
      RECT 39.61 1.96 39.685 2.22 ;
      RECT 39.59 1.94 39.595 2.22 ;
      RECT 38.91 1.725 39.015 2.02 ;
      RECT 33.355 1.7 33.425 1.96 ;
      RECT 39.25 1.575 39.255 1.946 ;
      RECT 39.24 1.63 39.245 1.946 ;
      RECT 39.545 0.8 39.605 1.06 ;
      RECT 39.6 1.955 39.61 2.22 ;
      RECT 39.595 1.945 39.6 2.22 ;
      RECT 39.515 1.892 39.59 2.22 ;
      RECT 39.54 0.8 39.545 1.08 ;
      RECT 39.53 0.8 39.54 1.1 ;
      RECT 39.515 0.8 39.53 1.13 ;
      RECT 39.5 0.8 39.515 1.173 ;
      RECT 39.495 1.835 39.515 2.22 ;
      RECT 39.485 0.8 39.5 1.21 ;
      RECT 39.48 1.815 39.495 2.22 ;
      RECT 39.48 0.8 39.485 1.233 ;
      RECT 39.47 0.8 39.48 1.258 ;
      RECT 39.44 1.782 39.48 2.22 ;
      RECT 39.445 0.8 39.47 1.308 ;
      RECT 39.44 0.8 39.445 1.363 ;
      RECT 39.435 0.8 39.44 1.405 ;
      RECT 39.425 1.745 39.44 2.22 ;
      RECT 39.43 0.8 39.435 1.448 ;
      RECT 39.425 0.8 39.43 1.513 ;
      RECT 39.42 0.8 39.425 1.535 ;
      RECT 39.42 1.733 39.425 2.085 ;
      RECT 39.415 0.8 39.42 1.603 ;
      RECT 39.415 1.725 39.42 2.068 ;
      RECT 39.41 0.8 39.415 1.648 ;
      RECT 39.405 1.707 39.415 2.045 ;
      RECT 39.405 0.8 39.41 1.685 ;
      RECT 39.395 0.8 39.405 2.025 ;
      RECT 39.39 0.8 39.395 2.008 ;
      RECT 39.385 0.8 39.39 1.993 ;
      RECT 39.38 0.8 39.385 1.978 ;
      RECT 39.36 0.8 39.38 1.968 ;
      RECT 39.355 0.8 39.36 1.958 ;
      RECT 39.345 0.8 39.355 1.954 ;
      RECT 39.34 1.077 39.345 1.953 ;
      RECT 39.335 1.1 39.34 1.952 ;
      RECT 39.33 1.13 39.335 1.951 ;
      RECT 39.325 1.157 39.33 1.95 ;
      RECT 39.32 1.185 39.325 1.95 ;
      RECT 39.315 1.212 39.32 1.95 ;
      RECT 39.31 1.232 39.315 1.95 ;
      RECT 39.305 1.26 39.31 1.95 ;
      RECT 39.295 1.302 39.305 1.95 ;
      RECT 39.285 1.347 39.295 1.949 ;
      RECT 39.28 1.4 39.285 1.948 ;
      RECT 39.275 1.432 39.28 1.947 ;
      RECT 39.27 1.452 39.275 1.946 ;
      RECT 39.265 1.49 39.27 1.946 ;
      RECT 39.26 1.512 39.265 1.946 ;
      RECT 39.255 1.537 39.26 1.946 ;
      RECT 39.245 1.602 39.25 1.946 ;
      RECT 39.23 1.662 39.24 1.946 ;
      RECT 39.215 1.672 39.23 1.946 ;
      RECT 39.195 1.682 39.215 1.946 ;
      RECT 39.165 1.687 39.195 1.943 ;
      RECT 39.105 1.697 39.165 1.94 ;
      RECT 39.085 1.706 39.105 1.945 ;
      RECT 39.06 1.712 39.085 1.958 ;
      RECT 39.04 1.717 39.06 1.973 ;
      RECT 39.015 1.722 39.04 2.02 ;
      RECT 38.886 1.724 38.91 2.02 ;
      RECT 38.8 1.719 38.886 2.02 ;
      RECT 38.76 1.716 38.8 2.02 ;
      RECT 38.71 1.718 38.76 2 ;
      RECT 38.68 1.722 38.71 2 ;
      RECT 38.601 1.732 38.68 2 ;
      RECT 38.515 1.747 38.601 2.001 ;
      RECT 38.465 1.757 38.515 2.002 ;
      RECT 38.457 1.76 38.465 2.002 ;
      RECT 38.371 1.762 38.457 2.003 ;
      RECT 38.285 1.766 38.371 2.003 ;
      RECT 38.199 1.77 38.285 2.004 ;
      RECT 38.113 1.773 38.199 2.005 ;
      RECT 38.027 1.777 38.113 2.005 ;
      RECT 37.941 1.781 38.027 2.006 ;
      RECT 37.855 1.784 37.941 2.007 ;
      RECT 37.769 1.788 37.855 2.007 ;
      RECT 37.683 1.792 37.769 2.008 ;
      RECT 37.597 1.796 37.683 2.009 ;
      RECT 37.511 1.799 37.597 2.009 ;
      RECT 37.425 1.803 37.511 2.01 ;
      RECT 37.395 1.805 37.425 2.01 ;
      RECT 37.309 1.808 37.395 2.011 ;
      RECT 37.223 1.812 37.309 2.012 ;
      RECT 37.137 1.816 37.223 2.013 ;
      RECT 37.051 1.819 37.137 2.013 ;
      RECT 36.965 1.823 37.051 2.014 ;
      RECT 36.93 1.828 36.965 2.015 ;
      RECT 36.875 1.838 36.93 2.022 ;
      RECT 36.85 1.85 36.875 2.032 ;
      RECT 36.815 1.863 36.85 2.04 ;
      RECT 36.775 1.88 36.815 2.063 ;
      RECT 36.755 1.893 36.775 2.09 ;
      RECT 36.725 1.905 36.755 2.118 ;
      RECT 36.72 1.913 36.725 2.138 ;
      RECT 36.715 1.916 36.72 2.148 ;
      RECT 36.665 1.928 36.715 2.182 ;
      RECT 36.655 1.943 36.665 2.215 ;
      RECT 36.645 1.949 36.655 2.228 ;
      RECT 36.635 1.956 36.645 2.24 ;
      RECT 36.61 1.969 36.635 2.258 ;
      RECT 36.595 1.984 36.61 2.28 ;
      RECT 36.585 1.992 36.595 2.296 ;
      RECT 36.57 2.001 36.585 2.311 ;
      RECT 36.56 2.011 36.57 2.325 ;
      RECT 36.541 2.024 36.56 2.342 ;
      RECT 36.455 2.069 36.541 2.407 ;
      RECT 36.44 2.114 36.455 2.465 ;
      RECT 36.435 2.123 36.44 2.478 ;
      RECT 36.425 2.13 36.435 2.483 ;
      RECT 36.42 2.135 36.425 2.487 ;
      RECT 36.4 2.145 36.42 2.494 ;
      RECT 36.375 2.165 36.4 2.508 ;
      RECT 36.34 2.19 36.375 2.528 ;
      RECT 36.325 2.213 36.34 2.543 ;
      RECT 36.315 2.223 36.325 2.548 ;
      RECT 36.305 2.231 36.315 2.555 ;
      RECT 36.295 2.24 36.305 2.561 ;
      RECT 36.275 2.252 36.295 2.563 ;
      RECT 36.265 2.265 36.275 2.565 ;
      RECT 36.24 2.28 36.265 2.568 ;
      RECT 36.22 2.297 36.24 2.572 ;
      RECT 36.18 2.325 36.22 2.578 ;
      RECT 36.115 2.372 36.18 2.587 ;
      RECT 36.1 2.405 36.115 2.595 ;
      RECT 36.095 2.412 36.1 2.597 ;
      RECT 36.045 2.437 36.095 2.602 ;
      RECT 36.03 2.461 36.045 2.609 ;
      RECT 35.98 2.466 36.03 2.61 ;
      RECT 35.894 2.47 35.98 2.61 ;
      RECT 35.808 2.47 35.894 2.61 ;
      RECT 35.722 2.47 35.808 2.611 ;
      RECT 35.636 2.47 35.722 2.611 ;
      RECT 35.55 2.47 35.636 2.611 ;
      RECT 35.484 2.47 35.55 2.611 ;
      RECT 35.398 2.47 35.484 2.612 ;
      RECT 35.312 2.47 35.398 2.612 ;
      RECT 35.226 2.471 35.312 2.613 ;
      RECT 35.14 2.471 35.226 2.613 ;
      RECT 35.054 2.471 35.14 2.613 ;
      RECT 34.968 2.471 35.054 2.614 ;
      RECT 34.882 2.471 34.968 2.614 ;
      RECT 34.796 2.472 34.882 2.615 ;
      RECT 34.71 2.472 34.796 2.615 ;
      RECT 34.69 2.472 34.71 2.615 ;
      RECT 34.604 2.472 34.69 2.615 ;
      RECT 34.518 2.472 34.604 2.615 ;
      RECT 34.432 2.473 34.518 2.615 ;
      RECT 34.346 2.473 34.432 2.615 ;
      RECT 34.26 2.473 34.346 2.615 ;
      RECT 34.174 2.474 34.26 2.615 ;
      RECT 34.088 2.474 34.174 2.615 ;
      RECT 34.002 2.474 34.088 2.615 ;
      RECT 33.916 2.474 34.002 2.615 ;
      RECT 33.83 2.475 33.916 2.615 ;
      RECT 33.78 2.472 33.83 2.615 ;
      RECT 33.77 2.47 33.78 2.614 ;
      RECT 33.766 2.47 33.77 2.613 ;
      RECT 33.68 2.465 33.766 2.608 ;
      RECT 33.658 2.458 33.68 2.602 ;
      RECT 33.572 2.449 33.658 2.596 ;
      RECT 33.486 2.436 33.572 2.587 ;
      RECT 33.4 2.422 33.486 2.577 ;
      RECT 33.355 2.412 33.4 2.57 ;
      RECT 33.335 1.7 33.355 1.978 ;
      RECT 33.335 2.405 33.355 2.566 ;
      RECT 33.305 1.7 33.335 2 ;
      RECT 33.295 2.372 33.335 2.563 ;
      RECT 33.29 1.7 33.305 2.02 ;
      RECT 33.29 2.337 33.295 2.561 ;
      RECT 33.285 1.7 33.29 2.145 ;
      RECT 33.285 2.297 33.29 2.561 ;
      RECT 33.275 1.7 33.285 2.561 ;
      RECT 33.2 1.7 33.275 2.555 ;
      RECT 33.17 1.7 33.2 2.545 ;
      RECT 33.165 1.7 33.17 2.537 ;
      RECT 33.16 1.742 33.165 2.53 ;
      RECT 33.15 1.811 33.16 2.521 ;
      RECT 33.145 1.881 33.15 2.473 ;
      RECT 33.14 1.945 33.145 2.37 ;
      RECT 33.135 1.98 33.14 2.325 ;
      RECT 33.133 2.017 33.135 2.217 ;
      RECT 33.13 2.025 33.133 2.21 ;
      RECT 33.125 2.09 33.13 2.153 ;
      RECT 37.2 1.18 37.48 1.46 ;
      RECT 37.19 1.18 37.48 1.323 ;
      RECT 37.145 1.045 37.405 1.305 ;
      RECT 37.145 1.16 37.46 1.305 ;
      RECT 37.145 1.13 37.455 1.305 ;
      RECT 37.145 1.117 37.445 1.305 ;
      RECT 37.145 1.107 37.44 1.305 ;
      RECT 33.12 1.09 33.38 1.35 ;
      RECT 36.89 0.64 37.15 0.9 ;
      RECT 36.88 0.665 37.15 0.86 ;
      RECT 36.875 0.665 36.88 0.859 ;
      RECT 36.805 0.66 36.875 0.851 ;
      RECT 36.72 0.647 36.805 0.834 ;
      RECT 36.716 0.639 36.72 0.824 ;
      RECT 36.63 0.632 36.716 0.814 ;
      RECT 36.621 0.624 36.63 0.804 ;
      RECT 36.535 0.617 36.621 0.792 ;
      RECT 36.515 0.608 36.535 0.778 ;
      RECT 36.46 0.603 36.515 0.77 ;
      RECT 36.45 0.597 36.46 0.764 ;
      RECT 36.43 0.595 36.45 0.76 ;
      RECT 36.422 0.594 36.43 0.756 ;
      RECT 36.336 0.586 36.422 0.745 ;
      RECT 36.25 0.572 36.336 0.725 ;
      RECT 36.19 0.56 36.25 0.71 ;
      RECT 36.18 0.555 36.19 0.705 ;
      RECT 36.13 0.555 36.18 0.707 ;
      RECT 36.083 0.557 36.13 0.711 ;
      RECT 35.997 0.564 36.083 0.716 ;
      RECT 35.911 0.572 35.997 0.722 ;
      RECT 35.825 0.581 35.911 0.728 ;
      RECT 35.766 0.587 35.825 0.733 ;
      RECT 35.68 0.592 35.766 0.739 ;
      RECT 35.605 0.597 35.68 0.745 ;
      RECT 35.566 0.599 35.605 0.75 ;
      RECT 35.48 0.596 35.566 0.755 ;
      RECT 35.395 0.594 35.48 0.762 ;
      RECT 35.363 0.593 35.395 0.765 ;
      RECT 35.277 0.592 35.363 0.766 ;
      RECT 35.191 0.591 35.277 0.767 ;
      RECT 35.105 0.59 35.191 0.767 ;
      RECT 35.019 0.589 35.105 0.768 ;
      RECT 34.933 0.588 35.019 0.769 ;
      RECT 34.847 0.587 34.933 0.77 ;
      RECT 34.761 0.586 34.847 0.77 ;
      RECT 34.675 0.585 34.761 0.771 ;
      RECT 34.625 0.585 34.675 0.772 ;
      RECT 34.611 0.586 34.625 0.772 ;
      RECT 34.525 0.593 34.611 0.773 ;
      RECT 34.451 0.604 34.525 0.774 ;
      RECT 34.365 0.613 34.451 0.775 ;
      RECT 34.33 0.62 34.365 0.79 ;
      RECT 34.305 0.623 34.33 0.82 ;
      RECT 34.28 0.632 34.305 0.849 ;
      RECT 34.27 0.643 34.28 0.869 ;
      RECT 34.26 0.651 34.27 0.883 ;
      RECT 34.255 0.657 34.26 0.893 ;
      RECT 34.23 0.674 34.255 0.91 ;
      RECT 34.215 0.696 34.23 0.938 ;
      RECT 34.185 0.722 34.215 0.968 ;
      RECT 34.165 0.751 34.185 0.998 ;
      RECT 34.16 0.766 34.165 1.015 ;
      RECT 34.14 0.781 34.16 1.03 ;
      RECT 34.13 0.799 34.14 1.048 ;
      RECT 34.12 0.81 34.13 1.063 ;
      RECT 34.07 0.842 34.12 1.089 ;
      RECT 34.065 0.872 34.07 1.109 ;
      RECT 34.055 0.885 34.065 1.115 ;
      RECT 34.046 0.895 34.055 1.123 ;
      RECT 34.035 0.906 34.046 1.131 ;
      RECT 34.03 0.916 34.035 1.137 ;
      RECT 34.015 0.937 34.03 1.144 ;
      RECT 34 0.967 34.015 1.152 ;
      RECT 33.965 0.997 34 1.158 ;
      RECT 33.94 1.015 33.965 1.165 ;
      RECT 33.89 1.023 33.94 1.174 ;
      RECT 33.865 1.028 33.89 1.183 ;
      RECT 33.81 1.034 33.865 1.193 ;
      RECT 33.805 1.039 33.81 1.201 ;
      RECT 33.791 1.042 33.805 1.203 ;
      RECT 33.705 1.054 33.791 1.215 ;
      RECT 33.695 1.066 33.705 1.228 ;
      RECT 33.61 1.079 33.695 1.24 ;
      RECT 33.566 1.096 33.61 1.254 ;
      RECT 33.48 1.113 33.566 1.27 ;
      RECT 33.45 1.127 33.48 1.284 ;
      RECT 33.44 1.132 33.45 1.289 ;
      RECT 33.38 1.135 33.44 1.298 ;
      RECT 36.27 1.405 36.53 1.665 ;
      RECT 36.27 1.405 36.55 1.518 ;
      RECT 36.27 1.405 36.575 1.485 ;
      RECT 36.27 1.405 36.58 1.465 ;
      RECT 36.32 1.18 36.6 1.46 ;
      RECT 35.875 1.915 36.135 2.175 ;
      RECT 35.865 1.772 36.06 2.113 ;
      RECT 35.86 1.88 36.075 2.105 ;
      RECT 35.855 1.93 36.135 2.095 ;
      RECT 35.845 2.007 36.135 2.08 ;
      RECT 35.865 1.855 36.075 2.113 ;
      RECT 35.875 1.73 36.06 2.175 ;
      RECT 35.875 1.625 36.04 2.175 ;
      RECT 35.885 1.612 36.04 2.175 ;
      RECT 35.885 1.57 36.03 2.175 ;
      RECT 35.89 1.495 36.03 2.175 ;
      RECT 35.92 1.145 36.03 2.175 ;
      RECT 35.925 0.875 36.05 1.498 ;
      RECT 35.895 1.45 36.05 1.498 ;
      RECT 35.91 1.252 36.03 2.175 ;
      RECT 35.9 1.362 36.05 1.498 ;
      RECT 35.925 0.875 36.065 1.355 ;
      RECT 35.925 0.875 36.085 1.23 ;
      RECT 35.89 0.875 36.15 1.135 ;
      RECT 35.36 1.18 35.64 1.46 ;
      RECT 35.345 1.18 35.64 1.44 ;
      RECT 33.4 2.045 33.66 2.305 ;
      RECT 35.185 1.9 35.445 2.16 ;
      RECT 35.165 1.92 35.445 2.135 ;
      RECT 35.122 1.92 35.165 2.134 ;
      RECT 35.036 1.921 35.122 2.131 ;
      RECT 34.95 1.922 35.036 2.127 ;
      RECT 34.875 1.924 34.95 2.124 ;
      RECT 34.852 1.925 34.875 2.122 ;
      RECT 34.766 1.926 34.852 2.12 ;
      RECT 34.68 1.927 34.766 2.117 ;
      RECT 34.656 1.928 34.68 2.115 ;
      RECT 34.57 1.93 34.656 2.112 ;
      RECT 34.485 1.932 34.57 2.113 ;
      RECT 34.428 1.933 34.485 2.119 ;
      RECT 34.342 1.935 34.428 2.129 ;
      RECT 34.256 1.938 34.342 2.142 ;
      RECT 34.17 1.94 34.256 2.154 ;
      RECT 34.156 1.941 34.17 2.161 ;
      RECT 34.07 1.942 34.156 2.169 ;
      RECT 34.03 1.944 34.07 2.178 ;
      RECT 34.021 1.945 34.03 2.181 ;
      RECT 33.935 1.953 34.021 2.187 ;
      RECT 33.915 1.962 33.935 2.195 ;
      RECT 33.83 1.977 33.915 2.203 ;
      RECT 33.77 2 33.83 2.214 ;
      RECT 33.76 2.012 33.77 2.219 ;
      RECT 33.72 2.022 33.76 2.223 ;
      RECT 33.665 2.039 33.72 2.231 ;
      RECT 33.66 2.049 33.665 2.235 ;
      RECT 34.726 1.18 34.785 1.577 ;
      RECT 34.64 1.18 34.845 1.568 ;
      RECT 34.635 1.21 34.845 1.563 ;
      RECT 34.601 1.21 34.845 1.561 ;
      RECT 34.515 1.21 34.845 1.555 ;
      RECT 34.47 1.21 34.865 1.533 ;
      RECT 34.47 1.21 34.885 1.488 ;
      RECT 34.43 1.21 34.885 1.478 ;
      RECT 34.64 1.18 34.92 1.46 ;
      RECT 34.375 1.18 34.635 1.44 ;
      RECT 33.56 0.66 33.82 0.92 ;
      RECT 33.64 0.62 33.92 0.9 ;
      RECT 32.2 1.74 32.48 2.02 ;
      RECT 32.17 1.702 32.425 2.005 ;
      RECT 32.165 1.703 32.425 2.003 ;
      RECT 32.16 1.704 32.425 1.997 ;
      RECT 32.155 1.707 32.425 1.99 ;
      RECT 32.15 1.74 32.48 1.983 ;
      RECT 32.12 1.71 32.425 1.97 ;
      RECT 32.12 1.737 32.445 1.97 ;
      RECT 32.12 1.727 32.44 1.97 ;
      RECT 32.12 1.712 32.435 1.97 ;
      RECT 32.2 1.699 32.415 2.02 ;
      RECT 32.286 1.697 32.415 2.02 ;
      RECT 32.372 1.695 32.4 2.02 ;
      RECT 19.53 0.59 19.9 0.96 ;
      RECT 20.045 0.605 20.305 0.93 ;
      RECT 19.53 0.635 20.305 0.895 ;
      RECT 10.315 1.195 10.55 1.455 ;
      RECT 13.46 0.975 13.625 1.235 ;
      RECT 13.365 0.965 13.38 1.235 ;
      RECT 11.965 0.535 12.005 0.675 ;
      RECT 13.38 0.97 13.46 1.235 ;
      RECT 13.325 0.965 13.365 1.201 ;
      RECT 13.311 0.965 13.325 1.201 ;
      RECT 13.225 0.97 13.311 1.203 ;
      RECT 13.18 0.977 13.225 1.205 ;
      RECT 13.15 0.977 13.18 1.207 ;
      RECT 13.125 0.972 13.15 1.209 ;
      RECT 13.095 0.968 13.125 1.218 ;
      RECT 13.085 0.965 13.095 1.23 ;
      RECT 13.08 0.965 13.085 1.238 ;
      RECT 13.075 0.965 13.08 1.243 ;
      RECT 13.065 0.964 13.075 1.253 ;
      RECT 13.06 0.963 13.065 1.263 ;
      RECT 13.045 0.962 13.06 1.268 ;
      RECT 13.017 0.959 13.045 1.295 ;
      RECT 12.931 0.951 13.017 1.295 ;
      RECT 12.845 0.94 12.931 1.295 ;
      RECT 12.805 0.925 12.845 1.295 ;
      RECT 12.765 0.899 12.805 1.295 ;
      RECT 12.76 0.881 12.765 1.107 ;
      RECT 12.75 0.877 12.76 1.097 ;
      RECT 12.735 0.867 12.75 1.084 ;
      RECT 12.715 0.851 12.735 1.069 ;
      RECT 12.7 0.836 12.715 1.054 ;
      RECT 12.69 0.825 12.7 1.044 ;
      RECT 12.665 0.809 12.69 1.033 ;
      RECT 12.66 0.796 12.665 1.023 ;
      RECT 12.655 0.792 12.66 1.018 ;
      RECT 12.6 0.778 12.655 0.996 ;
      RECT 12.561 0.759 12.6 0.96 ;
      RECT 12.475 0.733 12.561 0.913 ;
      RECT 12.471 0.715 12.475 0.879 ;
      RECT 12.385 0.696 12.471 0.857 ;
      RECT 12.38 0.678 12.385 0.835 ;
      RECT 12.375 0.676 12.38 0.833 ;
      RECT 12.365 0.675 12.375 0.828 ;
      RECT 12.305 0.662 12.365 0.814 ;
      RECT 12.26 0.64 12.305 0.793 ;
      RECT 12.2 0.617 12.26 0.772 ;
      RECT 12.136 0.592 12.2 0.747 ;
      RECT 12.05 0.562 12.136 0.716 ;
      RECT 12.035 0.542 12.05 0.695 ;
      RECT 12.005 0.537 12.035 0.686 ;
      RECT 11.952 0.535 11.965 0.675 ;
      RECT 11.866 0.535 11.952 0.677 ;
      RECT 11.78 0.535 11.866 0.679 ;
      RECT 11.76 0.535 11.78 0.683 ;
      RECT 11.715 0.537 11.76 0.694 ;
      RECT 11.675 0.547 11.715 0.71 ;
      RECT 11.671 0.556 11.675 0.718 ;
      RECT 11.585 0.576 11.671 0.734 ;
      RECT 11.575 0.595 11.585 0.752 ;
      RECT 11.57 0.597 11.575 0.755 ;
      RECT 11.56 0.601 11.57 0.758 ;
      RECT 11.54 0.606 11.56 0.768 ;
      RECT 11.51 0.616 11.54 0.788 ;
      RECT 11.505 0.623 11.51 0.802 ;
      RECT 11.495 0.627 11.505 0.809 ;
      RECT 11.48 0.635 11.495 0.82 ;
      RECT 11.47 0.645 11.48 0.831 ;
      RECT 11.46 0.652 11.47 0.839 ;
      RECT 11.435 0.665 11.46 0.854 ;
      RECT 11.371 0.701 11.435 0.893 ;
      RECT 11.285 0.764 11.371 0.957 ;
      RECT 11.25 0.815 11.285 1.01 ;
      RECT 11.245 0.832 11.25 1.027 ;
      RECT 11.23 0.841 11.245 1.034 ;
      RECT 11.21 0.856 11.23 1.048 ;
      RECT 11.205 0.867 11.21 1.058 ;
      RECT 11.185 0.88 11.205 1.068 ;
      RECT 11.18 0.89 11.185 1.078 ;
      RECT 11.165 0.895 11.18 1.087 ;
      RECT 11.155 0.905 11.165 1.098 ;
      RECT 11.125 0.922 11.155 1.115 ;
      RECT 11.115 0.94 11.125 1.133 ;
      RECT 11.1 0.951 11.115 1.144 ;
      RECT 11.06 0.975 11.1 1.16 ;
      RECT 11.025 1.009 11.06 1.177 ;
      RECT 10.995 1.032 11.025 1.189 ;
      RECT 10.98 1.042 10.995 1.198 ;
      RECT 10.94 1.052 10.98 1.209 ;
      RECT 10.92 1.063 10.94 1.221 ;
      RECT 10.915 1.067 10.92 1.228 ;
      RECT 10.9 1.071 10.915 1.233 ;
      RECT 10.89 1.076 10.9 1.238 ;
      RECT 10.885 1.079 10.89 1.241 ;
      RECT 10.855 1.085 10.885 1.248 ;
      RECT 10.82 1.095 10.855 1.262 ;
      RECT 10.76 1.11 10.82 1.282 ;
      RECT 10.705 1.13 10.76 1.306 ;
      RECT 10.676 1.145 10.705 1.324 ;
      RECT 10.59 1.165 10.676 1.349 ;
      RECT 10.585 1.18 10.59 1.369 ;
      RECT 10.575 1.183 10.585 1.37 ;
      RECT 10.55 1.19 10.575 1.455 ;
      RECT 13.245 1.683 13.525 2.02 ;
      RECT 13.245 1.693 13.53 1.978 ;
      RECT 13.245 1.702 13.535 1.875 ;
      RECT 13.245 1.717 13.54 1.743 ;
      RECT 13.245 1.545 13.505 2.02 ;
      RECT 10.965 2.425 10.975 2.615 ;
      RECT 9.225 2.3 9.505 2.58 ;
      RECT 12.27 1.24 12.275 1.725 ;
      RECT 12.165 1.24 12.225 1.5 ;
      RECT 12.49 2.21 12.495 2.285 ;
      RECT 12.48 2.077 12.49 2.32 ;
      RECT 12.47 1.912 12.48 2.341 ;
      RECT 12.465 1.782 12.47 2.357 ;
      RECT 12.455 1.672 12.465 2.373 ;
      RECT 12.45 1.571 12.455 2.39 ;
      RECT 12.445 1.553 12.45 2.4 ;
      RECT 12.44 1.535 12.445 2.41 ;
      RECT 12.43 1.51 12.44 2.425 ;
      RECT 12.425 1.49 12.43 2.44 ;
      RECT 12.405 1.24 12.425 2.465 ;
      RECT 12.39 1.24 12.405 2.498 ;
      RECT 12.36 1.24 12.39 2.52 ;
      RECT 12.34 1.24 12.36 2.534 ;
      RECT 12.32 1.24 12.34 2.05 ;
      RECT 12.335 2.117 12.34 2.539 ;
      RECT 12.33 2.147 12.335 2.541 ;
      RECT 12.325 2.16 12.33 2.544 ;
      RECT 12.32 2.17 12.325 2.548 ;
      RECT 12.315 1.24 12.32 1.968 ;
      RECT 12.315 2.18 12.32 2.55 ;
      RECT 12.31 1.24 12.315 1.945 ;
      RECT 12.3 2.202 12.315 2.55 ;
      RECT 12.295 1.24 12.31 1.89 ;
      RECT 12.29 2.227 12.3 2.55 ;
      RECT 12.29 1.24 12.295 1.835 ;
      RECT 12.28 1.24 12.29 1.783 ;
      RECT 12.285 2.24 12.29 2.551 ;
      RECT 12.28 2.252 12.285 2.552 ;
      RECT 12.275 1.24 12.28 1.743 ;
      RECT 12.275 2.265 12.28 2.553 ;
      RECT 12.26 2.28 12.275 2.554 ;
      RECT 12.265 1.24 12.27 1.705 ;
      RECT 12.26 1.24 12.265 1.67 ;
      RECT 12.255 1.24 12.26 1.645 ;
      RECT 12.25 2.307 12.26 2.556 ;
      RECT 12.245 1.24 12.255 1.603 ;
      RECT 12.245 2.325 12.25 2.557 ;
      RECT 12.24 1.24 12.245 1.563 ;
      RECT 12.24 2.332 12.245 2.558 ;
      RECT 12.235 1.24 12.24 1.535 ;
      RECT 12.23 2.35 12.24 2.559 ;
      RECT 12.225 1.24 12.235 1.515 ;
      RECT 12.22 2.37 12.23 2.561 ;
      RECT 12.21 2.387 12.22 2.562 ;
      RECT 12.175 2.41 12.21 2.565 ;
      RECT 12.12 2.428 12.175 2.571 ;
      RECT 12.034 2.436 12.12 2.58 ;
      RECT 11.948 2.447 12.034 2.591 ;
      RECT 11.862 2.457 11.948 2.602 ;
      RECT 11.776 2.467 11.862 2.614 ;
      RECT 11.69 2.477 11.776 2.625 ;
      RECT 11.67 2.483 11.69 2.631 ;
      RECT 11.59 2.485 11.67 2.635 ;
      RECT 11.585 2.484 11.59 2.64 ;
      RECT 11.577 2.483 11.585 2.64 ;
      RECT 11.491 2.479 11.577 2.638 ;
      RECT 11.405 2.471 11.491 2.635 ;
      RECT 11.319 2.462 11.405 2.631 ;
      RECT 11.233 2.454 11.319 2.628 ;
      RECT 11.147 2.446 11.233 2.624 ;
      RECT 11.061 2.437 11.147 2.621 ;
      RECT 10.975 2.429 11.061 2.617 ;
      RECT 10.92 2.422 10.965 2.615 ;
      RECT 10.835 2.415 10.92 2.613 ;
      RECT 10.761 2.407 10.835 2.609 ;
      RECT 10.675 2.399 10.761 2.606 ;
      RECT 10.672 2.395 10.675 2.604 ;
      RECT 10.586 2.391 10.672 2.603 ;
      RECT 10.5 2.383 10.586 2.6 ;
      RECT 10.415 2.378 10.5 2.597 ;
      RECT 10.329 2.375 10.415 2.594 ;
      RECT 10.243 2.373 10.329 2.591 ;
      RECT 10.157 2.37 10.243 2.588 ;
      RECT 10.071 2.367 10.157 2.585 ;
      RECT 9.985 2.364 10.071 2.582 ;
      RECT 9.909 2.362 9.985 2.579 ;
      RECT 9.823 2.359 9.909 2.576 ;
      RECT 9.737 2.356 9.823 2.574 ;
      RECT 9.651 2.354 9.737 2.571 ;
      RECT 9.565 2.351 9.651 2.568 ;
      RECT 9.505 2.342 9.565 2.566 ;
      RECT 12.015 1.96 12.09 2.22 ;
      RECT 11.995 1.94 12 2.22 ;
      RECT 11.315 1.725 11.42 2.02 ;
      RECT 5.76 1.7 5.83 1.96 ;
      RECT 11.655 1.575 11.66 1.946 ;
      RECT 11.645 1.63 11.65 1.946 ;
      RECT 11.95 0.8 12.01 1.06 ;
      RECT 12.005 1.955 12.015 2.22 ;
      RECT 12 1.945 12.005 2.22 ;
      RECT 11.92 1.892 11.995 2.22 ;
      RECT 11.945 0.8 11.95 1.08 ;
      RECT 11.935 0.8 11.945 1.1 ;
      RECT 11.92 0.8 11.935 1.13 ;
      RECT 11.905 0.8 11.92 1.173 ;
      RECT 11.9 1.835 11.92 2.22 ;
      RECT 11.89 0.8 11.905 1.21 ;
      RECT 11.885 1.815 11.9 2.22 ;
      RECT 11.885 0.8 11.89 1.233 ;
      RECT 11.875 0.8 11.885 1.258 ;
      RECT 11.845 1.782 11.885 2.22 ;
      RECT 11.85 0.8 11.875 1.308 ;
      RECT 11.845 0.8 11.85 1.363 ;
      RECT 11.84 0.8 11.845 1.405 ;
      RECT 11.83 1.745 11.845 2.22 ;
      RECT 11.835 0.8 11.84 1.448 ;
      RECT 11.83 0.8 11.835 1.513 ;
      RECT 11.825 0.8 11.83 1.535 ;
      RECT 11.825 1.733 11.83 2.085 ;
      RECT 11.82 0.8 11.825 1.603 ;
      RECT 11.82 1.725 11.825 2.068 ;
      RECT 11.815 0.8 11.82 1.648 ;
      RECT 11.81 1.707 11.82 2.045 ;
      RECT 11.81 0.8 11.815 1.685 ;
      RECT 11.8 0.8 11.81 2.025 ;
      RECT 11.795 0.8 11.8 2.008 ;
      RECT 11.79 0.8 11.795 1.993 ;
      RECT 11.785 0.8 11.79 1.978 ;
      RECT 11.765 0.8 11.785 1.968 ;
      RECT 11.76 0.8 11.765 1.958 ;
      RECT 11.75 0.8 11.76 1.954 ;
      RECT 11.745 1.077 11.75 1.953 ;
      RECT 11.74 1.1 11.745 1.952 ;
      RECT 11.735 1.13 11.74 1.951 ;
      RECT 11.73 1.157 11.735 1.95 ;
      RECT 11.725 1.185 11.73 1.95 ;
      RECT 11.72 1.212 11.725 1.95 ;
      RECT 11.715 1.232 11.72 1.95 ;
      RECT 11.71 1.26 11.715 1.95 ;
      RECT 11.7 1.302 11.71 1.95 ;
      RECT 11.69 1.347 11.7 1.949 ;
      RECT 11.685 1.4 11.69 1.948 ;
      RECT 11.68 1.432 11.685 1.947 ;
      RECT 11.675 1.452 11.68 1.946 ;
      RECT 11.67 1.49 11.675 1.946 ;
      RECT 11.665 1.512 11.67 1.946 ;
      RECT 11.66 1.537 11.665 1.946 ;
      RECT 11.65 1.602 11.655 1.946 ;
      RECT 11.635 1.662 11.645 1.946 ;
      RECT 11.62 1.672 11.635 1.946 ;
      RECT 11.6 1.682 11.62 1.946 ;
      RECT 11.57 1.687 11.6 1.943 ;
      RECT 11.51 1.697 11.57 1.94 ;
      RECT 11.49 1.706 11.51 1.945 ;
      RECT 11.465 1.712 11.49 1.958 ;
      RECT 11.445 1.717 11.465 1.973 ;
      RECT 11.42 1.722 11.445 2.02 ;
      RECT 11.291 1.724 11.315 2.02 ;
      RECT 11.205 1.719 11.291 2.02 ;
      RECT 11.165 1.716 11.205 2.02 ;
      RECT 11.115 1.718 11.165 2 ;
      RECT 11.085 1.722 11.115 2 ;
      RECT 11.006 1.732 11.085 2 ;
      RECT 10.92 1.747 11.006 2.001 ;
      RECT 10.87 1.757 10.92 2.002 ;
      RECT 10.862 1.76 10.87 2.002 ;
      RECT 10.776 1.762 10.862 2.003 ;
      RECT 10.69 1.766 10.776 2.003 ;
      RECT 10.604 1.77 10.69 2.004 ;
      RECT 10.518 1.773 10.604 2.005 ;
      RECT 10.432 1.777 10.518 2.005 ;
      RECT 10.346 1.781 10.432 2.006 ;
      RECT 10.26 1.784 10.346 2.007 ;
      RECT 10.174 1.788 10.26 2.007 ;
      RECT 10.088 1.792 10.174 2.008 ;
      RECT 10.002 1.796 10.088 2.009 ;
      RECT 9.916 1.799 10.002 2.009 ;
      RECT 9.83 1.803 9.916 2.01 ;
      RECT 9.8 1.805 9.83 2.01 ;
      RECT 9.714 1.808 9.8 2.011 ;
      RECT 9.628 1.812 9.714 2.012 ;
      RECT 9.542 1.816 9.628 2.013 ;
      RECT 9.456 1.819 9.542 2.013 ;
      RECT 9.37 1.823 9.456 2.014 ;
      RECT 9.335 1.828 9.37 2.015 ;
      RECT 9.28 1.838 9.335 2.022 ;
      RECT 9.255 1.85 9.28 2.032 ;
      RECT 9.22 1.863 9.255 2.04 ;
      RECT 9.18 1.88 9.22 2.063 ;
      RECT 9.16 1.893 9.18 2.09 ;
      RECT 9.13 1.905 9.16 2.118 ;
      RECT 9.125 1.913 9.13 2.138 ;
      RECT 9.12 1.916 9.125 2.148 ;
      RECT 9.07 1.928 9.12 2.182 ;
      RECT 9.06 1.943 9.07 2.215 ;
      RECT 9.05 1.949 9.06 2.228 ;
      RECT 9.04 1.956 9.05 2.24 ;
      RECT 9.015 1.969 9.04 2.258 ;
      RECT 9 1.984 9.015 2.28 ;
      RECT 8.99 1.992 9 2.296 ;
      RECT 8.975 2.001 8.99 2.311 ;
      RECT 8.965 2.011 8.975 2.325 ;
      RECT 8.946 2.024 8.965 2.342 ;
      RECT 8.86 2.069 8.946 2.407 ;
      RECT 8.845 2.114 8.86 2.465 ;
      RECT 8.84 2.123 8.845 2.478 ;
      RECT 8.83 2.13 8.84 2.483 ;
      RECT 8.825 2.135 8.83 2.487 ;
      RECT 8.805 2.145 8.825 2.494 ;
      RECT 8.78 2.165 8.805 2.508 ;
      RECT 8.745 2.19 8.78 2.528 ;
      RECT 8.73 2.213 8.745 2.543 ;
      RECT 8.72 2.223 8.73 2.548 ;
      RECT 8.71 2.231 8.72 2.555 ;
      RECT 8.7 2.24 8.71 2.561 ;
      RECT 8.68 2.252 8.7 2.563 ;
      RECT 8.67 2.265 8.68 2.565 ;
      RECT 8.645 2.28 8.67 2.568 ;
      RECT 8.625 2.297 8.645 2.572 ;
      RECT 8.585 2.325 8.625 2.578 ;
      RECT 8.52 2.372 8.585 2.587 ;
      RECT 8.505 2.405 8.52 2.595 ;
      RECT 8.5 2.412 8.505 2.597 ;
      RECT 8.45 2.437 8.5 2.602 ;
      RECT 8.435 2.461 8.45 2.609 ;
      RECT 8.385 2.466 8.435 2.61 ;
      RECT 8.299 2.47 8.385 2.61 ;
      RECT 8.213 2.47 8.299 2.61 ;
      RECT 8.127 2.47 8.213 2.611 ;
      RECT 8.041 2.47 8.127 2.611 ;
      RECT 7.955 2.47 8.041 2.611 ;
      RECT 7.889 2.47 7.955 2.611 ;
      RECT 7.803 2.47 7.889 2.612 ;
      RECT 7.717 2.47 7.803 2.612 ;
      RECT 7.631 2.471 7.717 2.613 ;
      RECT 7.545 2.471 7.631 2.613 ;
      RECT 7.459 2.471 7.545 2.613 ;
      RECT 7.373 2.471 7.459 2.614 ;
      RECT 7.287 2.471 7.373 2.614 ;
      RECT 7.201 2.472 7.287 2.615 ;
      RECT 7.115 2.472 7.201 2.615 ;
      RECT 7.095 2.472 7.115 2.615 ;
      RECT 7.009 2.472 7.095 2.615 ;
      RECT 6.923 2.472 7.009 2.615 ;
      RECT 6.837 2.473 6.923 2.615 ;
      RECT 6.751 2.473 6.837 2.615 ;
      RECT 6.665 2.473 6.751 2.615 ;
      RECT 6.579 2.474 6.665 2.615 ;
      RECT 6.493 2.474 6.579 2.615 ;
      RECT 6.407 2.474 6.493 2.615 ;
      RECT 6.321 2.474 6.407 2.615 ;
      RECT 6.235 2.475 6.321 2.615 ;
      RECT 6.185 2.472 6.235 2.615 ;
      RECT 6.175 2.47 6.185 2.614 ;
      RECT 6.171 2.47 6.175 2.613 ;
      RECT 6.085 2.465 6.171 2.608 ;
      RECT 6.063 2.458 6.085 2.602 ;
      RECT 5.977 2.449 6.063 2.596 ;
      RECT 5.891 2.436 5.977 2.587 ;
      RECT 5.805 2.422 5.891 2.577 ;
      RECT 5.76 2.412 5.805 2.57 ;
      RECT 5.74 1.7 5.76 1.978 ;
      RECT 5.74 2.405 5.76 2.566 ;
      RECT 5.71 1.7 5.74 2 ;
      RECT 5.7 2.372 5.74 2.563 ;
      RECT 5.695 1.7 5.71 2.02 ;
      RECT 5.695 2.337 5.7 2.561 ;
      RECT 5.69 1.7 5.695 2.145 ;
      RECT 5.69 2.297 5.695 2.561 ;
      RECT 5.68 1.7 5.69 2.561 ;
      RECT 5.605 1.7 5.68 2.555 ;
      RECT 5.575 1.7 5.605 2.545 ;
      RECT 5.57 1.7 5.575 2.537 ;
      RECT 5.565 1.742 5.57 2.53 ;
      RECT 5.555 1.811 5.565 2.521 ;
      RECT 5.55 1.881 5.555 2.473 ;
      RECT 5.545 1.945 5.55 2.37 ;
      RECT 5.54 1.98 5.545 2.325 ;
      RECT 5.538 2.017 5.54 2.217 ;
      RECT 5.535 2.025 5.538 2.21 ;
      RECT 5.53 2.09 5.535 2.153 ;
      RECT 9.605 1.18 9.885 1.46 ;
      RECT 9.595 1.18 9.885 1.323 ;
      RECT 9.55 1.045 9.81 1.305 ;
      RECT 9.55 1.16 9.865 1.305 ;
      RECT 9.55 1.13 9.86 1.305 ;
      RECT 9.55 1.117 9.85 1.305 ;
      RECT 9.55 1.107 9.845 1.305 ;
      RECT 5.525 1.09 5.785 1.35 ;
      RECT 9.295 0.64 9.555 0.9 ;
      RECT 9.285 0.665 9.555 0.86 ;
      RECT 9.28 0.665 9.285 0.859 ;
      RECT 9.21 0.66 9.28 0.851 ;
      RECT 9.125 0.647 9.21 0.834 ;
      RECT 9.121 0.639 9.125 0.824 ;
      RECT 9.035 0.632 9.121 0.814 ;
      RECT 9.026 0.624 9.035 0.804 ;
      RECT 8.94 0.617 9.026 0.792 ;
      RECT 8.92 0.608 8.94 0.778 ;
      RECT 8.865 0.603 8.92 0.77 ;
      RECT 8.855 0.597 8.865 0.764 ;
      RECT 8.835 0.595 8.855 0.76 ;
      RECT 8.827 0.594 8.835 0.756 ;
      RECT 8.741 0.586 8.827 0.745 ;
      RECT 8.655 0.572 8.741 0.725 ;
      RECT 8.595 0.56 8.655 0.71 ;
      RECT 8.585 0.555 8.595 0.705 ;
      RECT 8.535 0.555 8.585 0.707 ;
      RECT 8.488 0.557 8.535 0.711 ;
      RECT 8.402 0.564 8.488 0.716 ;
      RECT 8.316 0.572 8.402 0.722 ;
      RECT 8.23 0.581 8.316 0.728 ;
      RECT 8.171 0.587 8.23 0.733 ;
      RECT 8.085 0.592 8.171 0.739 ;
      RECT 8.01 0.597 8.085 0.745 ;
      RECT 7.971 0.599 8.01 0.75 ;
      RECT 7.885 0.596 7.971 0.755 ;
      RECT 7.8 0.594 7.885 0.762 ;
      RECT 7.768 0.593 7.8 0.765 ;
      RECT 7.682 0.592 7.768 0.766 ;
      RECT 7.596 0.591 7.682 0.767 ;
      RECT 7.51 0.59 7.596 0.767 ;
      RECT 7.424 0.589 7.51 0.768 ;
      RECT 7.338 0.588 7.424 0.769 ;
      RECT 7.252 0.587 7.338 0.77 ;
      RECT 7.166 0.586 7.252 0.77 ;
      RECT 7.08 0.585 7.166 0.771 ;
      RECT 7.03 0.585 7.08 0.772 ;
      RECT 7.016 0.586 7.03 0.772 ;
      RECT 6.93 0.593 7.016 0.773 ;
      RECT 6.856 0.604 6.93 0.774 ;
      RECT 6.77 0.613 6.856 0.775 ;
      RECT 6.735 0.62 6.77 0.79 ;
      RECT 6.71 0.623 6.735 0.82 ;
      RECT 6.685 0.632 6.71 0.849 ;
      RECT 6.675 0.643 6.685 0.869 ;
      RECT 6.665 0.651 6.675 0.883 ;
      RECT 6.66 0.657 6.665 0.893 ;
      RECT 6.635 0.674 6.66 0.91 ;
      RECT 6.62 0.696 6.635 0.938 ;
      RECT 6.59 0.722 6.62 0.968 ;
      RECT 6.57 0.751 6.59 0.998 ;
      RECT 6.565 0.766 6.57 1.015 ;
      RECT 6.545 0.781 6.565 1.03 ;
      RECT 6.535 0.799 6.545 1.048 ;
      RECT 6.525 0.81 6.535 1.063 ;
      RECT 6.475 0.842 6.525 1.089 ;
      RECT 6.47 0.872 6.475 1.109 ;
      RECT 6.46 0.885 6.47 1.115 ;
      RECT 6.451 0.895 6.46 1.123 ;
      RECT 6.44 0.906 6.451 1.131 ;
      RECT 6.435 0.916 6.44 1.137 ;
      RECT 6.42 0.937 6.435 1.144 ;
      RECT 6.405 0.967 6.42 1.152 ;
      RECT 6.37 0.997 6.405 1.158 ;
      RECT 6.345 1.015 6.37 1.165 ;
      RECT 6.295 1.023 6.345 1.174 ;
      RECT 6.27 1.028 6.295 1.183 ;
      RECT 6.215 1.034 6.27 1.193 ;
      RECT 6.21 1.039 6.215 1.201 ;
      RECT 6.196 1.042 6.21 1.203 ;
      RECT 6.11 1.054 6.196 1.215 ;
      RECT 6.1 1.066 6.11 1.228 ;
      RECT 6.015 1.079 6.1 1.24 ;
      RECT 5.971 1.096 6.015 1.254 ;
      RECT 5.885 1.113 5.971 1.27 ;
      RECT 5.855 1.127 5.885 1.284 ;
      RECT 5.845 1.132 5.855 1.289 ;
      RECT 5.785 1.135 5.845 1.298 ;
      RECT 8.675 1.405 8.935 1.665 ;
      RECT 8.675 1.405 8.955 1.518 ;
      RECT 8.675 1.405 8.98 1.485 ;
      RECT 8.675 1.405 8.985 1.465 ;
      RECT 8.725 1.18 9.005 1.46 ;
      RECT 8.28 1.915 8.54 2.175 ;
      RECT 8.27 1.772 8.465 2.113 ;
      RECT 8.265 1.88 8.48 2.105 ;
      RECT 8.26 1.93 8.54 2.095 ;
      RECT 8.25 2.007 8.54 2.08 ;
      RECT 8.27 1.855 8.48 2.113 ;
      RECT 8.28 1.73 8.465 2.175 ;
      RECT 8.28 1.625 8.445 2.175 ;
      RECT 8.29 1.612 8.445 2.175 ;
      RECT 8.29 1.57 8.435 2.175 ;
      RECT 8.295 1.495 8.435 2.175 ;
      RECT 8.325 1.145 8.435 2.175 ;
      RECT 8.33 0.875 8.455 1.498 ;
      RECT 8.3 1.45 8.455 1.498 ;
      RECT 8.315 1.252 8.435 2.175 ;
      RECT 8.305 1.362 8.455 1.498 ;
      RECT 8.33 0.875 8.47 1.355 ;
      RECT 8.33 0.875 8.49 1.23 ;
      RECT 8.295 0.875 8.555 1.135 ;
      RECT 7.765 1.18 8.045 1.46 ;
      RECT 7.75 1.18 8.045 1.44 ;
      RECT 5.805 2.045 6.065 2.305 ;
      RECT 7.59 1.9 7.85 2.16 ;
      RECT 7.57 1.92 7.85 2.135 ;
      RECT 7.527 1.92 7.57 2.134 ;
      RECT 7.441 1.921 7.527 2.131 ;
      RECT 7.355 1.922 7.441 2.127 ;
      RECT 7.28 1.924 7.355 2.124 ;
      RECT 7.257 1.925 7.28 2.122 ;
      RECT 7.171 1.926 7.257 2.12 ;
      RECT 7.085 1.927 7.171 2.117 ;
      RECT 7.061 1.928 7.085 2.115 ;
      RECT 6.975 1.93 7.061 2.112 ;
      RECT 6.89 1.932 6.975 2.113 ;
      RECT 6.833 1.933 6.89 2.119 ;
      RECT 6.747 1.935 6.833 2.129 ;
      RECT 6.661 1.938 6.747 2.142 ;
      RECT 6.575 1.94 6.661 2.154 ;
      RECT 6.561 1.941 6.575 2.161 ;
      RECT 6.475 1.942 6.561 2.169 ;
      RECT 6.435 1.944 6.475 2.178 ;
      RECT 6.426 1.945 6.435 2.181 ;
      RECT 6.34 1.953 6.426 2.187 ;
      RECT 6.32 1.962 6.34 2.195 ;
      RECT 6.235 1.977 6.32 2.203 ;
      RECT 6.175 2 6.235 2.214 ;
      RECT 6.165 2.012 6.175 2.219 ;
      RECT 6.125 2.022 6.165 2.223 ;
      RECT 6.07 2.039 6.125 2.231 ;
      RECT 6.065 2.049 6.07 2.235 ;
      RECT 7.131 1.18 7.19 1.577 ;
      RECT 7.045 1.18 7.25 1.568 ;
      RECT 7.04 1.21 7.25 1.563 ;
      RECT 7.006 1.21 7.25 1.561 ;
      RECT 6.92 1.21 7.25 1.555 ;
      RECT 6.875 1.21 7.27 1.533 ;
      RECT 6.875 1.21 7.29 1.488 ;
      RECT 6.835 1.21 7.29 1.478 ;
      RECT 7.045 1.18 7.325 1.46 ;
      RECT 6.78 1.18 7.04 1.44 ;
      RECT 5.965 0.66 6.225 0.92 ;
      RECT 6.045 0.62 6.325 0.9 ;
      RECT 4.605 1.74 4.885 2.02 ;
      RECT 4.575 1.702 4.83 2.005 ;
      RECT 4.57 1.703 4.83 2.003 ;
      RECT 4.565 1.704 4.83 1.997 ;
      RECT 4.56 1.707 4.83 1.99 ;
      RECT 4.555 1.74 4.885 1.983 ;
      RECT 4.525 1.71 4.83 1.97 ;
      RECT 4.525 1.737 4.85 1.97 ;
      RECT 4.525 1.727 4.845 1.97 ;
      RECT 4.525 1.712 4.84 1.97 ;
      RECT 4.605 1.699 4.82 2.02 ;
      RECT 4.691 1.697 4.82 2.02 ;
      RECT 4.777 1.695 4.805 2.02 ;
      RECT 134.735 0.8 135.105 1.175 ;
      RECT 131.705 1.61 132.055 1.98 ;
      RECT 130.895 0.74 131.175 1.11 ;
      RECT 127.57 1.61 127.92 1.98 ;
      RECT 126.355 0.68 126.635 1.05 ;
      RECT 125.895 1.4 126.265 1.77 ;
      RECT 124.21 0.06 124.58 0.43 ;
      RECT 113.77 1.61 114.12 1.98 ;
      RECT 112.96 0.67 113.24 1.04 ;
      RECT 110.53 1.71 110.9 2.08 ;
      RECT 104.11 1.61 104.46 1.98 ;
      RECT 103.3 0.74 103.58 1.11 ;
      RECT 99.975 1.61 100.325 1.98 ;
      RECT 98.76 0.68 99.04 1.05 ;
      RECT 98.3 1.4 98.67 1.77 ;
      RECT 96.615 0.06 96.985 0.43 ;
      RECT 86.175 1.61 86.525 1.98 ;
      RECT 85.365 0.67 85.645 1.04 ;
      RECT 82.935 1.71 83.305 2.08 ;
      RECT 76.515 1.61 76.865 1.98 ;
      RECT 75.705 0.74 75.985 1.11 ;
      RECT 72.38 1.61 72.73 1.98 ;
      RECT 71.165 0.68 71.445 1.05 ;
      RECT 70.705 1.4 71.075 1.77 ;
      RECT 69.02 0.06 69.39 0.43 ;
      RECT 58.58 1.61 58.93 1.98 ;
      RECT 57.77 0.67 58.05 1.04 ;
      RECT 55.34 1.71 55.71 2.08 ;
      RECT 48.92 1.61 49.27 1.98 ;
      RECT 48.11 0.74 48.39 1.11 ;
      RECT 44.785 1.61 45.135 1.98 ;
      RECT 43.57 0.68 43.85 1.05 ;
      RECT 43.11 1.4 43.48 1.77 ;
      RECT 41.425 0.06 41.795 0.43 ;
      RECT 30.985 1.61 31.335 1.98 ;
      RECT 30.175 0.67 30.455 1.04 ;
      RECT 27.745 1.71 28.115 2.08 ;
      RECT 21.325 1.61 21.675 1.98 ;
      RECT 20.515 0.74 20.795 1.11 ;
      RECT 17.19 1.61 17.54 1.98 ;
      RECT 15.975 0.68 16.255 1.05 ;
      RECT 15.515 1.4 15.885 1.77 ;
      RECT 13.83 0.06 14.2 0.43 ;
      RECT 3.39 1.61 3.74 1.98 ;
      RECT 2.58 0.67 2.86 1.04 ;
      RECT 0.15 1.71 0.52 2.08 ;
      RECT -2.025 0.595 -1.655 0.965 ;
    LAYER via1 ;
      RECT 134.835 0.9 134.985 1.05 ;
      RECT 131.805 1.71 131.955 1.86 ;
      RECT 130.95 0.84 131.1 0.99 ;
      RECT 130.48 0.69 130.63 0.84 ;
      RECT 127.67 1.71 127.82 1.86 ;
      RECT 126.41 0.78 126.56 0.93 ;
      RECT 125.995 1.5 126.145 1.65 ;
      RECT 124.32 0.17 124.47 0.32 ;
      RECT 123.8 1.03 123.95 1.18 ;
      RECT 123.68 1.6 123.83 1.75 ;
      RECT 122.6 1.295 122.75 1.445 ;
      RECT 122.265 2.015 122.415 2.165 ;
      RECT 122.185 0.855 122.335 1.005 ;
      RECT 120.75 1.25 120.9 1.4 ;
      RECT 119.985 1.1 120.135 1.25 ;
      RECT 119.73 0.695 119.88 0.845 ;
      RECT 119.11 1.46 119.26 1.61 ;
      RECT 118.73 0.93 118.88 1.08 ;
      RECT 118.715 1.97 118.865 2.12 ;
      RECT 118.185 1.235 118.335 1.385 ;
      RECT 118.025 1.955 118.175 2.105 ;
      RECT 117.215 1.235 117.365 1.385 ;
      RECT 116.4 0.715 116.55 0.865 ;
      RECT 116.24 2.1 116.39 2.25 ;
      RECT 116.005 1.755 116.155 1.905 ;
      RECT 115.96 1.145 116.11 1.295 ;
      RECT 114.96 1.765 115.11 1.915 ;
      RECT 113.87 1.71 114.02 1.86 ;
      RECT 113.015 0.77 113.165 0.92 ;
      RECT 110.65 1.81 110.8 1.96 ;
      RECT 104.21 1.71 104.36 1.86 ;
      RECT 103.355 0.84 103.505 0.99 ;
      RECT 102.885 0.69 103.035 0.84 ;
      RECT 100.075 1.71 100.225 1.86 ;
      RECT 98.815 0.78 98.965 0.93 ;
      RECT 98.4 1.5 98.55 1.65 ;
      RECT 96.725 0.17 96.875 0.32 ;
      RECT 96.205 1.03 96.355 1.18 ;
      RECT 96.085 1.6 96.235 1.75 ;
      RECT 95.005 1.295 95.155 1.445 ;
      RECT 94.67 2.015 94.82 2.165 ;
      RECT 94.59 0.855 94.74 1.005 ;
      RECT 93.155 1.25 93.305 1.4 ;
      RECT 92.39 1.1 92.54 1.25 ;
      RECT 92.135 0.695 92.285 0.845 ;
      RECT 91.515 1.46 91.665 1.61 ;
      RECT 91.135 0.93 91.285 1.08 ;
      RECT 91.12 1.97 91.27 2.12 ;
      RECT 90.59 1.235 90.74 1.385 ;
      RECT 90.43 1.955 90.58 2.105 ;
      RECT 89.62 1.235 89.77 1.385 ;
      RECT 88.805 0.715 88.955 0.865 ;
      RECT 88.645 2.1 88.795 2.25 ;
      RECT 88.41 1.755 88.56 1.905 ;
      RECT 88.365 1.145 88.515 1.295 ;
      RECT 87.365 1.765 87.515 1.915 ;
      RECT 86.275 1.71 86.425 1.86 ;
      RECT 85.42 0.77 85.57 0.92 ;
      RECT 83.055 1.81 83.205 1.96 ;
      RECT 76.615 1.71 76.765 1.86 ;
      RECT 75.76 0.84 75.91 0.99 ;
      RECT 75.29 0.69 75.44 0.84 ;
      RECT 72.48 1.71 72.63 1.86 ;
      RECT 71.22 0.78 71.37 0.93 ;
      RECT 70.805 1.5 70.955 1.65 ;
      RECT 69.13 0.17 69.28 0.32 ;
      RECT 68.61 1.03 68.76 1.18 ;
      RECT 68.49 1.6 68.64 1.75 ;
      RECT 67.41 1.295 67.56 1.445 ;
      RECT 67.075 2.015 67.225 2.165 ;
      RECT 66.995 0.855 67.145 1.005 ;
      RECT 65.56 1.25 65.71 1.4 ;
      RECT 64.795 1.1 64.945 1.25 ;
      RECT 64.54 0.695 64.69 0.845 ;
      RECT 63.92 1.46 64.07 1.61 ;
      RECT 63.54 0.93 63.69 1.08 ;
      RECT 63.525 1.97 63.675 2.12 ;
      RECT 62.995 1.235 63.145 1.385 ;
      RECT 62.835 1.955 62.985 2.105 ;
      RECT 62.025 1.235 62.175 1.385 ;
      RECT 61.21 0.715 61.36 0.865 ;
      RECT 61.05 2.1 61.2 2.25 ;
      RECT 60.815 1.755 60.965 1.905 ;
      RECT 60.77 1.145 60.92 1.295 ;
      RECT 59.77 1.765 59.92 1.915 ;
      RECT 58.68 1.71 58.83 1.86 ;
      RECT 57.825 0.77 57.975 0.92 ;
      RECT 55.46 1.81 55.61 1.96 ;
      RECT 49.02 1.71 49.17 1.86 ;
      RECT 48.165 0.84 48.315 0.99 ;
      RECT 47.695 0.69 47.845 0.84 ;
      RECT 44.885 1.71 45.035 1.86 ;
      RECT 43.625 0.78 43.775 0.93 ;
      RECT 43.21 1.5 43.36 1.65 ;
      RECT 41.535 0.17 41.685 0.32 ;
      RECT 41.015 1.03 41.165 1.18 ;
      RECT 40.895 1.6 41.045 1.75 ;
      RECT 39.815 1.295 39.965 1.445 ;
      RECT 39.48 2.015 39.63 2.165 ;
      RECT 39.4 0.855 39.55 1.005 ;
      RECT 37.965 1.25 38.115 1.4 ;
      RECT 37.2 1.1 37.35 1.25 ;
      RECT 36.945 0.695 37.095 0.845 ;
      RECT 36.325 1.46 36.475 1.61 ;
      RECT 35.945 0.93 36.095 1.08 ;
      RECT 35.93 1.97 36.08 2.12 ;
      RECT 35.4 1.235 35.55 1.385 ;
      RECT 35.24 1.955 35.39 2.105 ;
      RECT 34.43 1.235 34.58 1.385 ;
      RECT 33.615 0.715 33.765 0.865 ;
      RECT 33.455 2.1 33.605 2.25 ;
      RECT 33.22 1.755 33.37 1.905 ;
      RECT 33.175 1.145 33.325 1.295 ;
      RECT 32.175 1.765 32.325 1.915 ;
      RECT 31.085 1.71 31.235 1.86 ;
      RECT 30.23 0.77 30.38 0.92 ;
      RECT 27.865 1.81 28.015 1.96 ;
      RECT 21.425 1.71 21.575 1.86 ;
      RECT 20.57 0.84 20.72 0.99 ;
      RECT 20.1 0.69 20.25 0.84 ;
      RECT 17.29 1.71 17.44 1.86 ;
      RECT 16.03 0.78 16.18 0.93 ;
      RECT 15.615 1.5 15.765 1.65 ;
      RECT 13.94 0.17 14.09 0.32 ;
      RECT 13.42 1.03 13.57 1.18 ;
      RECT 13.3 1.6 13.45 1.75 ;
      RECT 12.22 1.295 12.37 1.445 ;
      RECT 11.885 2.015 12.035 2.165 ;
      RECT 11.805 0.855 11.955 1.005 ;
      RECT 10.37 1.25 10.52 1.4 ;
      RECT 9.605 1.1 9.755 1.25 ;
      RECT 9.35 0.695 9.5 0.845 ;
      RECT 8.73 1.46 8.88 1.61 ;
      RECT 8.35 0.93 8.5 1.08 ;
      RECT 8.335 1.97 8.485 2.12 ;
      RECT 7.805 1.235 7.955 1.385 ;
      RECT 7.645 1.955 7.795 2.105 ;
      RECT 6.835 1.235 6.985 1.385 ;
      RECT 6.02 0.715 6.17 0.865 ;
      RECT 5.86 2.1 6.01 2.25 ;
      RECT 5.625 1.755 5.775 1.905 ;
      RECT 5.58 1.145 5.73 1.295 ;
      RECT 4.58 1.765 4.73 1.915 ;
      RECT 3.49 1.71 3.64 1.86 ;
      RECT 2.635 0.77 2.785 0.92 ;
      RECT 0.27 1.81 0.42 1.96 ;
      RECT -1.915 0.705 -1.765 0.855 ;
    LAYER met1 ;
      RECT -3.95 2.72 138.165 3.2 ;
      RECT -1.495 1.67 -1.32 3.2 ;
      RECT -1.555 1.67 -1.265 1.9 ;
      RECT 124.4 2.125 124.705 2.355 ;
      RECT 132.54 2.155 135.955 2.33 ;
      RECT 135.78 1.305 135.955 2.33 ;
      RECT 124.4 2.155 135.955 2.325 ;
      RECT 135.725 1.305 136.055 1.555 ;
      RECT 132.985 1.315 133.275 1.555 ;
      RECT 128.535 1.285 128.795 1.52 ;
      RECT 128.535 1.315 133.275 1.485 ;
      RECT 131.72 1.655 132.04 1.915 ;
      RECT 131.705 1.7 132.04 1.87 ;
      RECT 130.425 0.635 130.72 0.925 ;
      RECT 130.39 0.635 130.72 0.895 ;
      RECT 127.585 1.655 127.905 1.915 ;
      RECT 127.57 1.7 127.905 1.87 ;
      RECT 125.91 1.445 126.23 1.705 ;
      RECT 125.895 1.445 126.25 1.68 ;
      RECT 123.21 1.205 123.395 1.415 ;
      RECT 123.2 1.21 123.41 1.408 ;
      RECT 123.2 1.21 123.496 1.385 ;
      RECT 123.2 1.21 123.555 1.36 ;
      RECT 123.2 1.21 123.61 1.34 ;
      RECT 123.2 1.21 123.62 1.328 ;
      RECT 123.2 1.21 123.815 1.267 ;
      RECT 123.2 1.21 123.845 1.25 ;
      RECT 123.2 1.21 123.865 1.24 ;
      RECT 123.745 0.975 124.005 1.235 ;
      RECT 123.73 1.065 123.745 1.282 ;
      RECT 123.265 1.197 124.005 1.235 ;
      RECT 123.716 1.076 123.73 1.288 ;
      RECT 123.305 1.19 124.005 1.235 ;
      RECT 123.63 1.116 123.716 1.307 ;
      RECT 123.555 1.177 124.005 1.235 ;
      RECT 123.625 1.152 123.63 1.324 ;
      RECT 123.61 1.162 124.005 1.235 ;
      RECT 123.62 1.157 123.625 1.326 ;
      RECT 123.915 1.662 123.92 1.754 ;
      RECT 123.91 1.64 123.915 1.771 ;
      RECT 123.905 1.63 123.91 1.783 ;
      RECT 123.895 1.621 123.905 1.793 ;
      RECT 123.89 1.616 123.895 1.801 ;
      RECT 123.885 1.612 123.89 1.804 ;
      RECT 123.851 1.545 123.885 1.815 ;
      RECT 123.765 1.545 123.851 1.85 ;
      RECT 123.685 1.545 123.765 1.898 ;
      RECT 123.625 1.545 123.685 1.923 ;
      RECT 123.565 1.645 123.625 1.93 ;
      RECT 123.53 1.67 123.565 1.936 ;
      RECT 123.505 1.685 123.53 1.94 ;
      RECT 123.491 1.694 123.505 1.942 ;
      RECT 123.405 1.721 123.491 1.948 ;
      RECT 123.34 1.762 123.405 1.957 ;
      RECT 123.325 1.782 123.34 1.962 ;
      RECT 123.295 1.792 123.325 1.965 ;
      RECT 123.29 1.802 123.295 1.968 ;
      RECT 123.26 1.807 123.29 1.97 ;
      RECT 123.24 1.812 123.26 1.974 ;
      RECT 123.155 1.815 123.24 1.981 ;
      RECT 123.14 1.812 123.155 1.987 ;
      RECT 123.13 1.809 123.14 1.989 ;
      RECT 123.11 1.806 123.13 1.991 ;
      RECT 123.09 1.802 123.11 1.992 ;
      RECT 123.075 1.798 123.09 1.994 ;
      RECT 123.065 1.795 123.075 1.995 ;
      RECT 123.025 1.789 123.065 1.993 ;
      RECT 123.015 1.784 123.025 1.991 ;
      RECT 123 1.781 123.015 1.987 ;
      RECT 122.975 1.776 123 1.98 ;
      RECT 122.925 1.767 122.975 1.968 ;
      RECT 122.855 1.753 122.925 1.95 ;
      RECT 122.797 1.738 122.855 1.932 ;
      RECT 122.711 1.721 122.797 1.912 ;
      RECT 122.625 1.7 122.711 1.887 ;
      RECT 122.575 1.685 122.625 1.868 ;
      RECT 122.571 1.679 122.575 1.86 ;
      RECT 122.485 1.669 122.571 1.847 ;
      RECT 122.45 1.654 122.485 1.83 ;
      RECT 122.435 1.647 122.45 1.823 ;
      RECT 122.375 1.635 122.435 1.811 ;
      RECT 122.355 1.622 122.375 1.799 ;
      RECT 122.315 1.613 122.355 1.791 ;
      RECT 122.31 1.605 122.315 1.784 ;
      RECT 122.23 1.595 122.31 1.77 ;
      RECT 122.215 1.582 122.23 1.755 ;
      RECT 122.21 1.58 122.215 1.753 ;
      RECT 122.131 1.568 122.21 1.74 ;
      RECT 122.045 1.543 122.131 1.715 ;
      RECT 122.03 1.512 122.045 1.7 ;
      RECT 122.015 1.487 122.03 1.696 ;
      RECT 122 1.48 122.015 1.692 ;
      RECT 121.825 1.485 121.83 1.688 ;
      RECT 121.82 1.49 121.825 1.683 ;
      RECT 121.83 1.48 122 1.69 ;
      RECT 122.545 1.24 122.65 1.5 ;
      RECT 123.36 0.765 123.365 0.99 ;
      RECT 123.49 0.765 123.545 0.975 ;
      RECT 123.545 0.77 123.555 0.968 ;
      RECT 123.451 0.765 123.49 0.978 ;
      RECT 123.365 0.765 123.451 0.985 ;
      RECT 123.345 0.77 123.36 0.991 ;
      RECT 123.335 0.81 123.345 0.993 ;
      RECT 123.305 0.82 123.335 0.995 ;
      RECT 123.3 0.825 123.305 0.997 ;
      RECT 123.275 0.83 123.3 0.999 ;
      RECT 123.26 0.835 123.275 1.001 ;
      RECT 123.245 0.837 123.26 1.003 ;
      RECT 123.24 0.842 123.245 1.005 ;
      RECT 123.19 0.85 123.24 1.008 ;
      RECT 123.165 0.859 123.19 1.013 ;
      RECT 123.155 0.866 123.165 1.018 ;
      RECT 123.15 0.869 123.155 1.022 ;
      RECT 123.13 0.872 123.15 1.031 ;
      RECT 123.1 0.88 123.13 1.051 ;
      RECT 123.071 0.893 123.1 1.073 ;
      RECT 122.985 0.927 123.071 1.117 ;
      RECT 122.98 0.953 122.985 1.155 ;
      RECT 122.975 0.957 122.98 1.164 ;
      RECT 122.94 0.97 122.975 1.197 ;
      RECT 122.93 0.984 122.94 1.235 ;
      RECT 122.925 0.988 122.93 1.248 ;
      RECT 122.92 0.992 122.925 1.253 ;
      RECT 122.91 1 122.92 1.265 ;
      RECT 122.905 1.007 122.91 1.28 ;
      RECT 122.88 1.02 122.905 1.305 ;
      RECT 122.84 1.049 122.88 1.36 ;
      RECT 122.825 1.074 122.84 1.415 ;
      RECT 122.815 1.085 122.825 1.438 ;
      RECT 122.81 1.092 122.815 1.45 ;
      RECT 122.805 1.096 122.81 1.458 ;
      RECT 122.75 1.124 122.805 1.5 ;
      RECT 122.73 1.16 122.75 1.5 ;
      RECT 122.715 1.175 122.73 1.5 ;
      RECT 122.66 1.207 122.715 1.5 ;
      RECT 122.65 1.237 122.66 1.5 ;
      RECT 122.26 0.852 122.445 1.09 ;
      RECT 122.245 0.854 122.455 1.085 ;
      RECT 122.13 0.8 122.39 1.06 ;
      RECT 122.125 0.837 122.39 1.014 ;
      RECT 122.12 0.847 122.39 1.011 ;
      RECT 122.115 0.887 122.455 1.005 ;
      RECT 122.11 0.92 122.455 0.995 ;
      RECT 122.12 0.862 122.47 0.933 ;
      RECT 122.417 1.96 122.43 2.49 ;
      RECT 122.331 1.96 122.43 2.489 ;
      RECT 122.331 1.96 122.435 2.488 ;
      RECT 122.245 1.96 122.435 2.486 ;
      RECT 122.24 1.96 122.435 2.483 ;
      RECT 122.24 1.96 122.445 2.481 ;
      RECT 122.235 2.252 122.445 2.478 ;
      RECT 122.235 2.262 122.45 2.475 ;
      RECT 122.235 2.33 122.455 2.471 ;
      RECT 122.225 2.335 122.455 2.47 ;
      RECT 122.225 2.427 122.46 2.467 ;
      RECT 122.21 1.96 122.47 2.22 ;
      RECT 121.44 0.95 121.485 2.485 ;
      RECT 121.64 0.95 121.67 1.165 ;
      RECT 120.015 0.69 120.135 0.9 ;
      RECT 119.675 0.64 119.935 0.9 ;
      RECT 119.675 0.685 119.97 0.89 ;
      RECT 121.68 0.966 121.685 1.02 ;
      RECT 121.675 0.959 121.68 1.153 ;
      RECT 121.67 0.953 121.675 1.16 ;
      RECT 121.625 0.95 121.64 1.173 ;
      RECT 121.62 0.95 121.625 1.195 ;
      RECT 121.615 0.95 121.62 1.243 ;
      RECT 121.61 0.95 121.615 1.263 ;
      RECT 121.6 0.95 121.61 1.37 ;
      RECT 121.595 0.95 121.6 1.433 ;
      RECT 121.59 0.95 121.595 1.49 ;
      RECT 121.585 0.95 121.59 1.498 ;
      RECT 121.57 0.95 121.585 1.605 ;
      RECT 121.56 0.95 121.57 1.74 ;
      RECT 121.55 0.95 121.56 1.85 ;
      RECT 121.54 0.95 121.55 1.907 ;
      RECT 121.535 0.95 121.54 1.947 ;
      RECT 121.53 0.95 121.535 1.983 ;
      RECT 121.52 0.95 121.53 2.023 ;
      RECT 121.515 0.95 121.52 2.065 ;
      RECT 121.495 0.95 121.515 2.13 ;
      RECT 121.5 2.275 121.505 2.455 ;
      RECT 121.495 2.257 121.5 2.463 ;
      RECT 121.49 0.95 121.495 2.193 ;
      RECT 121.49 2.237 121.495 2.47 ;
      RECT 121.485 0.95 121.49 2.48 ;
      RECT 121.43 0.95 121.44 1.25 ;
      RECT 121.435 1.497 121.44 2.485 ;
      RECT 121.43 1.562 121.435 2.485 ;
      RECT 121.425 0.951 121.43 1.24 ;
      RECT 121.42 1.627 121.43 2.485 ;
      RECT 121.415 0.952 121.425 1.23 ;
      RECT 121.405 1.74 121.42 2.485 ;
      RECT 121.41 0.953 121.415 1.22 ;
      RECT 121.39 0.954 121.41 1.198 ;
      RECT 121.395 1.837 121.405 2.485 ;
      RECT 121.39 1.912 121.395 2.485 ;
      RECT 121.38 0.953 121.39 1.175 ;
      RECT 121.385 1.955 121.39 2.485 ;
      RECT 121.38 1.982 121.385 2.485 ;
      RECT 121.37 0.951 121.38 1.163 ;
      RECT 121.375 2.025 121.38 2.485 ;
      RECT 121.37 2.052 121.375 2.485 ;
      RECT 121.36 0.95 121.37 1.15 ;
      RECT 121.365 2.067 121.37 2.485 ;
      RECT 121.325 2.125 121.365 2.485 ;
      RECT 121.355 0.949 121.36 1.135 ;
      RECT 121.35 0.947 121.355 1.128 ;
      RECT 121.34 0.944 121.35 1.118 ;
      RECT 121.335 0.941 121.34 1.103 ;
      RECT 121.32 0.937 121.335 1.096 ;
      RECT 121.315 2.18 121.325 2.485 ;
      RECT 121.315 0.934 121.32 1.091 ;
      RECT 121.3 0.93 121.315 1.085 ;
      RECT 121.31 2.197 121.315 2.485 ;
      RECT 121.3 2.26 121.31 2.485 ;
      RECT 121.22 0.915 121.3 1.065 ;
      RECT 121.295 2.267 121.3 2.48 ;
      RECT 121.29 2.275 121.295 2.47 ;
      RECT 121.21 0.901 121.22 1.049 ;
      RECT 121.195 0.897 121.21 1.047 ;
      RECT 121.185 0.892 121.195 1.043 ;
      RECT 121.16 0.885 121.185 1.035 ;
      RECT 121.155 0.88 121.16 1.03 ;
      RECT 121.145 0.88 121.155 1.028 ;
      RECT 121.135 0.878 121.145 1.026 ;
      RECT 121.105 0.87 121.135 1.02 ;
      RECT 121.09 0.862 121.105 1.013 ;
      RECT 121.07 0.857 121.09 1.006 ;
      RECT 121.065 0.853 121.07 1.001 ;
      RECT 121.035 0.846 121.065 0.995 ;
      RECT 121.01 0.837 121.035 0.985 ;
      RECT 120.98 0.83 121.01 0.977 ;
      RECT 120.955 0.82 120.98 0.968 ;
      RECT 120.94 0.812 120.955 0.962 ;
      RECT 120.915 0.807 120.94 0.957 ;
      RECT 120.905 0.803 120.915 0.952 ;
      RECT 120.885 0.798 120.905 0.947 ;
      RECT 120.85 0.793 120.885 0.94 ;
      RECT 120.79 0.788 120.85 0.933 ;
      RECT 120.777 0.784 120.79 0.931 ;
      RECT 120.691 0.779 120.777 0.928 ;
      RECT 120.605 0.769 120.691 0.924 ;
      RECT 120.564 0.762 120.605 0.921 ;
      RECT 120.478 0.755 120.564 0.918 ;
      RECT 120.392 0.745 120.478 0.914 ;
      RECT 120.306 0.735 120.392 0.909 ;
      RECT 120.22 0.725 120.306 0.905 ;
      RECT 120.21 0.71 120.22 0.903 ;
      RECT 120.2 0.695 120.21 0.903 ;
      RECT 120.135 0.69 120.2 0.902 ;
      RECT 119.97 0.687 120.015 0.895 ;
      RECT 121.215 1.592 121.22 1.783 ;
      RECT 121.21 1.587 121.215 1.79 ;
      RECT 121.196 1.585 121.21 1.796 ;
      RECT 121.11 1.585 121.196 1.798 ;
      RECT 121.106 1.585 121.11 1.801 ;
      RECT 121.02 1.585 121.106 1.819 ;
      RECT 121.01 1.59 121.02 1.838 ;
      RECT 121 1.645 121.01 1.842 ;
      RECT 120.975 1.66 121 1.849 ;
      RECT 120.935 1.68 120.975 1.862 ;
      RECT 120.93 1.692 120.935 1.872 ;
      RECT 120.915 1.698 120.93 1.877 ;
      RECT 120.91 1.703 120.915 1.881 ;
      RECT 120.89 1.71 120.91 1.886 ;
      RECT 120.82 1.735 120.89 1.903 ;
      RECT 120.78 1.763 120.82 1.923 ;
      RECT 120.775 1.773 120.78 1.931 ;
      RECT 120.755 1.78 120.775 1.933 ;
      RECT 120.75 1.787 120.755 1.936 ;
      RECT 120.72 1.795 120.75 1.939 ;
      RECT 120.715 1.8 120.72 1.943 ;
      RECT 120.641 1.804 120.715 1.951 ;
      RECT 120.555 1.813 120.641 1.967 ;
      RECT 120.551 1.818 120.555 1.976 ;
      RECT 120.465 1.823 120.551 1.986 ;
      RECT 120.425 1.831 120.465 1.998 ;
      RECT 120.375 1.837 120.425 2.005 ;
      RECT 120.29 1.846 120.375 2.02 ;
      RECT 120.215 1.857 120.29 2.038 ;
      RECT 120.18 1.864 120.215 2.048 ;
      RECT 120.105 1.872 120.18 2.053 ;
      RECT 120.05 1.881 120.105 2.053 ;
      RECT 120.025 1.886 120.05 2.051 ;
      RECT 120.015 1.889 120.025 2.049 ;
      RECT 119.98 1.891 120.015 2.047 ;
      RECT 119.95 1.893 119.98 2.043 ;
      RECT 119.905 1.892 119.95 2.039 ;
      RECT 119.885 1.887 119.905 2.036 ;
      RECT 119.835 1.872 119.885 2.033 ;
      RECT 119.825 1.857 119.835 2.028 ;
      RECT 119.775 1.842 119.825 2.018 ;
      RECT 119.725 1.817 119.775 1.998 ;
      RECT 119.715 1.802 119.725 1.98 ;
      RECT 119.71 1.8 119.715 1.974 ;
      RECT 119.69 1.795 119.71 1.969 ;
      RECT 119.685 1.787 119.69 1.963 ;
      RECT 119.67 1.781 119.685 1.956 ;
      RECT 119.665 1.776 119.67 1.948 ;
      RECT 119.645 1.771 119.665 1.94 ;
      RECT 119.63 1.764 119.645 1.933 ;
      RECT 119.615 1.758 119.63 1.924 ;
      RECT 119.61 1.752 119.615 1.917 ;
      RECT 119.565 1.727 119.61 1.903 ;
      RECT 119.55 1.697 119.565 1.885 ;
      RECT 119.535 1.68 119.55 1.876 ;
      RECT 119.51 1.66 119.535 1.864 ;
      RECT 119.47 1.63 119.51 1.844 ;
      RECT 119.46 1.6 119.47 1.829 ;
      RECT 119.445 1.59 119.46 1.822 ;
      RECT 119.39 1.555 119.445 1.801 ;
      RECT 119.375 1.518 119.39 1.78 ;
      RECT 119.365 1.505 119.375 1.772 ;
      RECT 119.315 1.475 119.365 1.754 ;
      RECT 119.3 1.405 119.315 1.735 ;
      RECT 119.255 1.405 119.3 1.718 ;
      RECT 119.23 1.405 119.255 1.7 ;
      RECT 119.22 1.405 119.23 1.693 ;
      RECT 119.141 1.405 119.22 1.686 ;
      RECT 119.055 1.405 119.141 1.678 ;
      RECT 119.04 1.437 119.055 1.673 ;
      RECT 118.965 1.447 119.04 1.669 ;
      RECT 118.945 1.457 118.965 1.664 ;
      RECT 118.92 1.457 118.945 1.661 ;
      RECT 118.91 1.447 118.92 1.66 ;
      RECT 118.9 1.42 118.91 1.659 ;
      RECT 118.86 1.415 118.9 1.657 ;
      RECT 118.815 1.415 118.86 1.653 ;
      RECT 118.79 1.415 118.815 1.648 ;
      RECT 118.74 1.415 118.79 1.635 ;
      RECT 118.7 1.42 118.71 1.62 ;
      RECT 118.71 1.415 118.74 1.625 ;
      RECT 120.695 1.195 120.955 1.455 ;
      RECT 120.69 1.217 120.955 1.413 ;
      RECT 119.93 1.045 120.15 1.41 ;
      RECT 119.912 1.132 120.15 1.409 ;
      RECT 119.895 1.137 120.15 1.406 ;
      RECT 119.895 1.137 120.17 1.405 ;
      RECT 119.865 1.147 120.17 1.403 ;
      RECT 119.86 1.162 120.17 1.399 ;
      RECT 119.86 1.162 120.175 1.398 ;
      RECT 119.855 1.22 120.175 1.396 ;
      RECT 119.855 1.22 120.185 1.393 ;
      RECT 119.85 1.285 120.185 1.388 ;
      RECT 119.93 1.045 120.19 1.305 ;
      RECT 118.675 0.875 118.935 1.135 ;
      RECT 118.675 0.918 119.021 1.109 ;
      RECT 118.675 0.918 119.065 1.108 ;
      RECT 118.675 0.918 119.085 1.106 ;
      RECT 118.675 0.918 119.185 1.105 ;
      RECT 118.675 0.918 119.205 1.103 ;
      RECT 118.675 0.918 119.215 1.098 ;
      RECT 119.085 0.885 119.275 1.095 ;
      RECT 119.085 0.887 119.28 1.093 ;
      RECT 119.075 0.892 119.285 1.085 ;
      RECT 119.021 0.916 119.285 1.085 ;
      RECT 119.065 0.91 119.075 1.107 ;
      RECT 119.075 0.89 119.28 1.093 ;
      RECT 118.03 1.95 118.235 2.18 ;
      RECT 117.97 1.9 118.025 2.16 ;
      RECT 118.03 1.9 118.23 2.18 ;
      RECT 119 2.215 119.005 2.242 ;
      RECT 118.99 2.125 119 2.247 ;
      RECT 118.985 2.047 118.99 2.253 ;
      RECT 118.975 2.037 118.985 2.26 ;
      RECT 118.97 2.027 118.975 2.266 ;
      RECT 118.96 2.022 118.97 2.268 ;
      RECT 118.945 2.014 118.96 2.276 ;
      RECT 118.93 2.005 118.945 2.288 ;
      RECT 118.92 1.997 118.93 2.298 ;
      RECT 118.885 1.915 118.92 2.316 ;
      RECT 118.85 1.915 118.885 2.335 ;
      RECT 118.835 1.915 118.85 2.343 ;
      RECT 118.78 1.915 118.835 2.343 ;
      RECT 118.746 1.915 118.78 2.334 ;
      RECT 118.66 1.915 118.746 2.31 ;
      RECT 118.65 1.975 118.66 2.292 ;
      RECT 118.61 1.977 118.65 2.283 ;
      RECT 118.605 1.979 118.61 2.273 ;
      RECT 118.585 1.981 118.605 2.268 ;
      RECT 118.575 1.984 118.585 2.263 ;
      RECT 118.565 1.985 118.575 2.258 ;
      RECT 118.541 1.986 118.565 2.25 ;
      RECT 118.455 1.991 118.541 2.228 ;
      RECT 118.4 1.99 118.455 2.201 ;
      RECT 118.385 1.983 118.4 2.188 ;
      RECT 118.35 1.978 118.385 2.184 ;
      RECT 118.295 1.97 118.35 2.183 ;
      RECT 118.235 1.957 118.295 2.181 ;
      RECT 118.025 1.9 118.03 2.168 ;
      RECT 118.1 1.27 118.285 1.48 ;
      RECT 118.09 1.275 118.3 1.473 ;
      RECT 118.13 1.18 118.39 1.44 ;
      RECT 118.085 1.337 118.39 1.363 ;
      RECT 117.43 1.13 117.435 1.93 ;
      RECT 117.375 1.18 117.405 1.93 ;
      RECT 117.365 1.18 117.37 1.49 ;
      RECT 117.35 1.18 117.355 1.485 ;
      RECT 116.895 1.225 116.91 1.44 ;
      RECT 116.825 1.225 116.91 1.435 ;
      RECT 118.09 0.805 118.16 1.015 ;
      RECT 118.16 0.812 118.17 1.01 ;
      RECT 118.056 0.805 118.09 1.022 ;
      RECT 117.97 0.805 118.056 1.046 ;
      RECT 117.96 0.81 117.97 1.065 ;
      RECT 117.955 0.822 117.96 1.068 ;
      RECT 117.94 0.837 117.955 1.072 ;
      RECT 117.935 0.855 117.94 1.076 ;
      RECT 117.895 0.865 117.935 1.085 ;
      RECT 117.88 0.872 117.895 1.097 ;
      RECT 117.865 0.877 117.88 1.102 ;
      RECT 117.85 0.88 117.865 1.107 ;
      RECT 117.84 0.882 117.85 1.111 ;
      RECT 117.805 0.889 117.84 1.119 ;
      RECT 117.77 0.897 117.805 1.133 ;
      RECT 117.76 0.903 117.77 1.142 ;
      RECT 117.755 0.905 117.76 1.144 ;
      RECT 117.735 0.908 117.755 1.15 ;
      RECT 117.705 0.915 117.735 1.161 ;
      RECT 117.695 0.921 117.705 1.168 ;
      RECT 117.67 0.924 117.695 1.175 ;
      RECT 117.66 0.928 117.67 1.183 ;
      RECT 117.655 0.929 117.66 1.205 ;
      RECT 117.65 0.93 117.655 1.22 ;
      RECT 117.645 0.931 117.65 1.235 ;
      RECT 117.64 0.932 117.645 1.25 ;
      RECT 117.635 0.933 117.64 1.28 ;
      RECT 117.625 0.935 117.635 1.313 ;
      RECT 117.61 0.939 117.625 1.36 ;
      RECT 117.6 0.942 117.61 1.405 ;
      RECT 117.595 0.945 117.6 1.433 ;
      RECT 117.585 0.947 117.595 1.46 ;
      RECT 117.58 0.95 117.585 1.495 ;
      RECT 117.55 0.955 117.58 1.553 ;
      RECT 117.545 0.96 117.55 1.638 ;
      RECT 117.54 0.962 117.545 1.673 ;
      RECT 117.535 0.964 117.54 1.755 ;
      RECT 117.53 0.966 117.535 1.843 ;
      RECT 117.52 0.968 117.53 1.925 ;
      RECT 117.505 0.982 117.52 1.93 ;
      RECT 117.47 1.027 117.505 1.93 ;
      RECT 117.46 1.067 117.47 1.93 ;
      RECT 117.445 1.095 117.46 1.93 ;
      RECT 117.44 1.112 117.445 1.93 ;
      RECT 117.435 1.12 117.44 1.93 ;
      RECT 117.425 1.135 117.43 1.93 ;
      RECT 117.42 1.142 117.425 1.93 ;
      RECT 117.41 1.162 117.42 1.93 ;
      RECT 117.405 1.175 117.41 1.93 ;
      RECT 117.37 1.18 117.375 1.515 ;
      RECT 117.355 1.57 117.375 1.93 ;
      RECT 117.355 1.18 117.365 1.488 ;
      RECT 117.35 1.61 117.355 1.93 ;
      RECT 117.3 1.18 117.35 1.483 ;
      RECT 117.345 1.647 117.35 1.93 ;
      RECT 117.335 1.67 117.345 1.93 ;
      RECT 117.33 1.715 117.335 1.93 ;
      RECT 117.32 1.725 117.33 1.923 ;
      RECT 117.246 1.18 117.3 1.477 ;
      RECT 117.16 1.18 117.246 1.47 ;
      RECT 117.111 1.227 117.16 1.463 ;
      RECT 117.025 1.235 117.111 1.456 ;
      RECT 117.01 1.232 117.025 1.451 ;
      RECT 116.996 1.225 117.01 1.45 ;
      RECT 116.91 1.225 116.996 1.445 ;
      RECT 116.815 1.23 116.825 1.43 ;
      RECT 116.405 0.66 116.42 1.06 ;
      RECT 116.6 0.66 116.605 0.92 ;
      RECT 116.345 0.66 116.39 0.92 ;
      RECT 116.8 1.965 116.805 2.17 ;
      RECT 116.795 1.955 116.8 2.175 ;
      RECT 116.79 1.942 116.795 2.18 ;
      RECT 116.785 1.922 116.79 2.18 ;
      RECT 116.76 1.875 116.785 2.18 ;
      RECT 116.725 1.79 116.76 2.18 ;
      RECT 116.72 1.727 116.725 2.18 ;
      RECT 116.715 1.712 116.72 2.18 ;
      RECT 116.7 1.672 116.715 2.18 ;
      RECT 116.695 1.647 116.7 2.18 ;
      RECT 116.685 1.63 116.695 2.18 ;
      RECT 116.65 1.552 116.685 2.18 ;
      RECT 116.645 1.495 116.65 2.18 ;
      RECT 116.64 1.482 116.645 2.18 ;
      RECT 116.63 1.46 116.64 2.18 ;
      RECT 116.62 1.425 116.63 2.18 ;
      RECT 116.61 1.395 116.62 2.18 ;
      RECT 116.6 1.31 116.61 1.823 ;
      RECT 116.607 1.955 116.61 2.18 ;
      RECT 116.605 1.965 116.607 2.18 ;
      RECT 116.595 1.975 116.605 2.175 ;
      RECT 116.59 0.66 116.6 1.055 ;
      RECT 116.595 1.187 116.6 1.798 ;
      RECT 116.59 1.085 116.595 1.781 ;
      RECT 116.58 0.66 116.59 1.757 ;
      RECT 116.575 0.66 116.58 1.728 ;
      RECT 116.57 0.66 116.575 1.718 ;
      RECT 116.55 0.66 116.57 1.68 ;
      RECT 116.545 0.66 116.55 1.638 ;
      RECT 116.54 0.66 116.545 1.618 ;
      RECT 116.51 0.66 116.54 1.568 ;
      RECT 116.5 0.66 116.51 1.515 ;
      RECT 116.495 0.66 116.5 1.488 ;
      RECT 116.49 0.66 116.495 1.473 ;
      RECT 116.48 0.66 116.49 1.45 ;
      RECT 116.47 0.66 116.48 1.425 ;
      RECT 116.465 0.66 116.47 1.365 ;
      RECT 116.455 0.66 116.465 1.303 ;
      RECT 116.45 0.66 116.455 1.223 ;
      RECT 116.445 0.66 116.45 1.188 ;
      RECT 116.44 0.66 116.445 1.163 ;
      RECT 116.435 0.66 116.44 1.148 ;
      RECT 116.43 0.66 116.435 1.118 ;
      RECT 116.425 0.66 116.43 1.095 ;
      RECT 116.42 0.66 116.425 1.068 ;
      RECT 116.39 0.66 116.405 1.055 ;
      RECT 115.545 2.195 115.73 2.405 ;
      RECT 115.535 2.2 115.745 2.398 ;
      RECT 115.535 2.2 115.765 2.37 ;
      RECT 115.535 2.2 115.78 2.349 ;
      RECT 115.535 2.2 115.795 2.347 ;
      RECT 115.535 2.2 115.805 2.346 ;
      RECT 115.535 2.2 115.835 2.343 ;
      RECT 116.185 2.045 116.445 2.305 ;
      RECT 116.145 2.092 116.445 2.288 ;
      RECT 116.136 2.1 116.145 2.291 ;
      RECT 115.73 2.193 116.445 2.288 ;
      RECT 116.05 2.118 116.136 2.298 ;
      RECT 115.745 2.19 116.445 2.288 ;
      RECT 115.991 2.14 116.05 2.31 ;
      RECT 115.765 2.186 116.445 2.288 ;
      RECT 115.905 2.152 115.991 2.321 ;
      RECT 115.78 2.182 116.445 2.288 ;
      RECT 115.85 2.165 115.905 2.333 ;
      RECT 115.795 2.18 116.445 2.288 ;
      RECT 115.835 2.171 115.85 2.339 ;
      RECT 115.805 2.176 116.445 2.288 ;
      RECT 115.95 1.7 116.21 1.96 ;
      RECT 115.95 1.72 116.32 1.93 ;
      RECT 115.95 1.725 116.33 1.925 ;
      RECT 116.141 1.139 116.22 1.37 ;
      RECT 116.055 1.142 116.27 1.365 ;
      RECT 116.05 1.142 116.27 1.36 ;
      RECT 116.05 1.147 116.28 1.358 ;
      RECT 116.025 1.147 116.28 1.355 ;
      RECT 116.025 1.155 116.29 1.353 ;
      RECT 115.905 1.09 116.165 1.35 ;
      RECT 115.905 1.137 116.215 1.35 ;
      RECT 115.16 1.71 115.165 1.97 ;
      RECT 114.99 1.48 114.995 1.97 ;
      RECT 114.875 1.72 114.88 1.945 ;
      RECT 115.585 0.815 115.59 1.025 ;
      RECT 115.59 0.82 115.605 1.02 ;
      RECT 115.525 0.815 115.585 1.033 ;
      RECT 115.51 0.815 115.525 1.043 ;
      RECT 115.46 0.815 115.51 1.06 ;
      RECT 115.44 0.815 115.46 1.083 ;
      RECT 115.425 0.815 115.44 1.095 ;
      RECT 115.405 0.815 115.425 1.105 ;
      RECT 115.395 0.82 115.405 1.114 ;
      RECT 115.39 0.83 115.395 1.119 ;
      RECT 115.385 0.842 115.39 1.123 ;
      RECT 115.375 0.865 115.385 1.128 ;
      RECT 115.37 0.88 115.375 1.132 ;
      RECT 115.365 0.897 115.37 1.135 ;
      RECT 115.36 0.905 115.365 1.138 ;
      RECT 115.35 0.91 115.36 1.142 ;
      RECT 115.345 0.917 115.35 1.147 ;
      RECT 115.335 0.922 115.345 1.151 ;
      RECT 115.31 0.934 115.335 1.162 ;
      RECT 115.29 0.951 115.31 1.178 ;
      RECT 115.265 0.968 115.29 1.2 ;
      RECT 115.23 0.991 115.265 1.258 ;
      RECT 115.21 1.013 115.23 1.32 ;
      RECT 115.205 1.023 115.21 1.355 ;
      RECT 115.195 1.03 115.205 1.393 ;
      RECT 115.19 1.037 115.195 1.413 ;
      RECT 115.185 1.048 115.19 1.45 ;
      RECT 115.18 1.056 115.185 1.515 ;
      RECT 115.17 1.067 115.18 1.568 ;
      RECT 115.165 1.085 115.17 1.638 ;
      RECT 115.16 1.095 115.165 1.675 ;
      RECT 115.155 1.105 115.16 1.97 ;
      RECT 115.15 1.117 115.155 1.97 ;
      RECT 115.145 1.127 115.15 1.97 ;
      RECT 115.135 1.137 115.145 1.97 ;
      RECT 115.125 1.16 115.135 1.97 ;
      RECT 115.11 1.195 115.125 1.97 ;
      RECT 115.07 1.257 115.11 1.97 ;
      RECT 115.065 1.31 115.07 1.97 ;
      RECT 115.04 1.345 115.065 1.97 ;
      RECT 115.025 1.39 115.04 1.97 ;
      RECT 115.02 1.412 115.025 1.97 ;
      RECT 115.01 1.425 115.02 1.97 ;
      RECT 115 1.45 115.01 1.97 ;
      RECT 114.995 1.472 115 1.97 ;
      RECT 114.97 1.51 114.99 1.97 ;
      RECT 114.93 1.567 114.97 1.97 ;
      RECT 114.925 1.617 114.93 1.97 ;
      RECT 114.92 1.635 114.925 1.97 ;
      RECT 114.915 1.647 114.92 1.97 ;
      RECT 114.905 1.665 114.915 1.97 ;
      RECT 114.895 1.685 114.905 1.945 ;
      RECT 114.89 1.702 114.895 1.945 ;
      RECT 114.88 1.715 114.89 1.945 ;
      RECT 114.85 1.725 114.875 1.945 ;
      RECT 114.84 1.732 114.85 1.945 ;
      RECT 114.825 1.742 114.84 1.94 ;
      RECT 113.785 1.655 114.105 1.915 ;
      RECT 113.65 1.7 114.105 1.87 ;
      RECT 107.12 1.515 107.495 1.765 ;
      RECT 107.22 0.73 107.395 1.765 ;
      RECT 112.93 0.715 113.25 0.975 ;
      RECT 112.93 0.745 113.33 0.915 ;
      RECT 107.22 0.73 113.25 0.905 ;
      RECT 110.595 1.755 110.89 2.045 ;
      RECT 110.565 1.755 110.89 2.015 ;
      RECT 96.805 2.125 97.11 2.355 ;
      RECT 104.945 2.155 108.36 2.33 ;
      RECT 108.185 1.305 108.36 2.33 ;
      RECT 96.805 2.155 108.36 2.325 ;
      RECT 108.13 1.305 108.46 1.555 ;
      RECT 105.39 1.315 105.68 1.555 ;
      RECT 100.94 1.285 101.2 1.52 ;
      RECT 100.94 1.315 105.68 1.485 ;
      RECT 104.125 1.655 104.445 1.915 ;
      RECT 104.11 1.7 104.445 1.87 ;
      RECT 102.83 0.635 103.125 0.925 ;
      RECT 102.795 0.635 103.125 0.895 ;
      RECT 99.99 1.655 100.31 1.915 ;
      RECT 99.975 1.7 100.31 1.87 ;
      RECT 98.315 1.445 98.635 1.705 ;
      RECT 98.3 1.445 98.655 1.68 ;
      RECT 95.615 1.205 95.8 1.415 ;
      RECT 95.605 1.21 95.815 1.408 ;
      RECT 95.605 1.21 95.901 1.385 ;
      RECT 95.605 1.21 95.96 1.36 ;
      RECT 95.605 1.21 96.015 1.34 ;
      RECT 95.605 1.21 96.025 1.328 ;
      RECT 95.605 1.21 96.22 1.267 ;
      RECT 95.605 1.21 96.25 1.25 ;
      RECT 95.605 1.21 96.27 1.24 ;
      RECT 96.15 0.975 96.41 1.235 ;
      RECT 96.135 1.065 96.15 1.282 ;
      RECT 95.67 1.197 96.41 1.235 ;
      RECT 96.121 1.076 96.135 1.288 ;
      RECT 95.71 1.19 96.41 1.235 ;
      RECT 96.035 1.116 96.121 1.307 ;
      RECT 95.96 1.177 96.41 1.235 ;
      RECT 96.03 1.152 96.035 1.324 ;
      RECT 96.015 1.162 96.41 1.235 ;
      RECT 96.025 1.157 96.03 1.326 ;
      RECT 96.32 1.662 96.325 1.754 ;
      RECT 96.315 1.64 96.32 1.771 ;
      RECT 96.31 1.63 96.315 1.783 ;
      RECT 96.3 1.621 96.31 1.793 ;
      RECT 96.295 1.616 96.3 1.801 ;
      RECT 96.29 1.612 96.295 1.804 ;
      RECT 96.256 1.545 96.29 1.815 ;
      RECT 96.17 1.545 96.256 1.85 ;
      RECT 96.09 1.545 96.17 1.898 ;
      RECT 96.03 1.545 96.09 1.923 ;
      RECT 95.97 1.645 96.03 1.93 ;
      RECT 95.935 1.67 95.97 1.936 ;
      RECT 95.91 1.685 95.935 1.94 ;
      RECT 95.896 1.694 95.91 1.942 ;
      RECT 95.81 1.721 95.896 1.948 ;
      RECT 95.745 1.762 95.81 1.957 ;
      RECT 95.73 1.782 95.745 1.962 ;
      RECT 95.7 1.792 95.73 1.965 ;
      RECT 95.695 1.802 95.7 1.968 ;
      RECT 95.665 1.807 95.695 1.97 ;
      RECT 95.645 1.812 95.665 1.974 ;
      RECT 95.56 1.815 95.645 1.981 ;
      RECT 95.545 1.812 95.56 1.987 ;
      RECT 95.535 1.809 95.545 1.989 ;
      RECT 95.515 1.806 95.535 1.991 ;
      RECT 95.495 1.802 95.515 1.992 ;
      RECT 95.48 1.798 95.495 1.994 ;
      RECT 95.47 1.795 95.48 1.995 ;
      RECT 95.43 1.789 95.47 1.993 ;
      RECT 95.42 1.784 95.43 1.991 ;
      RECT 95.405 1.781 95.42 1.987 ;
      RECT 95.38 1.776 95.405 1.98 ;
      RECT 95.33 1.767 95.38 1.968 ;
      RECT 95.26 1.753 95.33 1.95 ;
      RECT 95.202 1.738 95.26 1.932 ;
      RECT 95.116 1.721 95.202 1.912 ;
      RECT 95.03 1.7 95.116 1.887 ;
      RECT 94.98 1.685 95.03 1.868 ;
      RECT 94.976 1.679 94.98 1.86 ;
      RECT 94.89 1.669 94.976 1.847 ;
      RECT 94.855 1.654 94.89 1.83 ;
      RECT 94.84 1.647 94.855 1.823 ;
      RECT 94.78 1.635 94.84 1.811 ;
      RECT 94.76 1.622 94.78 1.799 ;
      RECT 94.72 1.613 94.76 1.791 ;
      RECT 94.715 1.605 94.72 1.784 ;
      RECT 94.635 1.595 94.715 1.77 ;
      RECT 94.62 1.582 94.635 1.755 ;
      RECT 94.615 1.58 94.62 1.753 ;
      RECT 94.536 1.568 94.615 1.74 ;
      RECT 94.45 1.543 94.536 1.715 ;
      RECT 94.435 1.512 94.45 1.7 ;
      RECT 94.42 1.487 94.435 1.696 ;
      RECT 94.405 1.48 94.42 1.692 ;
      RECT 94.23 1.485 94.235 1.688 ;
      RECT 94.225 1.49 94.23 1.683 ;
      RECT 94.235 1.48 94.405 1.69 ;
      RECT 94.95 1.24 95.055 1.5 ;
      RECT 95.765 0.765 95.77 0.99 ;
      RECT 95.895 0.765 95.95 0.975 ;
      RECT 95.95 0.77 95.96 0.968 ;
      RECT 95.856 0.765 95.895 0.978 ;
      RECT 95.77 0.765 95.856 0.985 ;
      RECT 95.75 0.77 95.765 0.991 ;
      RECT 95.74 0.81 95.75 0.993 ;
      RECT 95.71 0.82 95.74 0.995 ;
      RECT 95.705 0.825 95.71 0.997 ;
      RECT 95.68 0.83 95.705 0.999 ;
      RECT 95.665 0.835 95.68 1.001 ;
      RECT 95.65 0.837 95.665 1.003 ;
      RECT 95.645 0.842 95.65 1.005 ;
      RECT 95.595 0.85 95.645 1.008 ;
      RECT 95.57 0.859 95.595 1.013 ;
      RECT 95.56 0.866 95.57 1.018 ;
      RECT 95.555 0.869 95.56 1.022 ;
      RECT 95.535 0.872 95.555 1.031 ;
      RECT 95.505 0.88 95.535 1.051 ;
      RECT 95.476 0.893 95.505 1.073 ;
      RECT 95.39 0.927 95.476 1.117 ;
      RECT 95.385 0.953 95.39 1.155 ;
      RECT 95.38 0.957 95.385 1.164 ;
      RECT 95.345 0.97 95.38 1.197 ;
      RECT 95.335 0.984 95.345 1.235 ;
      RECT 95.33 0.988 95.335 1.248 ;
      RECT 95.325 0.992 95.33 1.253 ;
      RECT 95.315 1 95.325 1.265 ;
      RECT 95.31 1.007 95.315 1.28 ;
      RECT 95.285 1.02 95.31 1.305 ;
      RECT 95.245 1.049 95.285 1.36 ;
      RECT 95.23 1.074 95.245 1.415 ;
      RECT 95.22 1.085 95.23 1.438 ;
      RECT 95.215 1.092 95.22 1.45 ;
      RECT 95.21 1.096 95.215 1.458 ;
      RECT 95.155 1.124 95.21 1.5 ;
      RECT 95.135 1.16 95.155 1.5 ;
      RECT 95.12 1.175 95.135 1.5 ;
      RECT 95.065 1.207 95.12 1.5 ;
      RECT 95.055 1.237 95.065 1.5 ;
      RECT 94.665 0.852 94.85 1.09 ;
      RECT 94.65 0.854 94.86 1.085 ;
      RECT 94.535 0.8 94.795 1.06 ;
      RECT 94.53 0.837 94.795 1.014 ;
      RECT 94.525 0.847 94.795 1.011 ;
      RECT 94.52 0.887 94.86 1.005 ;
      RECT 94.515 0.92 94.86 0.995 ;
      RECT 94.525 0.862 94.875 0.933 ;
      RECT 94.822 1.96 94.835 2.49 ;
      RECT 94.736 1.96 94.835 2.489 ;
      RECT 94.736 1.96 94.84 2.488 ;
      RECT 94.65 1.96 94.84 2.486 ;
      RECT 94.645 1.96 94.84 2.483 ;
      RECT 94.645 1.96 94.85 2.481 ;
      RECT 94.64 2.252 94.85 2.478 ;
      RECT 94.64 2.262 94.855 2.475 ;
      RECT 94.64 2.33 94.86 2.471 ;
      RECT 94.63 2.335 94.86 2.47 ;
      RECT 94.63 2.427 94.865 2.467 ;
      RECT 94.615 1.96 94.875 2.22 ;
      RECT 93.845 0.95 93.89 2.485 ;
      RECT 94.045 0.95 94.075 1.165 ;
      RECT 92.42 0.69 92.54 0.9 ;
      RECT 92.08 0.64 92.34 0.9 ;
      RECT 92.08 0.685 92.375 0.89 ;
      RECT 94.085 0.966 94.09 1.02 ;
      RECT 94.08 0.959 94.085 1.153 ;
      RECT 94.075 0.953 94.08 1.16 ;
      RECT 94.03 0.95 94.045 1.173 ;
      RECT 94.025 0.95 94.03 1.195 ;
      RECT 94.02 0.95 94.025 1.243 ;
      RECT 94.015 0.95 94.02 1.263 ;
      RECT 94.005 0.95 94.015 1.37 ;
      RECT 94 0.95 94.005 1.433 ;
      RECT 93.995 0.95 94 1.49 ;
      RECT 93.99 0.95 93.995 1.498 ;
      RECT 93.975 0.95 93.99 1.605 ;
      RECT 93.965 0.95 93.975 1.74 ;
      RECT 93.955 0.95 93.965 1.85 ;
      RECT 93.945 0.95 93.955 1.907 ;
      RECT 93.94 0.95 93.945 1.947 ;
      RECT 93.935 0.95 93.94 1.983 ;
      RECT 93.925 0.95 93.935 2.023 ;
      RECT 93.92 0.95 93.925 2.065 ;
      RECT 93.9 0.95 93.92 2.13 ;
      RECT 93.905 2.275 93.91 2.455 ;
      RECT 93.9 2.257 93.905 2.463 ;
      RECT 93.895 0.95 93.9 2.193 ;
      RECT 93.895 2.237 93.9 2.47 ;
      RECT 93.89 0.95 93.895 2.48 ;
      RECT 93.835 0.95 93.845 1.25 ;
      RECT 93.84 1.497 93.845 2.485 ;
      RECT 93.835 1.562 93.84 2.485 ;
      RECT 93.83 0.951 93.835 1.24 ;
      RECT 93.825 1.627 93.835 2.485 ;
      RECT 93.82 0.952 93.83 1.23 ;
      RECT 93.81 1.74 93.825 2.485 ;
      RECT 93.815 0.953 93.82 1.22 ;
      RECT 93.795 0.954 93.815 1.198 ;
      RECT 93.8 1.837 93.81 2.485 ;
      RECT 93.795 1.912 93.8 2.485 ;
      RECT 93.785 0.953 93.795 1.175 ;
      RECT 93.79 1.955 93.795 2.485 ;
      RECT 93.785 1.982 93.79 2.485 ;
      RECT 93.775 0.951 93.785 1.163 ;
      RECT 93.78 2.025 93.785 2.485 ;
      RECT 93.775 2.052 93.78 2.485 ;
      RECT 93.765 0.95 93.775 1.15 ;
      RECT 93.77 2.067 93.775 2.485 ;
      RECT 93.73 2.125 93.77 2.485 ;
      RECT 93.76 0.949 93.765 1.135 ;
      RECT 93.755 0.947 93.76 1.128 ;
      RECT 93.745 0.944 93.755 1.118 ;
      RECT 93.74 0.941 93.745 1.103 ;
      RECT 93.725 0.937 93.74 1.096 ;
      RECT 93.72 2.18 93.73 2.485 ;
      RECT 93.72 0.934 93.725 1.091 ;
      RECT 93.705 0.93 93.72 1.085 ;
      RECT 93.715 2.197 93.72 2.485 ;
      RECT 93.705 2.26 93.715 2.485 ;
      RECT 93.625 0.915 93.705 1.065 ;
      RECT 93.7 2.267 93.705 2.48 ;
      RECT 93.695 2.275 93.7 2.47 ;
      RECT 93.615 0.901 93.625 1.049 ;
      RECT 93.6 0.897 93.615 1.047 ;
      RECT 93.59 0.892 93.6 1.043 ;
      RECT 93.565 0.885 93.59 1.035 ;
      RECT 93.56 0.88 93.565 1.03 ;
      RECT 93.55 0.88 93.56 1.028 ;
      RECT 93.54 0.878 93.55 1.026 ;
      RECT 93.51 0.87 93.54 1.02 ;
      RECT 93.495 0.862 93.51 1.013 ;
      RECT 93.475 0.857 93.495 1.006 ;
      RECT 93.47 0.853 93.475 1.001 ;
      RECT 93.44 0.846 93.47 0.995 ;
      RECT 93.415 0.837 93.44 0.985 ;
      RECT 93.385 0.83 93.415 0.977 ;
      RECT 93.36 0.82 93.385 0.968 ;
      RECT 93.345 0.812 93.36 0.962 ;
      RECT 93.32 0.807 93.345 0.957 ;
      RECT 93.31 0.803 93.32 0.952 ;
      RECT 93.29 0.798 93.31 0.947 ;
      RECT 93.255 0.793 93.29 0.94 ;
      RECT 93.195 0.788 93.255 0.933 ;
      RECT 93.182 0.784 93.195 0.931 ;
      RECT 93.096 0.779 93.182 0.928 ;
      RECT 93.01 0.769 93.096 0.924 ;
      RECT 92.969 0.762 93.01 0.921 ;
      RECT 92.883 0.755 92.969 0.918 ;
      RECT 92.797 0.745 92.883 0.914 ;
      RECT 92.711 0.735 92.797 0.909 ;
      RECT 92.625 0.725 92.711 0.905 ;
      RECT 92.615 0.71 92.625 0.903 ;
      RECT 92.605 0.695 92.615 0.903 ;
      RECT 92.54 0.69 92.605 0.902 ;
      RECT 92.375 0.687 92.42 0.895 ;
      RECT 93.62 1.592 93.625 1.783 ;
      RECT 93.615 1.587 93.62 1.79 ;
      RECT 93.601 1.585 93.615 1.796 ;
      RECT 93.515 1.585 93.601 1.798 ;
      RECT 93.511 1.585 93.515 1.801 ;
      RECT 93.425 1.585 93.511 1.819 ;
      RECT 93.415 1.59 93.425 1.838 ;
      RECT 93.405 1.645 93.415 1.842 ;
      RECT 93.38 1.66 93.405 1.849 ;
      RECT 93.34 1.68 93.38 1.862 ;
      RECT 93.335 1.692 93.34 1.872 ;
      RECT 93.32 1.698 93.335 1.877 ;
      RECT 93.315 1.703 93.32 1.881 ;
      RECT 93.295 1.71 93.315 1.886 ;
      RECT 93.225 1.735 93.295 1.903 ;
      RECT 93.185 1.763 93.225 1.923 ;
      RECT 93.18 1.773 93.185 1.931 ;
      RECT 93.16 1.78 93.18 1.933 ;
      RECT 93.155 1.787 93.16 1.936 ;
      RECT 93.125 1.795 93.155 1.939 ;
      RECT 93.12 1.8 93.125 1.943 ;
      RECT 93.046 1.804 93.12 1.951 ;
      RECT 92.96 1.813 93.046 1.967 ;
      RECT 92.956 1.818 92.96 1.976 ;
      RECT 92.87 1.823 92.956 1.986 ;
      RECT 92.83 1.831 92.87 1.998 ;
      RECT 92.78 1.837 92.83 2.005 ;
      RECT 92.695 1.846 92.78 2.02 ;
      RECT 92.62 1.857 92.695 2.038 ;
      RECT 92.585 1.864 92.62 2.048 ;
      RECT 92.51 1.872 92.585 2.053 ;
      RECT 92.455 1.881 92.51 2.053 ;
      RECT 92.43 1.886 92.455 2.051 ;
      RECT 92.42 1.889 92.43 2.049 ;
      RECT 92.385 1.891 92.42 2.047 ;
      RECT 92.355 1.893 92.385 2.043 ;
      RECT 92.31 1.892 92.355 2.039 ;
      RECT 92.29 1.887 92.31 2.036 ;
      RECT 92.24 1.872 92.29 2.033 ;
      RECT 92.23 1.857 92.24 2.028 ;
      RECT 92.18 1.842 92.23 2.018 ;
      RECT 92.13 1.817 92.18 1.998 ;
      RECT 92.12 1.802 92.13 1.98 ;
      RECT 92.115 1.8 92.12 1.974 ;
      RECT 92.095 1.795 92.115 1.969 ;
      RECT 92.09 1.787 92.095 1.963 ;
      RECT 92.075 1.781 92.09 1.956 ;
      RECT 92.07 1.776 92.075 1.948 ;
      RECT 92.05 1.771 92.07 1.94 ;
      RECT 92.035 1.764 92.05 1.933 ;
      RECT 92.02 1.758 92.035 1.924 ;
      RECT 92.015 1.752 92.02 1.917 ;
      RECT 91.97 1.727 92.015 1.903 ;
      RECT 91.955 1.697 91.97 1.885 ;
      RECT 91.94 1.68 91.955 1.876 ;
      RECT 91.915 1.66 91.94 1.864 ;
      RECT 91.875 1.63 91.915 1.844 ;
      RECT 91.865 1.6 91.875 1.829 ;
      RECT 91.85 1.59 91.865 1.822 ;
      RECT 91.795 1.555 91.85 1.801 ;
      RECT 91.78 1.518 91.795 1.78 ;
      RECT 91.77 1.505 91.78 1.772 ;
      RECT 91.72 1.475 91.77 1.754 ;
      RECT 91.705 1.405 91.72 1.735 ;
      RECT 91.66 1.405 91.705 1.718 ;
      RECT 91.635 1.405 91.66 1.7 ;
      RECT 91.625 1.405 91.635 1.693 ;
      RECT 91.546 1.405 91.625 1.686 ;
      RECT 91.46 1.405 91.546 1.678 ;
      RECT 91.445 1.437 91.46 1.673 ;
      RECT 91.37 1.447 91.445 1.669 ;
      RECT 91.35 1.457 91.37 1.664 ;
      RECT 91.325 1.457 91.35 1.661 ;
      RECT 91.315 1.447 91.325 1.66 ;
      RECT 91.305 1.42 91.315 1.659 ;
      RECT 91.265 1.415 91.305 1.657 ;
      RECT 91.22 1.415 91.265 1.653 ;
      RECT 91.195 1.415 91.22 1.648 ;
      RECT 91.145 1.415 91.195 1.635 ;
      RECT 91.105 1.42 91.115 1.62 ;
      RECT 91.115 1.415 91.145 1.625 ;
      RECT 93.1 1.195 93.36 1.455 ;
      RECT 93.095 1.217 93.36 1.413 ;
      RECT 92.335 1.045 92.555 1.41 ;
      RECT 92.317 1.132 92.555 1.409 ;
      RECT 92.3 1.137 92.555 1.406 ;
      RECT 92.3 1.137 92.575 1.405 ;
      RECT 92.27 1.147 92.575 1.403 ;
      RECT 92.265 1.162 92.575 1.399 ;
      RECT 92.265 1.162 92.58 1.398 ;
      RECT 92.26 1.22 92.58 1.396 ;
      RECT 92.26 1.22 92.59 1.393 ;
      RECT 92.255 1.285 92.59 1.388 ;
      RECT 92.335 1.045 92.595 1.305 ;
      RECT 91.08 0.875 91.34 1.135 ;
      RECT 91.08 0.918 91.426 1.109 ;
      RECT 91.08 0.918 91.47 1.108 ;
      RECT 91.08 0.918 91.49 1.106 ;
      RECT 91.08 0.918 91.59 1.105 ;
      RECT 91.08 0.918 91.61 1.103 ;
      RECT 91.08 0.918 91.62 1.098 ;
      RECT 91.49 0.885 91.68 1.095 ;
      RECT 91.49 0.887 91.685 1.093 ;
      RECT 91.48 0.892 91.69 1.085 ;
      RECT 91.426 0.916 91.69 1.085 ;
      RECT 91.47 0.91 91.48 1.107 ;
      RECT 91.48 0.89 91.685 1.093 ;
      RECT 90.435 1.95 90.64 2.18 ;
      RECT 90.375 1.9 90.43 2.16 ;
      RECT 90.435 1.9 90.635 2.18 ;
      RECT 91.405 2.215 91.41 2.242 ;
      RECT 91.395 2.125 91.405 2.247 ;
      RECT 91.39 2.047 91.395 2.253 ;
      RECT 91.38 2.037 91.39 2.26 ;
      RECT 91.375 2.027 91.38 2.266 ;
      RECT 91.365 2.022 91.375 2.268 ;
      RECT 91.35 2.014 91.365 2.276 ;
      RECT 91.335 2.005 91.35 2.288 ;
      RECT 91.325 1.997 91.335 2.298 ;
      RECT 91.29 1.915 91.325 2.316 ;
      RECT 91.255 1.915 91.29 2.335 ;
      RECT 91.24 1.915 91.255 2.343 ;
      RECT 91.185 1.915 91.24 2.343 ;
      RECT 91.151 1.915 91.185 2.334 ;
      RECT 91.065 1.915 91.151 2.31 ;
      RECT 91.055 1.975 91.065 2.292 ;
      RECT 91.015 1.977 91.055 2.283 ;
      RECT 91.01 1.979 91.015 2.273 ;
      RECT 90.99 1.981 91.01 2.268 ;
      RECT 90.98 1.984 90.99 2.263 ;
      RECT 90.97 1.985 90.98 2.258 ;
      RECT 90.946 1.986 90.97 2.25 ;
      RECT 90.86 1.991 90.946 2.228 ;
      RECT 90.805 1.99 90.86 2.201 ;
      RECT 90.79 1.983 90.805 2.188 ;
      RECT 90.755 1.978 90.79 2.184 ;
      RECT 90.7 1.97 90.755 2.183 ;
      RECT 90.64 1.957 90.7 2.181 ;
      RECT 90.43 1.9 90.435 2.168 ;
      RECT 90.505 1.27 90.69 1.48 ;
      RECT 90.495 1.275 90.705 1.473 ;
      RECT 90.535 1.18 90.795 1.44 ;
      RECT 90.49 1.337 90.795 1.363 ;
      RECT 89.835 1.13 89.84 1.93 ;
      RECT 89.78 1.18 89.81 1.93 ;
      RECT 89.77 1.18 89.775 1.49 ;
      RECT 89.755 1.18 89.76 1.485 ;
      RECT 89.3 1.225 89.315 1.44 ;
      RECT 89.23 1.225 89.315 1.435 ;
      RECT 90.495 0.805 90.565 1.015 ;
      RECT 90.565 0.812 90.575 1.01 ;
      RECT 90.461 0.805 90.495 1.022 ;
      RECT 90.375 0.805 90.461 1.046 ;
      RECT 90.365 0.81 90.375 1.065 ;
      RECT 90.36 0.822 90.365 1.068 ;
      RECT 90.345 0.837 90.36 1.072 ;
      RECT 90.34 0.855 90.345 1.076 ;
      RECT 90.3 0.865 90.34 1.085 ;
      RECT 90.285 0.872 90.3 1.097 ;
      RECT 90.27 0.877 90.285 1.102 ;
      RECT 90.255 0.88 90.27 1.107 ;
      RECT 90.245 0.882 90.255 1.111 ;
      RECT 90.21 0.889 90.245 1.119 ;
      RECT 90.175 0.897 90.21 1.133 ;
      RECT 90.165 0.903 90.175 1.142 ;
      RECT 90.16 0.905 90.165 1.144 ;
      RECT 90.14 0.908 90.16 1.15 ;
      RECT 90.11 0.915 90.14 1.161 ;
      RECT 90.1 0.921 90.11 1.168 ;
      RECT 90.075 0.924 90.1 1.175 ;
      RECT 90.065 0.928 90.075 1.183 ;
      RECT 90.06 0.929 90.065 1.205 ;
      RECT 90.055 0.93 90.06 1.22 ;
      RECT 90.05 0.931 90.055 1.235 ;
      RECT 90.045 0.932 90.05 1.25 ;
      RECT 90.04 0.933 90.045 1.28 ;
      RECT 90.03 0.935 90.04 1.313 ;
      RECT 90.015 0.939 90.03 1.36 ;
      RECT 90.005 0.942 90.015 1.405 ;
      RECT 90 0.945 90.005 1.433 ;
      RECT 89.99 0.947 90 1.46 ;
      RECT 89.985 0.95 89.99 1.495 ;
      RECT 89.955 0.955 89.985 1.553 ;
      RECT 89.95 0.96 89.955 1.638 ;
      RECT 89.945 0.962 89.95 1.673 ;
      RECT 89.94 0.964 89.945 1.755 ;
      RECT 89.935 0.966 89.94 1.843 ;
      RECT 89.925 0.968 89.935 1.925 ;
      RECT 89.91 0.982 89.925 1.93 ;
      RECT 89.875 1.027 89.91 1.93 ;
      RECT 89.865 1.067 89.875 1.93 ;
      RECT 89.85 1.095 89.865 1.93 ;
      RECT 89.845 1.112 89.85 1.93 ;
      RECT 89.84 1.12 89.845 1.93 ;
      RECT 89.83 1.135 89.835 1.93 ;
      RECT 89.825 1.142 89.83 1.93 ;
      RECT 89.815 1.162 89.825 1.93 ;
      RECT 89.81 1.175 89.815 1.93 ;
      RECT 89.775 1.18 89.78 1.515 ;
      RECT 89.76 1.57 89.78 1.93 ;
      RECT 89.76 1.18 89.77 1.488 ;
      RECT 89.755 1.61 89.76 1.93 ;
      RECT 89.705 1.18 89.755 1.483 ;
      RECT 89.75 1.647 89.755 1.93 ;
      RECT 89.74 1.67 89.75 1.93 ;
      RECT 89.735 1.715 89.74 1.93 ;
      RECT 89.725 1.725 89.735 1.923 ;
      RECT 89.651 1.18 89.705 1.477 ;
      RECT 89.565 1.18 89.651 1.47 ;
      RECT 89.516 1.227 89.565 1.463 ;
      RECT 89.43 1.235 89.516 1.456 ;
      RECT 89.415 1.232 89.43 1.451 ;
      RECT 89.401 1.225 89.415 1.45 ;
      RECT 89.315 1.225 89.401 1.445 ;
      RECT 89.22 1.23 89.23 1.43 ;
      RECT 88.81 0.66 88.825 1.06 ;
      RECT 89.005 0.66 89.01 0.92 ;
      RECT 88.75 0.66 88.795 0.92 ;
      RECT 89.205 1.965 89.21 2.17 ;
      RECT 89.2 1.955 89.205 2.175 ;
      RECT 89.195 1.942 89.2 2.18 ;
      RECT 89.19 1.922 89.195 2.18 ;
      RECT 89.165 1.875 89.19 2.18 ;
      RECT 89.13 1.79 89.165 2.18 ;
      RECT 89.125 1.727 89.13 2.18 ;
      RECT 89.12 1.712 89.125 2.18 ;
      RECT 89.105 1.672 89.12 2.18 ;
      RECT 89.1 1.647 89.105 2.18 ;
      RECT 89.09 1.63 89.1 2.18 ;
      RECT 89.055 1.552 89.09 2.18 ;
      RECT 89.05 1.495 89.055 2.18 ;
      RECT 89.045 1.482 89.05 2.18 ;
      RECT 89.035 1.46 89.045 2.18 ;
      RECT 89.025 1.425 89.035 2.18 ;
      RECT 89.015 1.395 89.025 2.18 ;
      RECT 89.005 1.31 89.015 1.823 ;
      RECT 89.012 1.955 89.015 2.18 ;
      RECT 89.01 1.965 89.012 2.18 ;
      RECT 89 1.975 89.01 2.175 ;
      RECT 88.995 0.66 89.005 1.055 ;
      RECT 89 1.187 89.005 1.798 ;
      RECT 88.995 1.085 89 1.781 ;
      RECT 88.985 0.66 88.995 1.757 ;
      RECT 88.98 0.66 88.985 1.728 ;
      RECT 88.975 0.66 88.98 1.718 ;
      RECT 88.955 0.66 88.975 1.68 ;
      RECT 88.95 0.66 88.955 1.638 ;
      RECT 88.945 0.66 88.95 1.618 ;
      RECT 88.915 0.66 88.945 1.568 ;
      RECT 88.905 0.66 88.915 1.515 ;
      RECT 88.9 0.66 88.905 1.488 ;
      RECT 88.895 0.66 88.9 1.473 ;
      RECT 88.885 0.66 88.895 1.45 ;
      RECT 88.875 0.66 88.885 1.425 ;
      RECT 88.87 0.66 88.875 1.365 ;
      RECT 88.86 0.66 88.87 1.303 ;
      RECT 88.855 0.66 88.86 1.223 ;
      RECT 88.85 0.66 88.855 1.188 ;
      RECT 88.845 0.66 88.85 1.163 ;
      RECT 88.84 0.66 88.845 1.148 ;
      RECT 88.835 0.66 88.84 1.118 ;
      RECT 88.83 0.66 88.835 1.095 ;
      RECT 88.825 0.66 88.83 1.068 ;
      RECT 88.795 0.66 88.81 1.055 ;
      RECT 87.95 2.195 88.135 2.405 ;
      RECT 87.94 2.2 88.15 2.398 ;
      RECT 87.94 2.2 88.17 2.37 ;
      RECT 87.94 2.2 88.185 2.349 ;
      RECT 87.94 2.2 88.2 2.347 ;
      RECT 87.94 2.2 88.21 2.346 ;
      RECT 87.94 2.2 88.24 2.343 ;
      RECT 88.59 2.045 88.85 2.305 ;
      RECT 88.55 2.092 88.85 2.288 ;
      RECT 88.541 2.1 88.55 2.291 ;
      RECT 88.135 2.193 88.85 2.288 ;
      RECT 88.455 2.118 88.541 2.298 ;
      RECT 88.15 2.19 88.85 2.288 ;
      RECT 88.396 2.14 88.455 2.31 ;
      RECT 88.17 2.186 88.85 2.288 ;
      RECT 88.31 2.152 88.396 2.321 ;
      RECT 88.185 2.182 88.85 2.288 ;
      RECT 88.255 2.165 88.31 2.333 ;
      RECT 88.2 2.18 88.85 2.288 ;
      RECT 88.24 2.171 88.255 2.339 ;
      RECT 88.21 2.176 88.85 2.288 ;
      RECT 88.355 1.7 88.615 1.96 ;
      RECT 88.355 1.72 88.725 1.93 ;
      RECT 88.355 1.725 88.735 1.925 ;
      RECT 88.546 1.139 88.625 1.37 ;
      RECT 88.46 1.142 88.675 1.365 ;
      RECT 88.455 1.142 88.675 1.36 ;
      RECT 88.455 1.147 88.685 1.358 ;
      RECT 88.43 1.147 88.685 1.355 ;
      RECT 88.43 1.155 88.695 1.353 ;
      RECT 88.31 1.09 88.57 1.35 ;
      RECT 88.31 1.137 88.62 1.35 ;
      RECT 87.565 1.71 87.57 1.97 ;
      RECT 87.395 1.48 87.4 1.97 ;
      RECT 87.28 1.72 87.285 1.945 ;
      RECT 87.99 0.815 87.995 1.025 ;
      RECT 87.995 0.82 88.01 1.02 ;
      RECT 87.93 0.815 87.99 1.033 ;
      RECT 87.915 0.815 87.93 1.043 ;
      RECT 87.865 0.815 87.915 1.06 ;
      RECT 87.845 0.815 87.865 1.083 ;
      RECT 87.83 0.815 87.845 1.095 ;
      RECT 87.81 0.815 87.83 1.105 ;
      RECT 87.8 0.82 87.81 1.114 ;
      RECT 87.795 0.83 87.8 1.119 ;
      RECT 87.79 0.842 87.795 1.123 ;
      RECT 87.78 0.865 87.79 1.128 ;
      RECT 87.775 0.88 87.78 1.132 ;
      RECT 87.77 0.897 87.775 1.135 ;
      RECT 87.765 0.905 87.77 1.138 ;
      RECT 87.755 0.91 87.765 1.142 ;
      RECT 87.75 0.917 87.755 1.147 ;
      RECT 87.74 0.922 87.75 1.151 ;
      RECT 87.715 0.934 87.74 1.162 ;
      RECT 87.695 0.951 87.715 1.178 ;
      RECT 87.67 0.968 87.695 1.2 ;
      RECT 87.635 0.991 87.67 1.258 ;
      RECT 87.615 1.013 87.635 1.32 ;
      RECT 87.61 1.023 87.615 1.355 ;
      RECT 87.6 1.03 87.61 1.393 ;
      RECT 87.595 1.037 87.6 1.413 ;
      RECT 87.59 1.048 87.595 1.45 ;
      RECT 87.585 1.056 87.59 1.515 ;
      RECT 87.575 1.067 87.585 1.568 ;
      RECT 87.57 1.085 87.575 1.638 ;
      RECT 87.565 1.095 87.57 1.675 ;
      RECT 87.56 1.105 87.565 1.97 ;
      RECT 87.555 1.117 87.56 1.97 ;
      RECT 87.55 1.127 87.555 1.97 ;
      RECT 87.54 1.137 87.55 1.97 ;
      RECT 87.53 1.16 87.54 1.97 ;
      RECT 87.515 1.195 87.53 1.97 ;
      RECT 87.475 1.257 87.515 1.97 ;
      RECT 87.47 1.31 87.475 1.97 ;
      RECT 87.445 1.345 87.47 1.97 ;
      RECT 87.43 1.39 87.445 1.97 ;
      RECT 87.425 1.412 87.43 1.97 ;
      RECT 87.415 1.425 87.425 1.97 ;
      RECT 87.405 1.45 87.415 1.97 ;
      RECT 87.4 1.472 87.405 1.97 ;
      RECT 87.375 1.51 87.395 1.97 ;
      RECT 87.335 1.567 87.375 1.97 ;
      RECT 87.33 1.617 87.335 1.97 ;
      RECT 87.325 1.635 87.33 1.97 ;
      RECT 87.32 1.647 87.325 1.97 ;
      RECT 87.31 1.665 87.32 1.97 ;
      RECT 87.3 1.685 87.31 1.945 ;
      RECT 87.295 1.702 87.3 1.945 ;
      RECT 87.285 1.715 87.295 1.945 ;
      RECT 87.255 1.725 87.28 1.945 ;
      RECT 87.245 1.732 87.255 1.945 ;
      RECT 87.23 1.742 87.245 1.94 ;
      RECT 86.19 1.655 86.51 1.915 ;
      RECT 86.055 1.7 86.51 1.87 ;
      RECT 79.54 1.515 79.915 1.765 ;
      RECT 79.64 0.73 79.815 1.765 ;
      RECT 85.335 0.715 85.655 0.975 ;
      RECT 85.335 0.745 85.735 0.915 ;
      RECT 79.64 0.73 85.655 0.905 ;
      RECT 83 1.755 83.295 2.045 ;
      RECT 82.97 1.755 83.295 2.015 ;
      RECT 69.21 2.125 69.515 2.355 ;
      RECT 77.35 2.155 80.765 2.33 ;
      RECT 80.59 1.305 80.765 2.33 ;
      RECT 69.21 2.155 80.765 2.325 ;
      RECT 80.535 1.305 80.865 1.555 ;
      RECT 77.795 1.315 78.085 1.555 ;
      RECT 73.345 1.285 73.605 1.52 ;
      RECT 73.345 1.315 78.085 1.485 ;
      RECT 76.53 1.655 76.85 1.915 ;
      RECT 76.515 1.7 76.85 1.87 ;
      RECT 75.235 0.635 75.53 0.925 ;
      RECT 75.2 0.635 75.53 0.895 ;
      RECT 72.395 1.655 72.715 1.915 ;
      RECT 72.38 1.7 72.715 1.87 ;
      RECT 70.72 1.445 71.04 1.705 ;
      RECT 70.705 1.445 71.06 1.68 ;
      RECT 68.02 1.205 68.205 1.415 ;
      RECT 68.01 1.21 68.22 1.408 ;
      RECT 68.01 1.21 68.306 1.385 ;
      RECT 68.01 1.21 68.365 1.36 ;
      RECT 68.01 1.21 68.42 1.34 ;
      RECT 68.01 1.21 68.43 1.328 ;
      RECT 68.01 1.21 68.625 1.267 ;
      RECT 68.01 1.21 68.655 1.25 ;
      RECT 68.01 1.21 68.675 1.24 ;
      RECT 68.555 0.975 68.815 1.235 ;
      RECT 68.54 1.065 68.555 1.282 ;
      RECT 68.075 1.197 68.815 1.235 ;
      RECT 68.526 1.076 68.54 1.288 ;
      RECT 68.115 1.19 68.815 1.235 ;
      RECT 68.44 1.116 68.526 1.307 ;
      RECT 68.365 1.177 68.815 1.235 ;
      RECT 68.435 1.152 68.44 1.324 ;
      RECT 68.42 1.162 68.815 1.235 ;
      RECT 68.43 1.157 68.435 1.326 ;
      RECT 68.725 1.662 68.73 1.754 ;
      RECT 68.72 1.64 68.725 1.771 ;
      RECT 68.715 1.63 68.72 1.783 ;
      RECT 68.705 1.621 68.715 1.793 ;
      RECT 68.7 1.616 68.705 1.801 ;
      RECT 68.695 1.612 68.7 1.804 ;
      RECT 68.661 1.545 68.695 1.815 ;
      RECT 68.575 1.545 68.661 1.85 ;
      RECT 68.495 1.545 68.575 1.898 ;
      RECT 68.435 1.545 68.495 1.923 ;
      RECT 68.375 1.645 68.435 1.93 ;
      RECT 68.34 1.67 68.375 1.936 ;
      RECT 68.315 1.685 68.34 1.94 ;
      RECT 68.301 1.694 68.315 1.942 ;
      RECT 68.215 1.721 68.301 1.948 ;
      RECT 68.15 1.762 68.215 1.957 ;
      RECT 68.135 1.782 68.15 1.962 ;
      RECT 68.105 1.792 68.135 1.965 ;
      RECT 68.1 1.802 68.105 1.968 ;
      RECT 68.07 1.807 68.1 1.97 ;
      RECT 68.05 1.812 68.07 1.974 ;
      RECT 67.965 1.815 68.05 1.981 ;
      RECT 67.95 1.812 67.965 1.987 ;
      RECT 67.94 1.809 67.95 1.989 ;
      RECT 67.92 1.806 67.94 1.991 ;
      RECT 67.9 1.802 67.92 1.992 ;
      RECT 67.885 1.798 67.9 1.994 ;
      RECT 67.875 1.795 67.885 1.995 ;
      RECT 67.835 1.789 67.875 1.993 ;
      RECT 67.825 1.784 67.835 1.991 ;
      RECT 67.81 1.781 67.825 1.987 ;
      RECT 67.785 1.776 67.81 1.98 ;
      RECT 67.735 1.767 67.785 1.968 ;
      RECT 67.665 1.753 67.735 1.95 ;
      RECT 67.607 1.738 67.665 1.932 ;
      RECT 67.521 1.721 67.607 1.912 ;
      RECT 67.435 1.7 67.521 1.887 ;
      RECT 67.385 1.685 67.435 1.868 ;
      RECT 67.381 1.679 67.385 1.86 ;
      RECT 67.295 1.669 67.381 1.847 ;
      RECT 67.26 1.654 67.295 1.83 ;
      RECT 67.245 1.647 67.26 1.823 ;
      RECT 67.185 1.635 67.245 1.811 ;
      RECT 67.165 1.622 67.185 1.799 ;
      RECT 67.125 1.613 67.165 1.791 ;
      RECT 67.12 1.605 67.125 1.784 ;
      RECT 67.04 1.595 67.12 1.77 ;
      RECT 67.025 1.582 67.04 1.755 ;
      RECT 67.02 1.58 67.025 1.753 ;
      RECT 66.941 1.568 67.02 1.74 ;
      RECT 66.855 1.543 66.941 1.715 ;
      RECT 66.84 1.512 66.855 1.7 ;
      RECT 66.825 1.487 66.84 1.696 ;
      RECT 66.81 1.48 66.825 1.692 ;
      RECT 66.635 1.485 66.64 1.688 ;
      RECT 66.63 1.49 66.635 1.683 ;
      RECT 66.64 1.48 66.81 1.69 ;
      RECT 67.355 1.24 67.46 1.5 ;
      RECT 68.17 0.765 68.175 0.99 ;
      RECT 68.3 0.765 68.355 0.975 ;
      RECT 68.355 0.77 68.365 0.968 ;
      RECT 68.261 0.765 68.3 0.978 ;
      RECT 68.175 0.765 68.261 0.985 ;
      RECT 68.155 0.77 68.17 0.991 ;
      RECT 68.145 0.81 68.155 0.993 ;
      RECT 68.115 0.82 68.145 0.995 ;
      RECT 68.11 0.825 68.115 0.997 ;
      RECT 68.085 0.83 68.11 0.999 ;
      RECT 68.07 0.835 68.085 1.001 ;
      RECT 68.055 0.837 68.07 1.003 ;
      RECT 68.05 0.842 68.055 1.005 ;
      RECT 68 0.85 68.05 1.008 ;
      RECT 67.975 0.859 68 1.013 ;
      RECT 67.965 0.866 67.975 1.018 ;
      RECT 67.96 0.869 67.965 1.022 ;
      RECT 67.94 0.872 67.96 1.031 ;
      RECT 67.91 0.88 67.94 1.051 ;
      RECT 67.881 0.893 67.91 1.073 ;
      RECT 67.795 0.927 67.881 1.117 ;
      RECT 67.79 0.953 67.795 1.155 ;
      RECT 67.785 0.957 67.79 1.164 ;
      RECT 67.75 0.97 67.785 1.197 ;
      RECT 67.74 0.984 67.75 1.235 ;
      RECT 67.735 0.988 67.74 1.248 ;
      RECT 67.73 0.992 67.735 1.253 ;
      RECT 67.72 1 67.73 1.265 ;
      RECT 67.715 1.007 67.72 1.28 ;
      RECT 67.69 1.02 67.715 1.305 ;
      RECT 67.65 1.049 67.69 1.36 ;
      RECT 67.635 1.074 67.65 1.415 ;
      RECT 67.625 1.085 67.635 1.438 ;
      RECT 67.62 1.092 67.625 1.45 ;
      RECT 67.615 1.096 67.62 1.458 ;
      RECT 67.56 1.124 67.615 1.5 ;
      RECT 67.54 1.16 67.56 1.5 ;
      RECT 67.525 1.175 67.54 1.5 ;
      RECT 67.47 1.207 67.525 1.5 ;
      RECT 67.46 1.237 67.47 1.5 ;
      RECT 67.07 0.852 67.255 1.09 ;
      RECT 67.055 0.854 67.265 1.085 ;
      RECT 66.94 0.8 67.2 1.06 ;
      RECT 66.935 0.837 67.2 1.014 ;
      RECT 66.93 0.847 67.2 1.011 ;
      RECT 66.925 0.887 67.265 1.005 ;
      RECT 66.92 0.92 67.265 0.995 ;
      RECT 66.93 0.862 67.28 0.933 ;
      RECT 67.227 1.96 67.24 2.49 ;
      RECT 67.141 1.96 67.24 2.489 ;
      RECT 67.141 1.96 67.245 2.488 ;
      RECT 67.055 1.96 67.245 2.486 ;
      RECT 67.05 1.96 67.245 2.483 ;
      RECT 67.05 1.96 67.255 2.481 ;
      RECT 67.045 2.252 67.255 2.478 ;
      RECT 67.045 2.262 67.26 2.475 ;
      RECT 67.045 2.33 67.265 2.471 ;
      RECT 67.035 2.335 67.265 2.47 ;
      RECT 67.035 2.427 67.27 2.467 ;
      RECT 67.02 1.96 67.28 2.22 ;
      RECT 66.25 0.95 66.295 2.485 ;
      RECT 66.45 0.95 66.48 1.165 ;
      RECT 64.825 0.69 64.945 0.9 ;
      RECT 64.485 0.64 64.745 0.9 ;
      RECT 64.485 0.685 64.78 0.89 ;
      RECT 66.49 0.966 66.495 1.02 ;
      RECT 66.485 0.959 66.49 1.153 ;
      RECT 66.48 0.953 66.485 1.16 ;
      RECT 66.435 0.95 66.45 1.173 ;
      RECT 66.43 0.95 66.435 1.195 ;
      RECT 66.425 0.95 66.43 1.243 ;
      RECT 66.42 0.95 66.425 1.263 ;
      RECT 66.41 0.95 66.42 1.37 ;
      RECT 66.405 0.95 66.41 1.433 ;
      RECT 66.4 0.95 66.405 1.49 ;
      RECT 66.395 0.95 66.4 1.498 ;
      RECT 66.38 0.95 66.395 1.605 ;
      RECT 66.37 0.95 66.38 1.74 ;
      RECT 66.36 0.95 66.37 1.85 ;
      RECT 66.35 0.95 66.36 1.907 ;
      RECT 66.345 0.95 66.35 1.947 ;
      RECT 66.34 0.95 66.345 1.983 ;
      RECT 66.33 0.95 66.34 2.023 ;
      RECT 66.325 0.95 66.33 2.065 ;
      RECT 66.305 0.95 66.325 2.13 ;
      RECT 66.31 2.275 66.315 2.455 ;
      RECT 66.305 2.257 66.31 2.463 ;
      RECT 66.3 0.95 66.305 2.193 ;
      RECT 66.3 2.237 66.305 2.47 ;
      RECT 66.295 0.95 66.3 2.48 ;
      RECT 66.24 0.95 66.25 1.25 ;
      RECT 66.245 1.497 66.25 2.485 ;
      RECT 66.24 1.562 66.245 2.485 ;
      RECT 66.235 0.951 66.24 1.24 ;
      RECT 66.23 1.627 66.24 2.485 ;
      RECT 66.225 0.952 66.235 1.23 ;
      RECT 66.215 1.74 66.23 2.485 ;
      RECT 66.22 0.953 66.225 1.22 ;
      RECT 66.2 0.954 66.22 1.198 ;
      RECT 66.205 1.837 66.215 2.485 ;
      RECT 66.2 1.912 66.205 2.485 ;
      RECT 66.19 0.953 66.2 1.175 ;
      RECT 66.195 1.955 66.2 2.485 ;
      RECT 66.19 1.982 66.195 2.485 ;
      RECT 66.18 0.951 66.19 1.163 ;
      RECT 66.185 2.025 66.19 2.485 ;
      RECT 66.18 2.052 66.185 2.485 ;
      RECT 66.17 0.95 66.18 1.15 ;
      RECT 66.175 2.067 66.18 2.485 ;
      RECT 66.135 2.125 66.175 2.485 ;
      RECT 66.165 0.949 66.17 1.135 ;
      RECT 66.16 0.947 66.165 1.128 ;
      RECT 66.15 0.944 66.16 1.118 ;
      RECT 66.145 0.941 66.15 1.103 ;
      RECT 66.13 0.937 66.145 1.096 ;
      RECT 66.125 2.18 66.135 2.485 ;
      RECT 66.125 0.934 66.13 1.091 ;
      RECT 66.11 0.93 66.125 1.085 ;
      RECT 66.12 2.197 66.125 2.485 ;
      RECT 66.11 2.26 66.12 2.485 ;
      RECT 66.03 0.915 66.11 1.065 ;
      RECT 66.105 2.267 66.11 2.48 ;
      RECT 66.1 2.275 66.105 2.47 ;
      RECT 66.02 0.901 66.03 1.049 ;
      RECT 66.005 0.897 66.02 1.047 ;
      RECT 65.995 0.892 66.005 1.043 ;
      RECT 65.97 0.885 65.995 1.035 ;
      RECT 65.965 0.88 65.97 1.03 ;
      RECT 65.955 0.88 65.965 1.028 ;
      RECT 65.945 0.878 65.955 1.026 ;
      RECT 65.915 0.87 65.945 1.02 ;
      RECT 65.9 0.862 65.915 1.013 ;
      RECT 65.88 0.857 65.9 1.006 ;
      RECT 65.875 0.853 65.88 1.001 ;
      RECT 65.845 0.846 65.875 0.995 ;
      RECT 65.82 0.837 65.845 0.985 ;
      RECT 65.79 0.83 65.82 0.977 ;
      RECT 65.765 0.82 65.79 0.968 ;
      RECT 65.75 0.812 65.765 0.962 ;
      RECT 65.725 0.807 65.75 0.957 ;
      RECT 65.715 0.803 65.725 0.952 ;
      RECT 65.695 0.798 65.715 0.947 ;
      RECT 65.66 0.793 65.695 0.94 ;
      RECT 65.6 0.788 65.66 0.933 ;
      RECT 65.587 0.784 65.6 0.931 ;
      RECT 65.501 0.779 65.587 0.928 ;
      RECT 65.415 0.769 65.501 0.924 ;
      RECT 65.374 0.762 65.415 0.921 ;
      RECT 65.288 0.755 65.374 0.918 ;
      RECT 65.202 0.745 65.288 0.914 ;
      RECT 65.116 0.735 65.202 0.909 ;
      RECT 65.03 0.725 65.116 0.905 ;
      RECT 65.02 0.71 65.03 0.903 ;
      RECT 65.01 0.695 65.02 0.903 ;
      RECT 64.945 0.69 65.01 0.902 ;
      RECT 64.78 0.687 64.825 0.895 ;
      RECT 66.025 1.592 66.03 1.783 ;
      RECT 66.02 1.587 66.025 1.79 ;
      RECT 66.006 1.585 66.02 1.796 ;
      RECT 65.92 1.585 66.006 1.798 ;
      RECT 65.916 1.585 65.92 1.801 ;
      RECT 65.83 1.585 65.916 1.819 ;
      RECT 65.82 1.59 65.83 1.838 ;
      RECT 65.81 1.645 65.82 1.842 ;
      RECT 65.785 1.66 65.81 1.849 ;
      RECT 65.745 1.68 65.785 1.862 ;
      RECT 65.74 1.692 65.745 1.872 ;
      RECT 65.725 1.698 65.74 1.877 ;
      RECT 65.72 1.703 65.725 1.881 ;
      RECT 65.7 1.71 65.72 1.886 ;
      RECT 65.63 1.735 65.7 1.903 ;
      RECT 65.59 1.763 65.63 1.923 ;
      RECT 65.585 1.773 65.59 1.931 ;
      RECT 65.565 1.78 65.585 1.933 ;
      RECT 65.56 1.787 65.565 1.936 ;
      RECT 65.53 1.795 65.56 1.939 ;
      RECT 65.525 1.8 65.53 1.943 ;
      RECT 65.451 1.804 65.525 1.951 ;
      RECT 65.365 1.813 65.451 1.967 ;
      RECT 65.361 1.818 65.365 1.976 ;
      RECT 65.275 1.823 65.361 1.986 ;
      RECT 65.235 1.831 65.275 1.998 ;
      RECT 65.185 1.837 65.235 2.005 ;
      RECT 65.1 1.846 65.185 2.02 ;
      RECT 65.025 1.857 65.1 2.038 ;
      RECT 64.99 1.864 65.025 2.048 ;
      RECT 64.915 1.872 64.99 2.053 ;
      RECT 64.86 1.881 64.915 2.053 ;
      RECT 64.835 1.886 64.86 2.051 ;
      RECT 64.825 1.889 64.835 2.049 ;
      RECT 64.79 1.891 64.825 2.047 ;
      RECT 64.76 1.893 64.79 2.043 ;
      RECT 64.715 1.892 64.76 2.039 ;
      RECT 64.695 1.887 64.715 2.036 ;
      RECT 64.645 1.872 64.695 2.033 ;
      RECT 64.635 1.857 64.645 2.028 ;
      RECT 64.585 1.842 64.635 2.018 ;
      RECT 64.535 1.817 64.585 1.998 ;
      RECT 64.525 1.802 64.535 1.98 ;
      RECT 64.52 1.8 64.525 1.974 ;
      RECT 64.5 1.795 64.52 1.969 ;
      RECT 64.495 1.787 64.5 1.963 ;
      RECT 64.48 1.781 64.495 1.956 ;
      RECT 64.475 1.776 64.48 1.948 ;
      RECT 64.455 1.771 64.475 1.94 ;
      RECT 64.44 1.764 64.455 1.933 ;
      RECT 64.425 1.758 64.44 1.924 ;
      RECT 64.42 1.752 64.425 1.917 ;
      RECT 64.375 1.727 64.42 1.903 ;
      RECT 64.36 1.697 64.375 1.885 ;
      RECT 64.345 1.68 64.36 1.876 ;
      RECT 64.32 1.66 64.345 1.864 ;
      RECT 64.28 1.63 64.32 1.844 ;
      RECT 64.27 1.6 64.28 1.829 ;
      RECT 64.255 1.59 64.27 1.822 ;
      RECT 64.2 1.555 64.255 1.801 ;
      RECT 64.185 1.518 64.2 1.78 ;
      RECT 64.175 1.505 64.185 1.772 ;
      RECT 64.125 1.475 64.175 1.754 ;
      RECT 64.11 1.405 64.125 1.735 ;
      RECT 64.065 1.405 64.11 1.718 ;
      RECT 64.04 1.405 64.065 1.7 ;
      RECT 64.03 1.405 64.04 1.693 ;
      RECT 63.951 1.405 64.03 1.686 ;
      RECT 63.865 1.405 63.951 1.678 ;
      RECT 63.85 1.437 63.865 1.673 ;
      RECT 63.775 1.447 63.85 1.669 ;
      RECT 63.755 1.457 63.775 1.664 ;
      RECT 63.73 1.457 63.755 1.661 ;
      RECT 63.72 1.447 63.73 1.66 ;
      RECT 63.71 1.42 63.72 1.659 ;
      RECT 63.67 1.415 63.71 1.657 ;
      RECT 63.625 1.415 63.67 1.653 ;
      RECT 63.6 1.415 63.625 1.648 ;
      RECT 63.55 1.415 63.6 1.635 ;
      RECT 63.51 1.42 63.52 1.62 ;
      RECT 63.52 1.415 63.55 1.625 ;
      RECT 65.505 1.195 65.765 1.455 ;
      RECT 65.5 1.217 65.765 1.413 ;
      RECT 64.74 1.045 64.96 1.41 ;
      RECT 64.722 1.132 64.96 1.409 ;
      RECT 64.705 1.137 64.96 1.406 ;
      RECT 64.705 1.137 64.98 1.405 ;
      RECT 64.675 1.147 64.98 1.403 ;
      RECT 64.67 1.162 64.98 1.399 ;
      RECT 64.67 1.162 64.985 1.398 ;
      RECT 64.665 1.22 64.985 1.396 ;
      RECT 64.665 1.22 64.995 1.393 ;
      RECT 64.66 1.285 64.995 1.388 ;
      RECT 64.74 1.045 65 1.305 ;
      RECT 63.485 0.875 63.745 1.135 ;
      RECT 63.485 0.918 63.831 1.109 ;
      RECT 63.485 0.918 63.875 1.108 ;
      RECT 63.485 0.918 63.895 1.106 ;
      RECT 63.485 0.918 63.995 1.105 ;
      RECT 63.485 0.918 64.015 1.103 ;
      RECT 63.485 0.918 64.025 1.098 ;
      RECT 63.895 0.885 64.085 1.095 ;
      RECT 63.895 0.887 64.09 1.093 ;
      RECT 63.885 0.892 64.095 1.085 ;
      RECT 63.831 0.916 64.095 1.085 ;
      RECT 63.875 0.91 63.885 1.107 ;
      RECT 63.885 0.89 64.09 1.093 ;
      RECT 62.84 1.95 63.045 2.18 ;
      RECT 62.78 1.9 62.835 2.16 ;
      RECT 62.84 1.9 63.04 2.18 ;
      RECT 63.81 2.215 63.815 2.242 ;
      RECT 63.8 2.125 63.81 2.247 ;
      RECT 63.795 2.047 63.8 2.253 ;
      RECT 63.785 2.037 63.795 2.26 ;
      RECT 63.78 2.027 63.785 2.266 ;
      RECT 63.77 2.022 63.78 2.268 ;
      RECT 63.755 2.014 63.77 2.276 ;
      RECT 63.74 2.005 63.755 2.288 ;
      RECT 63.73 1.997 63.74 2.298 ;
      RECT 63.695 1.915 63.73 2.316 ;
      RECT 63.66 1.915 63.695 2.335 ;
      RECT 63.645 1.915 63.66 2.343 ;
      RECT 63.59 1.915 63.645 2.343 ;
      RECT 63.556 1.915 63.59 2.334 ;
      RECT 63.47 1.915 63.556 2.31 ;
      RECT 63.46 1.975 63.47 2.292 ;
      RECT 63.42 1.977 63.46 2.283 ;
      RECT 63.415 1.979 63.42 2.273 ;
      RECT 63.395 1.981 63.415 2.268 ;
      RECT 63.385 1.984 63.395 2.263 ;
      RECT 63.375 1.985 63.385 2.258 ;
      RECT 63.351 1.986 63.375 2.25 ;
      RECT 63.265 1.991 63.351 2.228 ;
      RECT 63.21 1.99 63.265 2.201 ;
      RECT 63.195 1.983 63.21 2.188 ;
      RECT 63.16 1.978 63.195 2.184 ;
      RECT 63.105 1.97 63.16 2.183 ;
      RECT 63.045 1.957 63.105 2.181 ;
      RECT 62.835 1.9 62.84 2.168 ;
      RECT 62.91 1.27 63.095 1.48 ;
      RECT 62.9 1.275 63.11 1.473 ;
      RECT 62.94 1.18 63.2 1.44 ;
      RECT 62.895 1.337 63.2 1.363 ;
      RECT 62.24 1.13 62.245 1.93 ;
      RECT 62.185 1.18 62.215 1.93 ;
      RECT 62.175 1.18 62.18 1.49 ;
      RECT 62.16 1.18 62.165 1.485 ;
      RECT 61.705 1.225 61.72 1.44 ;
      RECT 61.635 1.225 61.72 1.435 ;
      RECT 62.9 0.805 62.97 1.015 ;
      RECT 62.97 0.812 62.98 1.01 ;
      RECT 62.866 0.805 62.9 1.022 ;
      RECT 62.78 0.805 62.866 1.046 ;
      RECT 62.77 0.81 62.78 1.065 ;
      RECT 62.765 0.822 62.77 1.068 ;
      RECT 62.75 0.837 62.765 1.072 ;
      RECT 62.745 0.855 62.75 1.076 ;
      RECT 62.705 0.865 62.745 1.085 ;
      RECT 62.69 0.872 62.705 1.097 ;
      RECT 62.675 0.877 62.69 1.102 ;
      RECT 62.66 0.88 62.675 1.107 ;
      RECT 62.65 0.882 62.66 1.111 ;
      RECT 62.615 0.889 62.65 1.119 ;
      RECT 62.58 0.897 62.615 1.133 ;
      RECT 62.57 0.903 62.58 1.142 ;
      RECT 62.565 0.905 62.57 1.144 ;
      RECT 62.545 0.908 62.565 1.15 ;
      RECT 62.515 0.915 62.545 1.161 ;
      RECT 62.505 0.921 62.515 1.168 ;
      RECT 62.48 0.924 62.505 1.175 ;
      RECT 62.47 0.928 62.48 1.183 ;
      RECT 62.465 0.929 62.47 1.205 ;
      RECT 62.46 0.93 62.465 1.22 ;
      RECT 62.455 0.931 62.46 1.235 ;
      RECT 62.45 0.932 62.455 1.25 ;
      RECT 62.445 0.933 62.45 1.28 ;
      RECT 62.435 0.935 62.445 1.313 ;
      RECT 62.42 0.939 62.435 1.36 ;
      RECT 62.41 0.942 62.42 1.405 ;
      RECT 62.405 0.945 62.41 1.433 ;
      RECT 62.395 0.947 62.405 1.46 ;
      RECT 62.39 0.95 62.395 1.495 ;
      RECT 62.36 0.955 62.39 1.553 ;
      RECT 62.355 0.96 62.36 1.638 ;
      RECT 62.35 0.962 62.355 1.673 ;
      RECT 62.345 0.964 62.35 1.755 ;
      RECT 62.34 0.966 62.345 1.843 ;
      RECT 62.33 0.968 62.34 1.925 ;
      RECT 62.315 0.982 62.33 1.93 ;
      RECT 62.28 1.027 62.315 1.93 ;
      RECT 62.27 1.067 62.28 1.93 ;
      RECT 62.255 1.095 62.27 1.93 ;
      RECT 62.25 1.112 62.255 1.93 ;
      RECT 62.245 1.12 62.25 1.93 ;
      RECT 62.235 1.135 62.24 1.93 ;
      RECT 62.23 1.142 62.235 1.93 ;
      RECT 62.22 1.162 62.23 1.93 ;
      RECT 62.215 1.175 62.22 1.93 ;
      RECT 62.18 1.18 62.185 1.515 ;
      RECT 62.165 1.57 62.185 1.93 ;
      RECT 62.165 1.18 62.175 1.488 ;
      RECT 62.16 1.61 62.165 1.93 ;
      RECT 62.11 1.18 62.16 1.483 ;
      RECT 62.155 1.647 62.16 1.93 ;
      RECT 62.145 1.67 62.155 1.93 ;
      RECT 62.14 1.715 62.145 1.93 ;
      RECT 62.13 1.725 62.14 1.923 ;
      RECT 62.056 1.18 62.11 1.477 ;
      RECT 61.97 1.18 62.056 1.47 ;
      RECT 61.921 1.227 61.97 1.463 ;
      RECT 61.835 1.235 61.921 1.456 ;
      RECT 61.82 1.232 61.835 1.451 ;
      RECT 61.806 1.225 61.82 1.45 ;
      RECT 61.72 1.225 61.806 1.445 ;
      RECT 61.625 1.23 61.635 1.43 ;
      RECT 61.215 0.66 61.23 1.06 ;
      RECT 61.41 0.66 61.415 0.92 ;
      RECT 61.155 0.66 61.2 0.92 ;
      RECT 61.61 1.965 61.615 2.17 ;
      RECT 61.605 1.955 61.61 2.175 ;
      RECT 61.6 1.942 61.605 2.18 ;
      RECT 61.595 1.922 61.6 2.18 ;
      RECT 61.57 1.875 61.595 2.18 ;
      RECT 61.535 1.79 61.57 2.18 ;
      RECT 61.53 1.727 61.535 2.18 ;
      RECT 61.525 1.712 61.53 2.18 ;
      RECT 61.51 1.672 61.525 2.18 ;
      RECT 61.505 1.647 61.51 2.18 ;
      RECT 61.495 1.63 61.505 2.18 ;
      RECT 61.46 1.552 61.495 2.18 ;
      RECT 61.455 1.495 61.46 2.18 ;
      RECT 61.45 1.482 61.455 2.18 ;
      RECT 61.44 1.46 61.45 2.18 ;
      RECT 61.43 1.425 61.44 2.18 ;
      RECT 61.42 1.395 61.43 2.18 ;
      RECT 61.41 1.31 61.42 1.823 ;
      RECT 61.417 1.955 61.42 2.18 ;
      RECT 61.415 1.965 61.417 2.18 ;
      RECT 61.405 1.975 61.415 2.175 ;
      RECT 61.4 0.66 61.41 1.055 ;
      RECT 61.405 1.187 61.41 1.798 ;
      RECT 61.4 1.085 61.405 1.781 ;
      RECT 61.39 0.66 61.4 1.757 ;
      RECT 61.385 0.66 61.39 1.728 ;
      RECT 61.38 0.66 61.385 1.718 ;
      RECT 61.36 0.66 61.38 1.68 ;
      RECT 61.355 0.66 61.36 1.638 ;
      RECT 61.35 0.66 61.355 1.618 ;
      RECT 61.32 0.66 61.35 1.568 ;
      RECT 61.31 0.66 61.32 1.515 ;
      RECT 61.305 0.66 61.31 1.488 ;
      RECT 61.3 0.66 61.305 1.473 ;
      RECT 61.29 0.66 61.3 1.45 ;
      RECT 61.28 0.66 61.29 1.425 ;
      RECT 61.275 0.66 61.28 1.365 ;
      RECT 61.265 0.66 61.275 1.303 ;
      RECT 61.26 0.66 61.265 1.223 ;
      RECT 61.255 0.66 61.26 1.188 ;
      RECT 61.25 0.66 61.255 1.163 ;
      RECT 61.245 0.66 61.25 1.148 ;
      RECT 61.24 0.66 61.245 1.118 ;
      RECT 61.235 0.66 61.24 1.095 ;
      RECT 61.23 0.66 61.235 1.068 ;
      RECT 61.2 0.66 61.215 1.055 ;
      RECT 60.355 2.195 60.54 2.405 ;
      RECT 60.345 2.2 60.555 2.398 ;
      RECT 60.345 2.2 60.575 2.37 ;
      RECT 60.345 2.2 60.59 2.349 ;
      RECT 60.345 2.2 60.605 2.347 ;
      RECT 60.345 2.2 60.615 2.346 ;
      RECT 60.345 2.2 60.645 2.343 ;
      RECT 60.995 2.045 61.255 2.305 ;
      RECT 60.955 2.092 61.255 2.288 ;
      RECT 60.946 2.1 60.955 2.291 ;
      RECT 60.54 2.193 61.255 2.288 ;
      RECT 60.86 2.118 60.946 2.298 ;
      RECT 60.555 2.19 61.255 2.288 ;
      RECT 60.801 2.14 60.86 2.31 ;
      RECT 60.575 2.186 61.255 2.288 ;
      RECT 60.715 2.152 60.801 2.321 ;
      RECT 60.59 2.182 61.255 2.288 ;
      RECT 60.66 2.165 60.715 2.333 ;
      RECT 60.605 2.18 61.255 2.288 ;
      RECT 60.645 2.171 60.66 2.339 ;
      RECT 60.615 2.176 61.255 2.288 ;
      RECT 60.76 1.7 61.02 1.96 ;
      RECT 60.76 1.72 61.13 1.93 ;
      RECT 60.76 1.725 61.14 1.925 ;
      RECT 60.951 1.139 61.03 1.37 ;
      RECT 60.865 1.142 61.08 1.365 ;
      RECT 60.86 1.142 61.08 1.36 ;
      RECT 60.86 1.147 61.09 1.358 ;
      RECT 60.835 1.147 61.09 1.355 ;
      RECT 60.835 1.155 61.1 1.353 ;
      RECT 60.715 1.09 60.975 1.35 ;
      RECT 60.715 1.137 61.025 1.35 ;
      RECT 59.97 1.71 59.975 1.97 ;
      RECT 59.8 1.48 59.805 1.97 ;
      RECT 59.685 1.72 59.69 1.945 ;
      RECT 60.395 0.815 60.4 1.025 ;
      RECT 60.4 0.82 60.415 1.02 ;
      RECT 60.335 0.815 60.395 1.033 ;
      RECT 60.32 0.815 60.335 1.043 ;
      RECT 60.27 0.815 60.32 1.06 ;
      RECT 60.25 0.815 60.27 1.083 ;
      RECT 60.235 0.815 60.25 1.095 ;
      RECT 60.215 0.815 60.235 1.105 ;
      RECT 60.205 0.82 60.215 1.114 ;
      RECT 60.2 0.83 60.205 1.119 ;
      RECT 60.195 0.842 60.2 1.123 ;
      RECT 60.185 0.865 60.195 1.128 ;
      RECT 60.18 0.88 60.185 1.132 ;
      RECT 60.175 0.897 60.18 1.135 ;
      RECT 60.17 0.905 60.175 1.138 ;
      RECT 60.16 0.91 60.17 1.142 ;
      RECT 60.155 0.917 60.16 1.147 ;
      RECT 60.145 0.922 60.155 1.151 ;
      RECT 60.12 0.934 60.145 1.162 ;
      RECT 60.1 0.951 60.12 1.178 ;
      RECT 60.075 0.968 60.1 1.2 ;
      RECT 60.04 0.991 60.075 1.258 ;
      RECT 60.02 1.013 60.04 1.32 ;
      RECT 60.015 1.023 60.02 1.355 ;
      RECT 60.005 1.03 60.015 1.393 ;
      RECT 60 1.037 60.005 1.413 ;
      RECT 59.995 1.048 60 1.45 ;
      RECT 59.99 1.056 59.995 1.515 ;
      RECT 59.98 1.067 59.99 1.568 ;
      RECT 59.975 1.085 59.98 1.638 ;
      RECT 59.97 1.095 59.975 1.675 ;
      RECT 59.965 1.105 59.97 1.97 ;
      RECT 59.96 1.117 59.965 1.97 ;
      RECT 59.955 1.127 59.96 1.97 ;
      RECT 59.945 1.137 59.955 1.97 ;
      RECT 59.935 1.16 59.945 1.97 ;
      RECT 59.92 1.195 59.935 1.97 ;
      RECT 59.88 1.257 59.92 1.97 ;
      RECT 59.875 1.31 59.88 1.97 ;
      RECT 59.85 1.345 59.875 1.97 ;
      RECT 59.835 1.39 59.85 1.97 ;
      RECT 59.83 1.412 59.835 1.97 ;
      RECT 59.82 1.425 59.83 1.97 ;
      RECT 59.81 1.45 59.82 1.97 ;
      RECT 59.805 1.472 59.81 1.97 ;
      RECT 59.78 1.51 59.8 1.97 ;
      RECT 59.74 1.567 59.78 1.97 ;
      RECT 59.735 1.617 59.74 1.97 ;
      RECT 59.73 1.635 59.735 1.97 ;
      RECT 59.725 1.647 59.73 1.97 ;
      RECT 59.715 1.665 59.725 1.97 ;
      RECT 59.705 1.685 59.715 1.945 ;
      RECT 59.7 1.702 59.705 1.945 ;
      RECT 59.69 1.715 59.7 1.945 ;
      RECT 59.66 1.725 59.685 1.945 ;
      RECT 59.65 1.732 59.66 1.945 ;
      RECT 59.635 1.742 59.65 1.94 ;
      RECT 58.595 1.655 58.915 1.915 ;
      RECT 58.46 1.7 58.915 1.87 ;
      RECT 51.96 1.515 52.335 1.765 ;
      RECT 52.06 0.73 52.235 1.765 ;
      RECT 57.74 0.715 58.06 0.975 ;
      RECT 57.74 0.745 58.14 0.915 ;
      RECT 52.06 0.73 58.06 0.905 ;
      RECT 55.405 1.755 55.7 2.045 ;
      RECT 55.375 1.755 55.7 2.015 ;
      RECT 41.615 2.125 41.92 2.355 ;
      RECT 49.755 2.155 53.17 2.33 ;
      RECT 52.995 1.305 53.17 2.33 ;
      RECT 41.615 2.155 53.17 2.325 ;
      RECT 52.94 1.305 53.27 1.555 ;
      RECT 50.2 1.315 50.49 1.555 ;
      RECT 45.75 1.285 46.01 1.52 ;
      RECT 45.75 1.315 50.49 1.485 ;
      RECT 48.935 1.655 49.255 1.915 ;
      RECT 48.92 1.7 49.255 1.87 ;
      RECT 47.64 0.635 47.935 0.925 ;
      RECT 47.605 0.635 47.935 0.895 ;
      RECT 44.8 1.655 45.12 1.915 ;
      RECT 44.785 1.7 45.12 1.87 ;
      RECT 43.125 1.445 43.445 1.705 ;
      RECT 43.11 1.445 43.465 1.68 ;
      RECT 40.425 1.205 40.61 1.415 ;
      RECT 40.415 1.21 40.625 1.408 ;
      RECT 40.415 1.21 40.711 1.385 ;
      RECT 40.415 1.21 40.77 1.36 ;
      RECT 40.415 1.21 40.825 1.34 ;
      RECT 40.415 1.21 40.835 1.328 ;
      RECT 40.415 1.21 41.03 1.267 ;
      RECT 40.415 1.21 41.06 1.25 ;
      RECT 40.415 1.21 41.08 1.24 ;
      RECT 40.96 0.975 41.22 1.235 ;
      RECT 40.945 1.065 40.96 1.282 ;
      RECT 40.48 1.197 41.22 1.235 ;
      RECT 40.931 1.076 40.945 1.288 ;
      RECT 40.52 1.19 41.22 1.235 ;
      RECT 40.845 1.116 40.931 1.307 ;
      RECT 40.77 1.177 41.22 1.235 ;
      RECT 40.84 1.152 40.845 1.324 ;
      RECT 40.825 1.162 41.22 1.235 ;
      RECT 40.835 1.157 40.84 1.326 ;
      RECT 41.13 1.662 41.135 1.754 ;
      RECT 41.125 1.64 41.13 1.771 ;
      RECT 41.12 1.63 41.125 1.783 ;
      RECT 41.11 1.621 41.12 1.793 ;
      RECT 41.105 1.616 41.11 1.801 ;
      RECT 41.1 1.612 41.105 1.804 ;
      RECT 41.066 1.545 41.1 1.815 ;
      RECT 40.98 1.545 41.066 1.85 ;
      RECT 40.9 1.545 40.98 1.898 ;
      RECT 40.84 1.545 40.9 1.923 ;
      RECT 40.78 1.645 40.84 1.93 ;
      RECT 40.745 1.67 40.78 1.936 ;
      RECT 40.72 1.685 40.745 1.94 ;
      RECT 40.706 1.694 40.72 1.942 ;
      RECT 40.62 1.721 40.706 1.948 ;
      RECT 40.555 1.762 40.62 1.957 ;
      RECT 40.54 1.782 40.555 1.962 ;
      RECT 40.51 1.792 40.54 1.965 ;
      RECT 40.505 1.802 40.51 1.968 ;
      RECT 40.475 1.807 40.505 1.97 ;
      RECT 40.455 1.812 40.475 1.974 ;
      RECT 40.37 1.815 40.455 1.981 ;
      RECT 40.355 1.812 40.37 1.987 ;
      RECT 40.345 1.809 40.355 1.989 ;
      RECT 40.325 1.806 40.345 1.991 ;
      RECT 40.305 1.802 40.325 1.992 ;
      RECT 40.29 1.798 40.305 1.994 ;
      RECT 40.28 1.795 40.29 1.995 ;
      RECT 40.24 1.789 40.28 1.993 ;
      RECT 40.23 1.784 40.24 1.991 ;
      RECT 40.215 1.781 40.23 1.987 ;
      RECT 40.19 1.776 40.215 1.98 ;
      RECT 40.14 1.767 40.19 1.968 ;
      RECT 40.07 1.753 40.14 1.95 ;
      RECT 40.012 1.738 40.07 1.932 ;
      RECT 39.926 1.721 40.012 1.912 ;
      RECT 39.84 1.7 39.926 1.887 ;
      RECT 39.79 1.685 39.84 1.868 ;
      RECT 39.786 1.679 39.79 1.86 ;
      RECT 39.7 1.669 39.786 1.847 ;
      RECT 39.665 1.654 39.7 1.83 ;
      RECT 39.65 1.647 39.665 1.823 ;
      RECT 39.59 1.635 39.65 1.811 ;
      RECT 39.57 1.622 39.59 1.799 ;
      RECT 39.53 1.613 39.57 1.791 ;
      RECT 39.525 1.605 39.53 1.784 ;
      RECT 39.445 1.595 39.525 1.77 ;
      RECT 39.43 1.582 39.445 1.755 ;
      RECT 39.425 1.58 39.43 1.753 ;
      RECT 39.346 1.568 39.425 1.74 ;
      RECT 39.26 1.543 39.346 1.715 ;
      RECT 39.245 1.512 39.26 1.7 ;
      RECT 39.23 1.487 39.245 1.696 ;
      RECT 39.215 1.48 39.23 1.692 ;
      RECT 39.04 1.485 39.045 1.688 ;
      RECT 39.035 1.49 39.04 1.683 ;
      RECT 39.045 1.48 39.215 1.69 ;
      RECT 39.76 1.24 39.865 1.5 ;
      RECT 40.575 0.765 40.58 0.99 ;
      RECT 40.705 0.765 40.76 0.975 ;
      RECT 40.76 0.77 40.77 0.968 ;
      RECT 40.666 0.765 40.705 0.978 ;
      RECT 40.58 0.765 40.666 0.985 ;
      RECT 40.56 0.77 40.575 0.991 ;
      RECT 40.55 0.81 40.56 0.993 ;
      RECT 40.52 0.82 40.55 0.995 ;
      RECT 40.515 0.825 40.52 0.997 ;
      RECT 40.49 0.83 40.515 0.999 ;
      RECT 40.475 0.835 40.49 1.001 ;
      RECT 40.46 0.837 40.475 1.003 ;
      RECT 40.455 0.842 40.46 1.005 ;
      RECT 40.405 0.85 40.455 1.008 ;
      RECT 40.38 0.859 40.405 1.013 ;
      RECT 40.37 0.866 40.38 1.018 ;
      RECT 40.365 0.869 40.37 1.022 ;
      RECT 40.345 0.872 40.365 1.031 ;
      RECT 40.315 0.88 40.345 1.051 ;
      RECT 40.286 0.893 40.315 1.073 ;
      RECT 40.2 0.927 40.286 1.117 ;
      RECT 40.195 0.953 40.2 1.155 ;
      RECT 40.19 0.957 40.195 1.164 ;
      RECT 40.155 0.97 40.19 1.197 ;
      RECT 40.145 0.984 40.155 1.235 ;
      RECT 40.14 0.988 40.145 1.248 ;
      RECT 40.135 0.992 40.14 1.253 ;
      RECT 40.125 1 40.135 1.265 ;
      RECT 40.12 1.007 40.125 1.28 ;
      RECT 40.095 1.02 40.12 1.305 ;
      RECT 40.055 1.049 40.095 1.36 ;
      RECT 40.04 1.074 40.055 1.415 ;
      RECT 40.03 1.085 40.04 1.438 ;
      RECT 40.025 1.092 40.03 1.45 ;
      RECT 40.02 1.096 40.025 1.458 ;
      RECT 39.965 1.124 40.02 1.5 ;
      RECT 39.945 1.16 39.965 1.5 ;
      RECT 39.93 1.175 39.945 1.5 ;
      RECT 39.875 1.207 39.93 1.5 ;
      RECT 39.865 1.237 39.875 1.5 ;
      RECT 39.475 0.852 39.66 1.09 ;
      RECT 39.46 0.854 39.67 1.085 ;
      RECT 39.345 0.8 39.605 1.06 ;
      RECT 39.34 0.837 39.605 1.014 ;
      RECT 39.335 0.847 39.605 1.011 ;
      RECT 39.33 0.887 39.67 1.005 ;
      RECT 39.325 0.92 39.67 0.995 ;
      RECT 39.335 0.862 39.685 0.933 ;
      RECT 39.632 1.96 39.645 2.49 ;
      RECT 39.546 1.96 39.645 2.489 ;
      RECT 39.546 1.96 39.65 2.488 ;
      RECT 39.46 1.96 39.65 2.486 ;
      RECT 39.455 1.96 39.65 2.483 ;
      RECT 39.455 1.96 39.66 2.481 ;
      RECT 39.45 2.252 39.66 2.478 ;
      RECT 39.45 2.262 39.665 2.475 ;
      RECT 39.45 2.33 39.67 2.471 ;
      RECT 39.44 2.335 39.67 2.47 ;
      RECT 39.44 2.427 39.675 2.467 ;
      RECT 39.425 1.96 39.685 2.22 ;
      RECT 38.655 0.95 38.7 2.485 ;
      RECT 38.855 0.95 38.885 1.165 ;
      RECT 37.23 0.69 37.35 0.9 ;
      RECT 36.89 0.64 37.15 0.9 ;
      RECT 36.89 0.685 37.185 0.89 ;
      RECT 38.895 0.966 38.9 1.02 ;
      RECT 38.89 0.959 38.895 1.153 ;
      RECT 38.885 0.953 38.89 1.16 ;
      RECT 38.84 0.95 38.855 1.173 ;
      RECT 38.835 0.95 38.84 1.195 ;
      RECT 38.83 0.95 38.835 1.243 ;
      RECT 38.825 0.95 38.83 1.263 ;
      RECT 38.815 0.95 38.825 1.37 ;
      RECT 38.81 0.95 38.815 1.433 ;
      RECT 38.805 0.95 38.81 1.49 ;
      RECT 38.8 0.95 38.805 1.498 ;
      RECT 38.785 0.95 38.8 1.605 ;
      RECT 38.775 0.95 38.785 1.74 ;
      RECT 38.765 0.95 38.775 1.85 ;
      RECT 38.755 0.95 38.765 1.907 ;
      RECT 38.75 0.95 38.755 1.947 ;
      RECT 38.745 0.95 38.75 1.983 ;
      RECT 38.735 0.95 38.745 2.023 ;
      RECT 38.73 0.95 38.735 2.065 ;
      RECT 38.71 0.95 38.73 2.13 ;
      RECT 38.715 2.275 38.72 2.455 ;
      RECT 38.71 2.257 38.715 2.463 ;
      RECT 38.705 0.95 38.71 2.193 ;
      RECT 38.705 2.237 38.71 2.47 ;
      RECT 38.7 0.95 38.705 2.48 ;
      RECT 38.645 0.95 38.655 1.25 ;
      RECT 38.65 1.497 38.655 2.485 ;
      RECT 38.645 1.562 38.65 2.485 ;
      RECT 38.64 0.951 38.645 1.24 ;
      RECT 38.635 1.627 38.645 2.485 ;
      RECT 38.63 0.952 38.64 1.23 ;
      RECT 38.62 1.74 38.635 2.485 ;
      RECT 38.625 0.953 38.63 1.22 ;
      RECT 38.605 0.954 38.625 1.198 ;
      RECT 38.61 1.837 38.62 2.485 ;
      RECT 38.605 1.912 38.61 2.485 ;
      RECT 38.595 0.953 38.605 1.175 ;
      RECT 38.6 1.955 38.605 2.485 ;
      RECT 38.595 1.982 38.6 2.485 ;
      RECT 38.585 0.951 38.595 1.163 ;
      RECT 38.59 2.025 38.595 2.485 ;
      RECT 38.585 2.052 38.59 2.485 ;
      RECT 38.575 0.95 38.585 1.15 ;
      RECT 38.58 2.067 38.585 2.485 ;
      RECT 38.54 2.125 38.58 2.485 ;
      RECT 38.57 0.949 38.575 1.135 ;
      RECT 38.565 0.947 38.57 1.128 ;
      RECT 38.555 0.944 38.565 1.118 ;
      RECT 38.55 0.941 38.555 1.103 ;
      RECT 38.535 0.937 38.55 1.096 ;
      RECT 38.53 2.18 38.54 2.485 ;
      RECT 38.53 0.934 38.535 1.091 ;
      RECT 38.515 0.93 38.53 1.085 ;
      RECT 38.525 2.197 38.53 2.485 ;
      RECT 38.515 2.26 38.525 2.485 ;
      RECT 38.435 0.915 38.515 1.065 ;
      RECT 38.51 2.267 38.515 2.48 ;
      RECT 38.505 2.275 38.51 2.47 ;
      RECT 38.425 0.901 38.435 1.049 ;
      RECT 38.41 0.897 38.425 1.047 ;
      RECT 38.4 0.892 38.41 1.043 ;
      RECT 38.375 0.885 38.4 1.035 ;
      RECT 38.37 0.88 38.375 1.03 ;
      RECT 38.36 0.88 38.37 1.028 ;
      RECT 38.35 0.878 38.36 1.026 ;
      RECT 38.32 0.87 38.35 1.02 ;
      RECT 38.305 0.862 38.32 1.013 ;
      RECT 38.285 0.857 38.305 1.006 ;
      RECT 38.28 0.853 38.285 1.001 ;
      RECT 38.25 0.846 38.28 0.995 ;
      RECT 38.225 0.837 38.25 0.985 ;
      RECT 38.195 0.83 38.225 0.977 ;
      RECT 38.17 0.82 38.195 0.968 ;
      RECT 38.155 0.812 38.17 0.962 ;
      RECT 38.13 0.807 38.155 0.957 ;
      RECT 38.12 0.803 38.13 0.952 ;
      RECT 38.1 0.798 38.12 0.947 ;
      RECT 38.065 0.793 38.1 0.94 ;
      RECT 38.005 0.788 38.065 0.933 ;
      RECT 37.992 0.784 38.005 0.931 ;
      RECT 37.906 0.779 37.992 0.928 ;
      RECT 37.82 0.769 37.906 0.924 ;
      RECT 37.779 0.762 37.82 0.921 ;
      RECT 37.693 0.755 37.779 0.918 ;
      RECT 37.607 0.745 37.693 0.914 ;
      RECT 37.521 0.735 37.607 0.909 ;
      RECT 37.435 0.725 37.521 0.905 ;
      RECT 37.425 0.71 37.435 0.903 ;
      RECT 37.415 0.695 37.425 0.903 ;
      RECT 37.35 0.69 37.415 0.902 ;
      RECT 37.185 0.687 37.23 0.895 ;
      RECT 38.43 1.592 38.435 1.783 ;
      RECT 38.425 1.587 38.43 1.79 ;
      RECT 38.411 1.585 38.425 1.796 ;
      RECT 38.325 1.585 38.411 1.798 ;
      RECT 38.321 1.585 38.325 1.801 ;
      RECT 38.235 1.585 38.321 1.819 ;
      RECT 38.225 1.59 38.235 1.838 ;
      RECT 38.215 1.645 38.225 1.842 ;
      RECT 38.19 1.66 38.215 1.849 ;
      RECT 38.15 1.68 38.19 1.862 ;
      RECT 38.145 1.692 38.15 1.872 ;
      RECT 38.13 1.698 38.145 1.877 ;
      RECT 38.125 1.703 38.13 1.881 ;
      RECT 38.105 1.71 38.125 1.886 ;
      RECT 38.035 1.735 38.105 1.903 ;
      RECT 37.995 1.763 38.035 1.923 ;
      RECT 37.99 1.773 37.995 1.931 ;
      RECT 37.97 1.78 37.99 1.933 ;
      RECT 37.965 1.787 37.97 1.936 ;
      RECT 37.935 1.795 37.965 1.939 ;
      RECT 37.93 1.8 37.935 1.943 ;
      RECT 37.856 1.804 37.93 1.951 ;
      RECT 37.77 1.813 37.856 1.967 ;
      RECT 37.766 1.818 37.77 1.976 ;
      RECT 37.68 1.823 37.766 1.986 ;
      RECT 37.64 1.831 37.68 1.998 ;
      RECT 37.59 1.837 37.64 2.005 ;
      RECT 37.505 1.846 37.59 2.02 ;
      RECT 37.43 1.857 37.505 2.038 ;
      RECT 37.395 1.864 37.43 2.048 ;
      RECT 37.32 1.872 37.395 2.053 ;
      RECT 37.265 1.881 37.32 2.053 ;
      RECT 37.24 1.886 37.265 2.051 ;
      RECT 37.23 1.889 37.24 2.049 ;
      RECT 37.195 1.891 37.23 2.047 ;
      RECT 37.165 1.893 37.195 2.043 ;
      RECT 37.12 1.892 37.165 2.039 ;
      RECT 37.1 1.887 37.12 2.036 ;
      RECT 37.05 1.872 37.1 2.033 ;
      RECT 37.04 1.857 37.05 2.028 ;
      RECT 36.99 1.842 37.04 2.018 ;
      RECT 36.94 1.817 36.99 1.998 ;
      RECT 36.93 1.802 36.94 1.98 ;
      RECT 36.925 1.8 36.93 1.974 ;
      RECT 36.905 1.795 36.925 1.969 ;
      RECT 36.9 1.787 36.905 1.963 ;
      RECT 36.885 1.781 36.9 1.956 ;
      RECT 36.88 1.776 36.885 1.948 ;
      RECT 36.86 1.771 36.88 1.94 ;
      RECT 36.845 1.764 36.86 1.933 ;
      RECT 36.83 1.758 36.845 1.924 ;
      RECT 36.825 1.752 36.83 1.917 ;
      RECT 36.78 1.727 36.825 1.903 ;
      RECT 36.765 1.697 36.78 1.885 ;
      RECT 36.75 1.68 36.765 1.876 ;
      RECT 36.725 1.66 36.75 1.864 ;
      RECT 36.685 1.63 36.725 1.844 ;
      RECT 36.675 1.6 36.685 1.829 ;
      RECT 36.66 1.59 36.675 1.822 ;
      RECT 36.605 1.555 36.66 1.801 ;
      RECT 36.59 1.518 36.605 1.78 ;
      RECT 36.58 1.505 36.59 1.772 ;
      RECT 36.53 1.475 36.58 1.754 ;
      RECT 36.515 1.405 36.53 1.735 ;
      RECT 36.47 1.405 36.515 1.718 ;
      RECT 36.445 1.405 36.47 1.7 ;
      RECT 36.435 1.405 36.445 1.693 ;
      RECT 36.356 1.405 36.435 1.686 ;
      RECT 36.27 1.405 36.356 1.678 ;
      RECT 36.255 1.437 36.27 1.673 ;
      RECT 36.18 1.447 36.255 1.669 ;
      RECT 36.16 1.457 36.18 1.664 ;
      RECT 36.135 1.457 36.16 1.661 ;
      RECT 36.125 1.447 36.135 1.66 ;
      RECT 36.115 1.42 36.125 1.659 ;
      RECT 36.075 1.415 36.115 1.657 ;
      RECT 36.03 1.415 36.075 1.653 ;
      RECT 36.005 1.415 36.03 1.648 ;
      RECT 35.955 1.415 36.005 1.635 ;
      RECT 35.915 1.42 35.925 1.62 ;
      RECT 35.925 1.415 35.955 1.625 ;
      RECT 37.91 1.195 38.17 1.455 ;
      RECT 37.905 1.217 38.17 1.413 ;
      RECT 37.145 1.045 37.365 1.41 ;
      RECT 37.127 1.132 37.365 1.409 ;
      RECT 37.11 1.137 37.365 1.406 ;
      RECT 37.11 1.137 37.385 1.405 ;
      RECT 37.08 1.147 37.385 1.403 ;
      RECT 37.075 1.162 37.385 1.399 ;
      RECT 37.075 1.162 37.39 1.398 ;
      RECT 37.07 1.22 37.39 1.396 ;
      RECT 37.07 1.22 37.4 1.393 ;
      RECT 37.065 1.285 37.4 1.388 ;
      RECT 37.145 1.045 37.405 1.305 ;
      RECT 35.89 0.875 36.15 1.135 ;
      RECT 35.89 0.918 36.236 1.109 ;
      RECT 35.89 0.918 36.28 1.108 ;
      RECT 35.89 0.918 36.3 1.106 ;
      RECT 35.89 0.918 36.4 1.105 ;
      RECT 35.89 0.918 36.42 1.103 ;
      RECT 35.89 0.918 36.43 1.098 ;
      RECT 36.3 0.885 36.49 1.095 ;
      RECT 36.3 0.887 36.495 1.093 ;
      RECT 36.29 0.892 36.5 1.085 ;
      RECT 36.236 0.916 36.5 1.085 ;
      RECT 36.28 0.91 36.29 1.107 ;
      RECT 36.29 0.89 36.495 1.093 ;
      RECT 35.245 1.95 35.45 2.18 ;
      RECT 35.185 1.9 35.24 2.16 ;
      RECT 35.245 1.9 35.445 2.18 ;
      RECT 36.215 2.215 36.22 2.242 ;
      RECT 36.205 2.125 36.215 2.247 ;
      RECT 36.2 2.047 36.205 2.253 ;
      RECT 36.19 2.037 36.2 2.26 ;
      RECT 36.185 2.027 36.19 2.266 ;
      RECT 36.175 2.022 36.185 2.268 ;
      RECT 36.16 2.014 36.175 2.276 ;
      RECT 36.145 2.005 36.16 2.288 ;
      RECT 36.135 1.997 36.145 2.298 ;
      RECT 36.1 1.915 36.135 2.316 ;
      RECT 36.065 1.915 36.1 2.335 ;
      RECT 36.05 1.915 36.065 2.343 ;
      RECT 35.995 1.915 36.05 2.343 ;
      RECT 35.961 1.915 35.995 2.334 ;
      RECT 35.875 1.915 35.961 2.31 ;
      RECT 35.865 1.975 35.875 2.292 ;
      RECT 35.825 1.977 35.865 2.283 ;
      RECT 35.82 1.979 35.825 2.273 ;
      RECT 35.8 1.981 35.82 2.268 ;
      RECT 35.79 1.984 35.8 2.263 ;
      RECT 35.78 1.985 35.79 2.258 ;
      RECT 35.756 1.986 35.78 2.25 ;
      RECT 35.67 1.991 35.756 2.228 ;
      RECT 35.615 1.99 35.67 2.201 ;
      RECT 35.6 1.983 35.615 2.188 ;
      RECT 35.565 1.978 35.6 2.184 ;
      RECT 35.51 1.97 35.565 2.183 ;
      RECT 35.45 1.957 35.51 2.181 ;
      RECT 35.24 1.9 35.245 2.168 ;
      RECT 35.315 1.27 35.5 1.48 ;
      RECT 35.305 1.275 35.515 1.473 ;
      RECT 35.345 1.18 35.605 1.44 ;
      RECT 35.3 1.337 35.605 1.363 ;
      RECT 34.645 1.13 34.65 1.93 ;
      RECT 34.59 1.18 34.62 1.93 ;
      RECT 34.58 1.18 34.585 1.49 ;
      RECT 34.565 1.18 34.57 1.485 ;
      RECT 34.11 1.225 34.125 1.44 ;
      RECT 34.04 1.225 34.125 1.435 ;
      RECT 35.305 0.805 35.375 1.015 ;
      RECT 35.375 0.812 35.385 1.01 ;
      RECT 35.271 0.805 35.305 1.022 ;
      RECT 35.185 0.805 35.271 1.046 ;
      RECT 35.175 0.81 35.185 1.065 ;
      RECT 35.17 0.822 35.175 1.068 ;
      RECT 35.155 0.837 35.17 1.072 ;
      RECT 35.15 0.855 35.155 1.076 ;
      RECT 35.11 0.865 35.15 1.085 ;
      RECT 35.095 0.872 35.11 1.097 ;
      RECT 35.08 0.877 35.095 1.102 ;
      RECT 35.065 0.88 35.08 1.107 ;
      RECT 35.055 0.882 35.065 1.111 ;
      RECT 35.02 0.889 35.055 1.119 ;
      RECT 34.985 0.897 35.02 1.133 ;
      RECT 34.975 0.903 34.985 1.142 ;
      RECT 34.97 0.905 34.975 1.144 ;
      RECT 34.95 0.908 34.97 1.15 ;
      RECT 34.92 0.915 34.95 1.161 ;
      RECT 34.91 0.921 34.92 1.168 ;
      RECT 34.885 0.924 34.91 1.175 ;
      RECT 34.875 0.928 34.885 1.183 ;
      RECT 34.87 0.929 34.875 1.205 ;
      RECT 34.865 0.93 34.87 1.22 ;
      RECT 34.86 0.931 34.865 1.235 ;
      RECT 34.855 0.932 34.86 1.25 ;
      RECT 34.85 0.933 34.855 1.28 ;
      RECT 34.84 0.935 34.85 1.313 ;
      RECT 34.825 0.939 34.84 1.36 ;
      RECT 34.815 0.942 34.825 1.405 ;
      RECT 34.81 0.945 34.815 1.433 ;
      RECT 34.8 0.947 34.81 1.46 ;
      RECT 34.795 0.95 34.8 1.495 ;
      RECT 34.765 0.955 34.795 1.553 ;
      RECT 34.76 0.96 34.765 1.638 ;
      RECT 34.755 0.962 34.76 1.673 ;
      RECT 34.75 0.964 34.755 1.755 ;
      RECT 34.745 0.966 34.75 1.843 ;
      RECT 34.735 0.968 34.745 1.925 ;
      RECT 34.72 0.982 34.735 1.93 ;
      RECT 34.685 1.027 34.72 1.93 ;
      RECT 34.675 1.067 34.685 1.93 ;
      RECT 34.66 1.095 34.675 1.93 ;
      RECT 34.655 1.112 34.66 1.93 ;
      RECT 34.65 1.12 34.655 1.93 ;
      RECT 34.64 1.135 34.645 1.93 ;
      RECT 34.635 1.142 34.64 1.93 ;
      RECT 34.625 1.162 34.635 1.93 ;
      RECT 34.62 1.175 34.625 1.93 ;
      RECT 34.585 1.18 34.59 1.515 ;
      RECT 34.57 1.57 34.59 1.93 ;
      RECT 34.57 1.18 34.58 1.488 ;
      RECT 34.565 1.61 34.57 1.93 ;
      RECT 34.515 1.18 34.565 1.483 ;
      RECT 34.56 1.647 34.565 1.93 ;
      RECT 34.55 1.67 34.56 1.93 ;
      RECT 34.545 1.715 34.55 1.93 ;
      RECT 34.535 1.725 34.545 1.923 ;
      RECT 34.461 1.18 34.515 1.477 ;
      RECT 34.375 1.18 34.461 1.47 ;
      RECT 34.326 1.227 34.375 1.463 ;
      RECT 34.24 1.235 34.326 1.456 ;
      RECT 34.225 1.232 34.24 1.451 ;
      RECT 34.211 1.225 34.225 1.45 ;
      RECT 34.125 1.225 34.211 1.445 ;
      RECT 34.03 1.23 34.04 1.43 ;
      RECT 33.62 0.66 33.635 1.06 ;
      RECT 33.815 0.66 33.82 0.92 ;
      RECT 33.56 0.66 33.605 0.92 ;
      RECT 34.015 1.965 34.02 2.17 ;
      RECT 34.01 1.955 34.015 2.175 ;
      RECT 34.005 1.942 34.01 2.18 ;
      RECT 34 1.922 34.005 2.18 ;
      RECT 33.975 1.875 34 2.18 ;
      RECT 33.94 1.79 33.975 2.18 ;
      RECT 33.935 1.727 33.94 2.18 ;
      RECT 33.93 1.712 33.935 2.18 ;
      RECT 33.915 1.672 33.93 2.18 ;
      RECT 33.91 1.647 33.915 2.18 ;
      RECT 33.9 1.63 33.91 2.18 ;
      RECT 33.865 1.552 33.9 2.18 ;
      RECT 33.86 1.495 33.865 2.18 ;
      RECT 33.855 1.482 33.86 2.18 ;
      RECT 33.845 1.46 33.855 2.18 ;
      RECT 33.835 1.425 33.845 2.18 ;
      RECT 33.825 1.395 33.835 2.18 ;
      RECT 33.815 1.31 33.825 1.823 ;
      RECT 33.822 1.955 33.825 2.18 ;
      RECT 33.82 1.965 33.822 2.18 ;
      RECT 33.81 1.975 33.82 2.175 ;
      RECT 33.805 0.66 33.815 1.055 ;
      RECT 33.81 1.187 33.815 1.798 ;
      RECT 33.805 1.085 33.81 1.781 ;
      RECT 33.795 0.66 33.805 1.757 ;
      RECT 33.79 0.66 33.795 1.728 ;
      RECT 33.785 0.66 33.79 1.718 ;
      RECT 33.765 0.66 33.785 1.68 ;
      RECT 33.76 0.66 33.765 1.638 ;
      RECT 33.755 0.66 33.76 1.618 ;
      RECT 33.725 0.66 33.755 1.568 ;
      RECT 33.715 0.66 33.725 1.515 ;
      RECT 33.71 0.66 33.715 1.488 ;
      RECT 33.705 0.66 33.71 1.473 ;
      RECT 33.695 0.66 33.705 1.45 ;
      RECT 33.685 0.66 33.695 1.425 ;
      RECT 33.68 0.66 33.685 1.365 ;
      RECT 33.67 0.66 33.68 1.303 ;
      RECT 33.665 0.66 33.67 1.223 ;
      RECT 33.66 0.66 33.665 1.188 ;
      RECT 33.655 0.66 33.66 1.163 ;
      RECT 33.65 0.66 33.655 1.148 ;
      RECT 33.645 0.66 33.65 1.118 ;
      RECT 33.64 0.66 33.645 1.095 ;
      RECT 33.635 0.66 33.64 1.068 ;
      RECT 33.605 0.66 33.62 1.055 ;
      RECT 32.76 2.195 32.945 2.405 ;
      RECT 32.75 2.2 32.96 2.398 ;
      RECT 32.75 2.2 32.98 2.37 ;
      RECT 32.75 2.2 32.995 2.349 ;
      RECT 32.75 2.2 33.01 2.347 ;
      RECT 32.75 2.2 33.02 2.346 ;
      RECT 32.75 2.2 33.05 2.343 ;
      RECT 33.4 2.045 33.66 2.305 ;
      RECT 33.36 2.092 33.66 2.288 ;
      RECT 33.351 2.1 33.36 2.291 ;
      RECT 32.945 2.193 33.66 2.288 ;
      RECT 33.265 2.118 33.351 2.298 ;
      RECT 32.96 2.19 33.66 2.288 ;
      RECT 33.206 2.14 33.265 2.31 ;
      RECT 32.98 2.186 33.66 2.288 ;
      RECT 33.12 2.152 33.206 2.321 ;
      RECT 32.995 2.182 33.66 2.288 ;
      RECT 33.065 2.165 33.12 2.333 ;
      RECT 33.01 2.18 33.66 2.288 ;
      RECT 33.05 2.171 33.065 2.339 ;
      RECT 33.02 2.176 33.66 2.288 ;
      RECT 33.165 1.7 33.425 1.96 ;
      RECT 33.165 1.72 33.535 1.93 ;
      RECT 33.165 1.725 33.545 1.925 ;
      RECT 33.356 1.139 33.435 1.37 ;
      RECT 33.27 1.142 33.485 1.365 ;
      RECT 33.265 1.142 33.485 1.36 ;
      RECT 33.265 1.147 33.495 1.358 ;
      RECT 33.24 1.147 33.495 1.355 ;
      RECT 33.24 1.155 33.505 1.353 ;
      RECT 33.12 1.09 33.38 1.35 ;
      RECT 33.12 1.137 33.43 1.35 ;
      RECT 32.375 1.71 32.38 1.97 ;
      RECT 32.205 1.48 32.21 1.97 ;
      RECT 32.09 1.72 32.095 1.945 ;
      RECT 32.8 0.815 32.805 1.025 ;
      RECT 32.805 0.82 32.82 1.02 ;
      RECT 32.74 0.815 32.8 1.033 ;
      RECT 32.725 0.815 32.74 1.043 ;
      RECT 32.675 0.815 32.725 1.06 ;
      RECT 32.655 0.815 32.675 1.083 ;
      RECT 32.64 0.815 32.655 1.095 ;
      RECT 32.62 0.815 32.64 1.105 ;
      RECT 32.61 0.82 32.62 1.114 ;
      RECT 32.605 0.83 32.61 1.119 ;
      RECT 32.6 0.842 32.605 1.123 ;
      RECT 32.59 0.865 32.6 1.128 ;
      RECT 32.585 0.88 32.59 1.132 ;
      RECT 32.58 0.897 32.585 1.135 ;
      RECT 32.575 0.905 32.58 1.138 ;
      RECT 32.565 0.91 32.575 1.142 ;
      RECT 32.56 0.917 32.565 1.147 ;
      RECT 32.55 0.922 32.56 1.151 ;
      RECT 32.525 0.934 32.55 1.162 ;
      RECT 32.505 0.951 32.525 1.178 ;
      RECT 32.48 0.968 32.505 1.2 ;
      RECT 32.445 0.991 32.48 1.258 ;
      RECT 32.425 1.013 32.445 1.32 ;
      RECT 32.42 1.023 32.425 1.355 ;
      RECT 32.41 1.03 32.42 1.393 ;
      RECT 32.405 1.037 32.41 1.413 ;
      RECT 32.4 1.048 32.405 1.45 ;
      RECT 32.395 1.056 32.4 1.515 ;
      RECT 32.385 1.067 32.395 1.568 ;
      RECT 32.38 1.085 32.385 1.638 ;
      RECT 32.375 1.095 32.38 1.675 ;
      RECT 32.37 1.105 32.375 1.97 ;
      RECT 32.365 1.117 32.37 1.97 ;
      RECT 32.36 1.127 32.365 1.97 ;
      RECT 32.35 1.137 32.36 1.97 ;
      RECT 32.34 1.16 32.35 1.97 ;
      RECT 32.325 1.195 32.34 1.97 ;
      RECT 32.285 1.257 32.325 1.97 ;
      RECT 32.28 1.31 32.285 1.97 ;
      RECT 32.255 1.345 32.28 1.97 ;
      RECT 32.24 1.39 32.255 1.97 ;
      RECT 32.235 1.412 32.24 1.97 ;
      RECT 32.225 1.425 32.235 1.97 ;
      RECT 32.215 1.45 32.225 1.97 ;
      RECT 32.21 1.472 32.215 1.97 ;
      RECT 32.185 1.51 32.205 1.97 ;
      RECT 32.145 1.567 32.185 1.97 ;
      RECT 32.14 1.617 32.145 1.97 ;
      RECT 32.135 1.635 32.14 1.97 ;
      RECT 32.13 1.647 32.135 1.97 ;
      RECT 32.12 1.665 32.13 1.97 ;
      RECT 32.11 1.685 32.12 1.945 ;
      RECT 32.105 1.702 32.11 1.945 ;
      RECT 32.095 1.715 32.105 1.945 ;
      RECT 32.065 1.725 32.09 1.945 ;
      RECT 32.055 1.732 32.065 1.945 ;
      RECT 32.04 1.742 32.055 1.94 ;
      RECT 31 1.655 31.32 1.915 ;
      RECT 30.865 1.7 31.32 1.87 ;
      RECT 24.37 1.475 24.745 1.725 ;
      RECT 24.465 0.73 24.64 1.725 ;
      RECT 30.145 0.715 30.465 0.975 ;
      RECT 30.145 0.745 30.545 0.915 ;
      RECT 24.465 0.73 30.465 0.905 ;
      RECT 27.81 1.755 28.105 2.045 ;
      RECT 27.78 1.755 28.105 2.015 ;
      RECT 14.02 2.125 14.325 2.355 ;
      RECT 22.16 2.155 25.575 2.33 ;
      RECT 25.4 1.305 25.575 2.33 ;
      RECT 14.02 2.155 25.575 2.325 ;
      RECT 25.345 1.305 25.675 1.555 ;
      RECT 22.605 1.315 22.895 1.555 ;
      RECT 18.155 1.285 18.415 1.52 ;
      RECT 18.155 1.315 22.895 1.485 ;
      RECT 21.34 1.655 21.66 1.915 ;
      RECT 21.325 1.7 21.66 1.87 ;
      RECT 20.045 0.635 20.34 0.925 ;
      RECT 20.01 0.635 20.34 0.895 ;
      RECT 17.205 1.655 17.525 1.915 ;
      RECT 17.19 1.7 17.525 1.87 ;
      RECT 15.53 1.445 15.85 1.705 ;
      RECT 15.515 1.445 15.87 1.68 ;
      RECT 12.83 1.205 13.015 1.415 ;
      RECT 12.82 1.21 13.03 1.408 ;
      RECT 12.82 1.21 13.116 1.385 ;
      RECT 12.82 1.21 13.175 1.36 ;
      RECT 12.82 1.21 13.23 1.34 ;
      RECT 12.82 1.21 13.24 1.328 ;
      RECT 12.82 1.21 13.435 1.267 ;
      RECT 12.82 1.21 13.465 1.25 ;
      RECT 12.82 1.21 13.485 1.24 ;
      RECT 13.365 0.975 13.625 1.235 ;
      RECT 13.35 1.065 13.365 1.282 ;
      RECT 12.885 1.197 13.625 1.235 ;
      RECT 13.336 1.076 13.35 1.288 ;
      RECT 12.925 1.19 13.625 1.235 ;
      RECT 13.25 1.116 13.336 1.307 ;
      RECT 13.175 1.177 13.625 1.235 ;
      RECT 13.245 1.152 13.25 1.324 ;
      RECT 13.23 1.162 13.625 1.235 ;
      RECT 13.24 1.157 13.245 1.326 ;
      RECT 13.535 1.662 13.54 1.754 ;
      RECT 13.53 1.64 13.535 1.771 ;
      RECT 13.525 1.63 13.53 1.783 ;
      RECT 13.515 1.621 13.525 1.793 ;
      RECT 13.51 1.616 13.515 1.801 ;
      RECT 13.505 1.612 13.51 1.804 ;
      RECT 13.471 1.545 13.505 1.815 ;
      RECT 13.385 1.545 13.471 1.85 ;
      RECT 13.305 1.545 13.385 1.898 ;
      RECT 13.245 1.545 13.305 1.923 ;
      RECT 13.185 1.645 13.245 1.93 ;
      RECT 13.15 1.67 13.185 1.936 ;
      RECT 13.125 1.685 13.15 1.94 ;
      RECT 13.111 1.694 13.125 1.942 ;
      RECT 13.025 1.721 13.111 1.948 ;
      RECT 12.96 1.762 13.025 1.957 ;
      RECT 12.945 1.782 12.96 1.962 ;
      RECT 12.915 1.792 12.945 1.965 ;
      RECT 12.91 1.802 12.915 1.968 ;
      RECT 12.88 1.807 12.91 1.97 ;
      RECT 12.86 1.812 12.88 1.974 ;
      RECT 12.775 1.815 12.86 1.981 ;
      RECT 12.76 1.812 12.775 1.987 ;
      RECT 12.75 1.809 12.76 1.989 ;
      RECT 12.73 1.806 12.75 1.991 ;
      RECT 12.71 1.802 12.73 1.992 ;
      RECT 12.695 1.798 12.71 1.994 ;
      RECT 12.685 1.795 12.695 1.995 ;
      RECT 12.645 1.789 12.685 1.993 ;
      RECT 12.635 1.784 12.645 1.991 ;
      RECT 12.62 1.781 12.635 1.987 ;
      RECT 12.595 1.776 12.62 1.98 ;
      RECT 12.545 1.767 12.595 1.968 ;
      RECT 12.475 1.753 12.545 1.95 ;
      RECT 12.417 1.738 12.475 1.932 ;
      RECT 12.331 1.721 12.417 1.912 ;
      RECT 12.245 1.7 12.331 1.887 ;
      RECT 12.195 1.685 12.245 1.868 ;
      RECT 12.191 1.679 12.195 1.86 ;
      RECT 12.105 1.669 12.191 1.847 ;
      RECT 12.07 1.654 12.105 1.83 ;
      RECT 12.055 1.647 12.07 1.823 ;
      RECT 11.995 1.635 12.055 1.811 ;
      RECT 11.975 1.622 11.995 1.799 ;
      RECT 11.935 1.613 11.975 1.791 ;
      RECT 11.93 1.605 11.935 1.784 ;
      RECT 11.85 1.595 11.93 1.77 ;
      RECT 11.835 1.582 11.85 1.755 ;
      RECT 11.83 1.58 11.835 1.753 ;
      RECT 11.751 1.568 11.83 1.74 ;
      RECT 11.665 1.543 11.751 1.715 ;
      RECT 11.65 1.512 11.665 1.7 ;
      RECT 11.635 1.487 11.65 1.696 ;
      RECT 11.62 1.48 11.635 1.692 ;
      RECT 11.445 1.485 11.45 1.688 ;
      RECT 11.44 1.49 11.445 1.683 ;
      RECT 11.45 1.48 11.62 1.69 ;
      RECT 12.165 1.24 12.27 1.5 ;
      RECT 12.98 0.765 12.985 0.99 ;
      RECT 13.11 0.765 13.165 0.975 ;
      RECT 13.165 0.77 13.175 0.968 ;
      RECT 13.071 0.765 13.11 0.978 ;
      RECT 12.985 0.765 13.071 0.985 ;
      RECT 12.965 0.77 12.98 0.991 ;
      RECT 12.955 0.81 12.965 0.993 ;
      RECT 12.925 0.82 12.955 0.995 ;
      RECT 12.92 0.825 12.925 0.997 ;
      RECT 12.895 0.83 12.92 0.999 ;
      RECT 12.88 0.835 12.895 1.001 ;
      RECT 12.865 0.837 12.88 1.003 ;
      RECT 12.86 0.842 12.865 1.005 ;
      RECT 12.81 0.85 12.86 1.008 ;
      RECT 12.785 0.859 12.81 1.013 ;
      RECT 12.775 0.866 12.785 1.018 ;
      RECT 12.77 0.869 12.775 1.022 ;
      RECT 12.75 0.872 12.77 1.031 ;
      RECT 12.72 0.88 12.75 1.051 ;
      RECT 12.691 0.893 12.72 1.073 ;
      RECT 12.605 0.927 12.691 1.117 ;
      RECT 12.6 0.953 12.605 1.155 ;
      RECT 12.595 0.957 12.6 1.164 ;
      RECT 12.56 0.97 12.595 1.197 ;
      RECT 12.55 0.984 12.56 1.235 ;
      RECT 12.545 0.988 12.55 1.248 ;
      RECT 12.54 0.992 12.545 1.253 ;
      RECT 12.53 1 12.54 1.265 ;
      RECT 12.525 1.007 12.53 1.28 ;
      RECT 12.5 1.02 12.525 1.305 ;
      RECT 12.46 1.049 12.5 1.36 ;
      RECT 12.445 1.074 12.46 1.415 ;
      RECT 12.435 1.085 12.445 1.438 ;
      RECT 12.43 1.092 12.435 1.45 ;
      RECT 12.425 1.096 12.43 1.458 ;
      RECT 12.37 1.124 12.425 1.5 ;
      RECT 12.35 1.16 12.37 1.5 ;
      RECT 12.335 1.175 12.35 1.5 ;
      RECT 12.28 1.207 12.335 1.5 ;
      RECT 12.27 1.237 12.28 1.5 ;
      RECT 11.88 0.852 12.065 1.09 ;
      RECT 11.865 0.854 12.075 1.085 ;
      RECT 11.75 0.8 12.01 1.06 ;
      RECT 11.745 0.837 12.01 1.014 ;
      RECT 11.74 0.847 12.01 1.011 ;
      RECT 11.735 0.887 12.075 1.005 ;
      RECT 11.73 0.92 12.075 0.995 ;
      RECT 11.74 0.862 12.09 0.933 ;
      RECT 12.037 1.96 12.05 2.49 ;
      RECT 11.951 1.96 12.05 2.489 ;
      RECT 11.951 1.96 12.055 2.488 ;
      RECT 11.865 1.96 12.055 2.486 ;
      RECT 11.86 1.96 12.055 2.483 ;
      RECT 11.86 1.96 12.065 2.481 ;
      RECT 11.855 2.252 12.065 2.478 ;
      RECT 11.855 2.262 12.07 2.475 ;
      RECT 11.855 2.33 12.075 2.471 ;
      RECT 11.845 2.335 12.075 2.47 ;
      RECT 11.845 2.427 12.08 2.467 ;
      RECT 11.83 1.96 12.09 2.22 ;
      RECT 11.06 0.95 11.105 2.485 ;
      RECT 11.26 0.95 11.29 1.165 ;
      RECT 9.635 0.69 9.755 0.9 ;
      RECT 9.295 0.64 9.555 0.9 ;
      RECT 9.295 0.685 9.59 0.89 ;
      RECT 11.3 0.966 11.305 1.02 ;
      RECT 11.295 0.959 11.3 1.153 ;
      RECT 11.29 0.953 11.295 1.16 ;
      RECT 11.245 0.95 11.26 1.173 ;
      RECT 11.24 0.95 11.245 1.195 ;
      RECT 11.235 0.95 11.24 1.243 ;
      RECT 11.23 0.95 11.235 1.263 ;
      RECT 11.22 0.95 11.23 1.37 ;
      RECT 11.215 0.95 11.22 1.433 ;
      RECT 11.21 0.95 11.215 1.49 ;
      RECT 11.205 0.95 11.21 1.498 ;
      RECT 11.19 0.95 11.205 1.605 ;
      RECT 11.18 0.95 11.19 1.74 ;
      RECT 11.17 0.95 11.18 1.85 ;
      RECT 11.16 0.95 11.17 1.907 ;
      RECT 11.155 0.95 11.16 1.947 ;
      RECT 11.15 0.95 11.155 1.983 ;
      RECT 11.14 0.95 11.15 2.023 ;
      RECT 11.135 0.95 11.14 2.065 ;
      RECT 11.115 0.95 11.135 2.13 ;
      RECT 11.12 2.275 11.125 2.455 ;
      RECT 11.115 2.257 11.12 2.463 ;
      RECT 11.11 0.95 11.115 2.193 ;
      RECT 11.11 2.237 11.115 2.47 ;
      RECT 11.105 0.95 11.11 2.48 ;
      RECT 11.05 0.95 11.06 1.25 ;
      RECT 11.055 1.497 11.06 2.485 ;
      RECT 11.05 1.562 11.055 2.485 ;
      RECT 11.045 0.951 11.05 1.24 ;
      RECT 11.04 1.627 11.05 2.485 ;
      RECT 11.035 0.952 11.045 1.23 ;
      RECT 11.025 1.74 11.04 2.485 ;
      RECT 11.03 0.953 11.035 1.22 ;
      RECT 11.01 0.954 11.03 1.198 ;
      RECT 11.015 1.837 11.025 2.485 ;
      RECT 11.01 1.912 11.015 2.485 ;
      RECT 11 0.953 11.01 1.175 ;
      RECT 11.005 1.955 11.01 2.485 ;
      RECT 11 1.982 11.005 2.485 ;
      RECT 10.99 0.951 11 1.163 ;
      RECT 10.995 2.025 11 2.485 ;
      RECT 10.99 2.052 10.995 2.485 ;
      RECT 10.98 0.95 10.99 1.15 ;
      RECT 10.985 2.067 10.99 2.485 ;
      RECT 10.945 2.125 10.985 2.485 ;
      RECT 10.975 0.949 10.98 1.135 ;
      RECT 10.97 0.947 10.975 1.128 ;
      RECT 10.96 0.944 10.97 1.118 ;
      RECT 10.955 0.941 10.96 1.103 ;
      RECT 10.94 0.937 10.955 1.096 ;
      RECT 10.935 2.18 10.945 2.485 ;
      RECT 10.935 0.934 10.94 1.091 ;
      RECT 10.92 0.93 10.935 1.085 ;
      RECT 10.93 2.197 10.935 2.485 ;
      RECT 10.92 2.26 10.93 2.485 ;
      RECT 10.84 0.915 10.92 1.065 ;
      RECT 10.915 2.267 10.92 2.48 ;
      RECT 10.91 2.275 10.915 2.47 ;
      RECT 10.83 0.901 10.84 1.049 ;
      RECT 10.815 0.897 10.83 1.047 ;
      RECT 10.805 0.892 10.815 1.043 ;
      RECT 10.78 0.885 10.805 1.035 ;
      RECT 10.775 0.88 10.78 1.03 ;
      RECT 10.765 0.88 10.775 1.028 ;
      RECT 10.755 0.878 10.765 1.026 ;
      RECT 10.725 0.87 10.755 1.02 ;
      RECT 10.71 0.862 10.725 1.013 ;
      RECT 10.69 0.857 10.71 1.006 ;
      RECT 10.685 0.853 10.69 1.001 ;
      RECT 10.655 0.846 10.685 0.995 ;
      RECT 10.63 0.837 10.655 0.985 ;
      RECT 10.6 0.83 10.63 0.977 ;
      RECT 10.575 0.82 10.6 0.968 ;
      RECT 10.56 0.812 10.575 0.962 ;
      RECT 10.535 0.807 10.56 0.957 ;
      RECT 10.525 0.803 10.535 0.952 ;
      RECT 10.505 0.798 10.525 0.947 ;
      RECT 10.47 0.793 10.505 0.94 ;
      RECT 10.41 0.788 10.47 0.933 ;
      RECT 10.397 0.784 10.41 0.931 ;
      RECT 10.311 0.779 10.397 0.928 ;
      RECT 10.225 0.769 10.311 0.924 ;
      RECT 10.184 0.762 10.225 0.921 ;
      RECT 10.098 0.755 10.184 0.918 ;
      RECT 10.012 0.745 10.098 0.914 ;
      RECT 9.926 0.735 10.012 0.909 ;
      RECT 9.84 0.725 9.926 0.905 ;
      RECT 9.83 0.71 9.84 0.903 ;
      RECT 9.82 0.695 9.83 0.903 ;
      RECT 9.755 0.69 9.82 0.902 ;
      RECT 9.59 0.687 9.635 0.895 ;
      RECT 10.835 1.592 10.84 1.783 ;
      RECT 10.83 1.587 10.835 1.79 ;
      RECT 10.816 1.585 10.83 1.796 ;
      RECT 10.73 1.585 10.816 1.798 ;
      RECT 10.726 1.585 10.73 1.801 ;
      RECT 10.64 1.585 10.726 1.819 ;
      RECT 10.63 1.59 10.64 1.838 ;
      RECT 10.62 1.645 10.63 1.842 ;
      RECT 10.595 1.66 10.62 1.849 ;
      RECT 10.555 1.68 10.595 1.862 ;
      RECT 10.55 1.692 10.555 1.872 ;
      RECT 10.535 1.698 10.55 1.877 ;
      RECT 10.53 1.703 10.535 1.881 ;
      RECT 10.51 1.71 10.53 1.886 ;
      RECT 10.44 1.735 10.51 1.903 ;
      RECT 10.4 1.763 10.44 1.923 ;
      RECT 10.395 1.773 10.4 1.931 ;
      RECT 10.375 1.78 10.395 1.933 ;
      RECT 10.37 1.787 10.375 1.936 ;
      RECT 10.34 1.795 10.37 1.939 ;
      RECT 10.335 1.8 10.34 1.943 ;
      RECT 10.261 1.804 10.335 1.951 ;
      RECT 10.175 1.813 10.261 1.967 ;
      RECT 10.171 1.818 10.175 1.976 ;
      RECT 10.085 1.823 10.171 1.986 ;
      RECT 10.045 1.831 10.085 1.998 ;
      RECT 9.995 1.837 10.045 2.005 ;
      RECT 9.91 1.846 9.995 2.02 ;
      RECT 9.835 1.857 9.91 2.038 ;
      RECT 9.8 1.864 9.835 2.048 ;
      RECT 9.725 1.872 9.8 2.053 ;
      RECT 9.67 1.881 9.725 2.053 ;
      RECT 9.645 1.886 9.67 2.051 ;
      RECT 9.635 1.889 9.645 2.049 ;
      RECT 9.6 1.891 9.635 2.047 ;
      RECT 9.57 1.893 9.6 2.043 ;
      RECT 9.525 1.892 9.57 2.039 ;
      RECT 9.505 1.887 9.525 2.036 ;
      RECT 9.455 1.872 9.505 2.033 ;
      RECT 9.445 1.857 9.455 2.028 ;
      RECT 9.395 1.842 9.445 2.018 ;
      RECT 9.345 1.817 9.395 1.998 ;
      RECT 9.335 1.802 9.345 1.98 ;
      RECT 9.33 1.8 9.335 1.974 ;
      RECT 9.31 1.795 9.33 1.969 ;
      RECT 9.305 1.787 9.31 1.963 ;
      RECT 9.29 1.781 9.305 1.956 ;
      RECT 9.285 1.776 9.29 1.948 ;
      RECT 9.265 1.771 9.285 1.94 ;
      RECT 9.25 1.764 9.265 1.933 ;
      RECT 9.235 1.758 9.25 1.924 ;
      RECT 9.23 1.752 9.235 1.917 ;
      RECT 9.185 1.727 9.23 1.903 ;
      RECT 9.17 1.697 9.185 1.885 ;
      RECT 9.155 1.68 9.17 1.876 ;
      RECT 9.13 1.66 9.155 1.864 ;
      RECT 9.09 1.63 9.13 1.844 ;
      RECT 9.08 1.6 9.09 1.829 ;
      RECT 9.065 1.59 9.08 1.822 ;
      RECT 9.01 1.555 9.065 1.801 ;
      RECT 8.995 1.518 9.01 1.78 ;
      RECT 8.985 1.505 8.995 1.772 ;
      RECT 8.935 1.475 8.985 1.754 ;
      RECT 8.92 1.405 8.935 1.735 ;
      RECT 8.875 1.405 8.92 1.718 ;
      RECT 8.85 1.405 8.875 1.7 ;
      RECT 8.84 1.405 8.85 1.693 ;
      RECT 8.761 1.405 8.84 1.686 ;
      RECT 8.675 1.405 8.761 1.678 ;
      RECT 8.66 1.437 8.675 1.673 ;
      RECT 8.585 1.447 8.66 1.669 ;
      RECT 8.565 1.457 8.585 1.664 ;
      RECT 8.54 1.457 8.565 1.661 ;
      RECT 8.53 1.447 8.54 1.66 ;
      RECT 8.52 1.42 8.53 1.659 ;
      RECT 8.48 1.415 8.52 1.657 ;
      RECT 8.435 1.415 8.48 1.653 ;
      RECT 8.41 1.415 8.435 1.648 ;
      RECT 8.36 1.415 8.41 1.635 ;
      RECT 8.32 1.42 8.33 1.62 ;
      RECT 8.33 1.415 8.36 1.625 ;
      RECT 10.315 1.195 10.575 1.455 ;
      RECT 10.31 1.217 10.575 1.413 ;
      RECT 9.55 1.045 9.77 1.41 ;
      RECT 9.532 1.132 9.77 1.409 ;
      RECT 9.515 1.137 9.77 1.406 ;
      RECT 9.515 1.137 9.79 1.405 ;
      RECT 9.485 1.147 9.79 1.403 ;
      RECT 9.48 1.162 9.79 1.399 ;
      RECT 9.48 1.162 9.795 1.398 ;
      RECT 9.475 1.22 9.795 1.396 ;
      RECT 9.475 1.22 9.805 1.393 ;
      RECT 9.47 1.285 9.805 1.388 ;
      RECT 9.55 1.045 9.81 1.305 ;
      RECT 8.295 0.875 8.555 1.135 ;
      RECT 8.295 0.918 8.641 1.109 ;
      RECT 8.295 0.918 8.685 1.108 ;
      RECT 8.295 0.918 8.705 1.106 ;
      RECT 8.295 0.918 8.805 1.105 ;
      RECT 8.295 0.918 8.825 1.103 ;
      RECT 8.295 0.918 8.835 1.098 ;
      RECT 8.705 0.885 8.895 1.095 ;
      RECT 8.705 0.887 8.9 1.093 ;
      RECT 8.695 0.892 8.905 1.085 ;
      RECT 8.641 0.916 8.905 1.085 ;
      RECT 8.685 0.91 8.695 1.107 ;
      RECT 8.695 0.89 8.9 1.093 ;
      RECT 7.65 1.95 7.855 2.18 ;
      RECT 7.59 1.9 7.645 2.16 ;
      RECT 7.65 1.9 7.85 2.18 ;
      RECT 8.62 2.215 8.625 2.242 ;
      RECT 8.61 2.125 8.62 2.247 ;
      RECT 8.605 2.047 8.61 2.253 ;
      RECT 8.595 2.037 8.605 2.26 ;
      RECT 8.59 2.027 8.595 2.266 ;
      RECT 8.58 2.022 8.59 2.268 ;
      RECT 8.565 2.014 8.58 2.276 ;
      RECT 8.55 2.005 8.565 2.288 ;
      RECT 8.54 1.997 8.55 2.298 ;
      RECT 8.505 1.915 8.54 2.316 ;
      RECT 8.47 1.915 8.505 2.335 ;
      RECT 8.455 1.915 8.47 2.343 ;
      RECT 8.4 1.915 8.455 2.343 ;
      RECT 8.366 1.915 8.4 2.334 ;
      RECT 8.28 1.915 8.366 2.31 ;
      RECT 8.27 1.975 8.28 2.292 ;
      RECT 8.23 1.977 8.27 2.283 ;
      RECT 8.225 1.979 8.23 2.273 ;
      RECT 8.205 1.981 8.225 2.268 ;
      RECT 8.195 1.984 8.205 2.263 ;
      RECT 8.185 1.985 8.195 2.258 ;
      RECT 8.161 1.986 8.185 2.25 ;
      RECT 8.075 1.991 8.161 2.228 ;
      RECT 8.02 1.99 8.075 2.201 ;
      RECT 8.005 1.983 8.02 2.188 ;
      RECT 7.97 1.978 8.005 2.184 ;
      RECT 7.915 1.97 7.97 2.183 ;
      RECT 7.855 1.957 7.915 2.181 ;
      RECT 7.645 1.9 7.65 2.168 ;
      RECT 7.72 1.27 7.905 1.48 ;
      RECT 7.71 1.275 7.92 1.473 ;
      RECT 7.75 1.18 8.01 1.44 ;
      RECT 7.705 1.337 8.01 1.363 ;
      RECT 7.05 1.13 7.055 1.93 ;
      RECT 6.995 1.18 7.025 1.93 ;
      RECT 6.985 1.18 6.99 1.49 ;
      RECT 6.97 1.18 6.975 1.485 ;
      RECT 6.515 1.225 6.53 1.44 ;
      RECT 6.445 1.225 6.53 1.435 ;
      RECT 7.71 0.805 7.78 1.015 ;
      RECT 7.78 0.812 7.79 1.01 ;
      RECT 7.676 0.805 7.71 1.022 ;
      RECT 7.59 0.805 7.676 1.046 ;
      RECT 7.58 0.81 7.59 1.065 ;
      RECT 7.575 0.822 7.58 1.068 ;
      RECT 7.56 0.837 7.575 1.072 ;
      RECT 7.555 0.855 7.56 1.076 ;
      RECT 7.515 0.865 7.555 1.085 ;
      RECT 7.5 0.872 7.515 1.097 ;
      RECT 7.485 0.877 7.5 1.102 ;
      RECT 7.47 0.88 7.485 1.107 ;
      RECT 7.46 0.882 7.47 1.111 ;
      RECT 7.425 0.889 7.46 1.119 ;
      RECT 7.39 0.897 7.425 1.133 ;
      RECT 7.38 0.903 7.39 1.142 ;
      RECT 7.375 0.905 7.38 1.144 ;
      RECT 7.355 0.908 7.375 1.15 ;
      RECT 7.325 0.915 7.355 1.161 ;
      RECT 7.315 0.921 7.325 1.168 ;
      RECT 7.29 0.924 7.315 1.175 ;
      RECT 7.28 0.928 7.29 1.183 ;
      RECT 7.275 0.929 7.28 1.205 ;
      RECT 7.27 0.93 7.275 1.22 ;
      RECT 7.265 0.931 7.27 1.235 ;
      RECT 7.26 0.932 7.265 1.25 ;
      RECT 7.255 0.933 7.26 1.28 ;
      RECT 7.245 0.935 7.255 1.313 ;
      RECT 7.23 0.939 7.245 1.36 ;
      RECT 7.22 0.942 7.23 1.405 ;
      RECT 7.215 0.945 7.22 1.433 ;
      RECT 7.205 0.947 7.215 1.46 ;
      RECT 7.2 0.95 7.205 1.495 ;
      RECT 7.17 0.955 7.2 1.553 ;
      RECT 7.165 0.96 7.17 1.638 ;
      RECT 7.16 0.962 7.165 1.673 ;
      RECT 7.155 0.964 7.16 1.755 ;
      RECT 7.15 0.966 7.155 1.843 ;
      RECT 7.14 0.968 7.15 1.925 ;
      RECT 7.125 0.982 7.14 1.93 ;
      RECT 7.09 1.027 7.125 1.93 ;
      RECT 7.08 1.067 7.09 1.93 ;
      RECT 7.065 1.095 7.08 1.93 ;
      RECT 7.06 1.112 7.065 1.93 ;
      RECT 7.055 1.12 7.06 1.93 ;
      RECT 7.045 1.135 7.05 1.93 ;
      RECT 7.04 1.142 7.045 1.93 ;
      RECT 7.03 1.162 7.04 1.93 ;
      RECT 7.025 1.175 7.03 1.93 ;
      RECT 6.99 1.18 6.995 1.515 ;
      RECT 6.975 1.57 6.995 1.93 ;
      RECT 6.975 1.18 6.985 1.488 ;
      RECT 6.97 1.61 6.975 1.93 ;
      RECT 6.92 1.18 6.97 1.483 ;
      RECT 6.965 1.647 6.97 1.93 ;
      RECT 6.955 1.67 6.965 1.93 ;
      RECT 6.95 1.715 6.955 1.93 ;
      RECT 6.94 1.725 6.95 1.923 ;
      RECT 6.866 1.18 6.92 1.477 ;
      RECT 6.78 1.18 6.866 1.47 ;
      RECT 6.731 1.227 6.78 1.463 ;
      RECT 6.645 1.235 6.731 1.456 ;
      RECT 6.63 1.232 6.645 1.451 ;
      RECT 6.616 1.225 6.63 1.45 ;
      RECT 6.53 1.225 6.616 1.445 ;
      RECT 6.435 1.23 6.445 1.43 ;
      RECT 6.025 0.66 6.04 1.06 ;
      RECT 6.22 0.66 6.225 0.92 ;
      RECT 5.965 0.66 6.01 0.92 ;
      RECT 6.42 1.965 6.425 2.17 ;
      RECT 6.415 1.955 6.42 2.175 ;
      RECT 6.41 1.942 6.415 2.18 ;
      RECT 6.405 1.922 6.41 2.18 ;
      RECT 6.38 1.875 6.405 2.18 ;
      RECT 6.345 1.79 6.38 2.18 ;
      RECT 6.34 1.727 6.345 2.18 ;
      RECT 6.335 1.712 6.34 2.18 ;
      RECT 6.32 1.672 6.335 2.18 ;
      RECT 6.315 1.647 6.32 2.18 ;
      RECT 6.305 1.63 6.315 2.18 ;
      RECT 6.27 1.552 6.305 2.18 ;
      RECT 6.265 1.495 6.27 2.18 ;
      RECT 6.26 1.482 6.265 2.18 ;
      RECT 6.25 1.46 6.26 2.18 ;
      RECT 6.24 1.425 6.25 2.18 ;
      RECT 6.23 1.395 6.24 2.18 ;
      RECT 6.22 1.31 6.23 1.823 ;
      RECT 6.227 1.955 6.23 2.18 ;
      RECT 6.225 1.965 6.227 2.18 ;
      RECT 6.215 1.975 6.225 2.175 ;
      RECT 6.21 0.66 6.22 1.055 ;
      RECT 6.215 1.187 6.22 1.798 ;
      RECT 6.21 1.085 6.215 1.781 ;
      RECT 6.2 0.66 6.21 1.757 ;
      RECT 6.195 0.66 6.2 1.728 ;
      RECT 6.19 0.66 6.195 1.718 ;
      RECT 6.17 0.66 6.19 1.68 ;
      RECT 6.165 0.66 6.17 1.638 ;
      RECT 6.16 0.66 6.165 1.618 ;
      RECT 6.13 0.66 6.16 1.568 ;
      RECT 6.12 0.66 6.13 1.515 ;
      RECT 6.115 0.66 6.12 1.488 ;
      RECT 6.11 0.66 6.115 1.473 ;
      RECT 6.1 0.66 6.11 1.45 ;
      RECT 6.09 0.66 6.1 1.425 ;
      RECT 6.085 0.66 6.09 1.365 ;
      RECT 6.075 0.66 6.085 1.303 ;
      RECT 6.07 0.66 6.075 1.223 ;
      RECT 6.065 0.66 6.07 1.188 ;
      RECT 6.06 0.66 6.065 1.163 ;
      RECT 6.055 0.66 6.06 1.148 ;
      RECT 6.05 0.66 6.055 1.118 ;
      RECT 6.045 0.66 6.05 1.095 ;
      RECT 6.04 0.66 6.045 1.068 ;
      RECT 6.01 0.66 6.025 1.055 ;
      RECT 5.165 2.195 5.35 2.405 ;
      RECT 5.155 2.2 5.365 2.398 ;
      RECT 5.155 2.2 5.385 2.37 ;
      RECT 5.155 2.2 5.4 2.349 ;
      RECT 5.155 2.2 5.415 2.347 ;
      RECT 5.155 2.2 5.425 2.346 ;
      RECT 5.155 2.2 5.455 2.343 ;
      RECT 5.805 2.045 6.065 2.305 ;
      RECT 5.765 2.092 6.065 2.288 ;
      RECT 5.756 2.1 5.765 2.291 ;
      RECT 5.35 2.193 6.065 2.288 ;
      RECT 5.67 2.118 5.756 2.298 ;
      RECT 5.365 2.19 6.065 2.288 ;
      RECT 5.611 2.14 5.67 2.31 ;
      RECT 5.385 2.186 6.065 2.288 ;
      RECT 5.525 2.152 5.611 2.321 ;
      RECT 5.4 2.182 6.065 2.288 ;
      RECT 5.47 2.165 5.525 2.333 ;
      RECT 5.415 2.18 6.065 2.288 ;
      RECT 5.455 2.171 5.47 2.339 ;
      RECT 5.425 2.176 6.065 2.288 ;
      RECT 5.57 1.7 5.83 1.96 ;
      RECT 5.57 1.72 5.94 1.93 ;
      RECT 5.57 1.725 5.95 1.925 ;
      RECT 5.761 1.139 5.84 1.37 ;
      RECT 5.675 1.142 5.89 1.365 ;
      RECT 5.67 1.142 5.89 1.36 ;
      RECT 5.67 1.147 5.9 1.358 ;
      RECT 5.645 1.147 5.9 1.355 ;
      RECT 5.645 1.155 5.91 1.353 ;
      RECT 5.525 1.09 5.785 1.35 ;
      RECT 5.525 1.137 5.835 1.35 ;
      RECT 4.78 1.71 4.785 1.97 ;
      RECT 4.61 1.48 4.615 1.97 ;
      RECT 4.495 1.72 4.5 1.945 ;
      RECT 5.205 0.815 5.21 1.025 ;
      RECT 5.21 0.82 5.225 1.02 ;
      RECT 5.145 0.815 5.205 1.033 ;
      RECT 5.13 0.815 5.145 1.043 ;
      RECT 5.08 0.815 5.13 1.06 ;
      RECT 5.06 0.815 5.08 1.083 ;
      RECT 5.045 0.815 5.06 1.095 ;
      RECT 5.025 0.815 5.045 1.105 ;
      RECT 5.015 0.82 5.025 1.114 ;
      RECT 5.01 0.83 5.015 1.119 ;
      RECT 5.005 0.842 5.01 1.123 ;
      RECT 4.995 0.865 5.005 1.128 ;
      RECT 4.99 0.88 4.995 1.132 ;
      RECT 4.985 0.897 4.99 1.135 ;
      RECT 4.98 0.905 4.985 1.138 ;
      RECT 4.97 0.91 4.98 1.142 ;
      RECT 4.965 0.917 4.97 1.147 ;
      RECT 4.955 0.922 4.965 1.151 ;
      RECT 4.93 0.934 4.955 1.162 ;
      RECT 4.91 0.951 4.93 1.178 ;
      RECT 4.885 0.968 4.91 1.2 ;
      RECT 4.85 0.991 4.885 1.258 ;
      RECT 4.83 1.013 4.85 1.32 ;
      RECT 4.825 1.023 4.83 1.355 ;
      RECT 4.815 1.03 4.825 1.393 ;
      RECT 4.81 1.037 4.815 1.413 ;
      RECT 4.805 1.048 4.81 1.45 ;
      RECT 4.8 1.056 4.805 1.515 ;
      RECT 4.79 1.067 4.8 1.568 ;
      RECT 4.785 1.085 4.79 1.638 ;
      RECT 4.78 1.095 4.785 1.675 ;
      RECT 4.775 1.105 4.78 1.97 ;
      RECT 4.77 1.117 4.775 1.97 ;
      RECT 4.765 1.127 4.77 1.97 ;
      RECT 4.755 1.137 4.765 1.97 ;
      RECT 4.745 1.16 4.755 1.97 ;
      RECT 4.73 1.195 4.745 1.97 ;
      RECT 4.69 1.257 4.73 1.97 ;
      RECT 4.685 1.31 4.69 1.97 ;
      RECT 4.66 1.345 4.685 1.97 ;
      RECT 4.645 1.39 4.66 1.97 ;
      RECT 4.64 1.412 4.645 1.97 ;
      RECT 4.63 1.425 4.64 1.97 ;
      RECT 4.62 1.45 4.63 1.97 ;
      RECT 4.615 1.472 4.62 1.97 ;
      RECT 4.59 1.51 4.61 1.97 ;
      RECT 4.55 1.567 4.59 1.97 ;
      RECT 4.545 1.617 4.55 1.97 ;
      RECT 4.54 1.635 4.545 1.97 ;
      RECT 4.535 1.647 4.54 1.97 ;
      RECT 4.525 1.665 4.535 1.97 ;
      RECT 4.515 1.685 4.525 1.945 ;
      RECT 4.51 1.702 4.515 1.945 ;
      RECT 4.5 1.715 4.51 1.945 ;
      RECT 4.47 1.725 4.495 1.945 ;
      RECT 4.46 1.732 4.47 1.945 ;
      RECT 4.445 1.742 4.46 1.94 ;
      RECT 3.405 1.655 3.725 1.915 ;
      RECT 3.27 1.7 3.725 1.87 ;
      RECT -3.835 1.78 -3.545 2.02 ;
      RECT -3.775 1.595 -3.6 2.02 ;
      RECT -3.77 1.135 -3.6 2.02 ;
      RECT -3.77 1.135 2.81 1.305 ;
      RECT 2.64 0.715 2.81 1.305 ;
      RECT 2.55 0.715 2.87 0.975 ;
      RECT 2.55 0.745 2.95 0.915 ;
      RECT 0.215 1.755 0.51 2.045 ;
      RECT 0.185 1.755 0.51 2.015 ;
      RECT -3.95 0 138.165 0.48 ;
      RECT 134.745 0.845 135.075 1.115 ;
      RECT 130.865 0.785 131.185 1.045 ;
      RECT 126.325 0.725 126.645 0.985 ;
      RECT 103.27 0.785 103.59 1.045 ;
      RECT 98.73 0.725 99.05 0.985 ;
      RECT 75.675 0.785 75.995 1.045 ;
      RECT 71.135 0.725 71.455 0.985 ;
      RECT 48.08 0.785 48.4 1.045 ;
      RECT 43.54 0.725 43.86 0.985 ;
      RECT 20.485 0.785 20.805 1.045 ;
      RECT 15.945 0.725 16.265 0.985 ;
      RECT -2 0.65 -1.68 0.91 ;
    LAYER mcon ;
      RECT 137.85 0.155 138.02 0.325 ;
      RECT 137.85 2.875 138.02 3.045 ;
      RECT 137.39 0.155 137.56 0.325 ;
      RECT 137.39 2.875 137.56 3.045 ;
      RECT 136.93 0.155 137.1 0.325 ;
      RECT 136.93 2.875 137.1 3.045 ;
      RECT 136.47 0.155 136.64 0.325 ;
      RECT 136.47 2.875 136.64 3.045 ;
      RECT 136.01 0.155 136.18 0.325 ;
      RECT 136.01 2.875 136.18 3.045 ;
      RECT 135.805 1.34 135.975 1.51 ;
      RECT 135.55 0.155 135.72 0.325 ;
      RECT 135.55 2.875 135.72 3.045 ;
      RECT 135.09 0.155 135.26 0.325 ;
      RECT 135.09 2.875 135.26 3.045 ;
      RECT 134.825 0.895 134.995 1.065 ;
      RECT 134.63 0.155 134.8 0.325 ;
      RECT 134.63 2.875 134.8 3.045 ;
      RECT 134.17 0.155 134.34 0.325 ;
      RECT 134.17 2.875 134.34 3.045 ;
      RECT 133.71 0.155 133.88 0.325 ;
      RECT 133.71 2.875 133.88 3.045 ;
      RECT 133.25 0.155 133.42 0.325 ;
      RECT 133.25 2.875 133.42 3.045 ;
      RECT 133.045 1.345 133.215 1.515 ;
      RECT 132.79 0.155 132.96 0.325 ;
      RECT 132.79 2.875 132.96 3.045 ;
      RECT 132.33 0.155 132.5 0.325 ;
      RECT 132.33 2.875 132.5 3.045 ;
      RECT 131.87 0.155 132.04 0.325 ;
      RECT 131.87 2.875 132.04 3.045 ;
      RECT 131.8 1.7 131.97 1.87 ;
      RECT 131.41 0.155 131.58 0.325 ;
      RECT 131.41 2.875 131.58 3.045 ;
      RECT 130.95 0.155 131.12 0.325 ;
      RECT 130.95 2.875 131.12 3.045 ;
      RECT 130.94 0.815 131.11 0.985 ;
      RECT 130.495 0.695 130.665 0.865 ;
      RECT 130.49 0.155 130.66 0.325 ;
      RECT 130.49 2.875 130.66 3.045 ;
      RECT 130.03 0.155 130.2 0.325 ;
      RECT 130.03 2.875 130.2 3.045 ;
      RECT 129.57 0.155 129.74 0.325 ;
      RECT 129.57 2.875 129.74 3.045 ;
      RECT 129.11 0.155 129.28 0.325 ;
      RECT 129.11 2.875 129.28 3.045 ;
      RECT 128.65 0.155 128.82 0.325 ;
      RECT 128.65 2.875 128.82 3.045 ;
      RECT 128.595 1.315 128.765 1.485 ;
      RECT 128.195 0.155 128.365 0.325 ;
      RECT 128.195 2.875 128.365 3.045 ;
      RECT 127.735 0.155 127.905 0.325 ;
      RECT 127.735 2.875 127.905 3.045 ;
      RECT 127.665 1.7 127.835 1.87 ;
      RECT 127.275 0.155 127.445 0.325 ;
      RECT 127.275 2.875 127.445 3.045 ;
      RECT 126.815 0.155 126.985 0.325 ;
      RECT 126.815 2.875 126.985 3.045 ;
      RECT 126.4 0.755 126.57 0.925 ;
      RECT 126.355 0.155 126.525 0.325 ;
      RECT 126.355 2.875 126.525 3.045 ;
      RECT 125.985 1.48 126.155 1.65 ;
      RECT 125.895 0.155 126.065 0.325 ;
      RECT 125.895 2.875 126.065 3.045 ;
      RECT 125.435 0.155 125.605 0.325 ;
      RECT 125.435 2.875 125.605 3.045 ;
      RECT 124.975 0.155 125.145 0.325 ;
      RECT 124.975 2.875 125.145 3.045 ;
      RECT 124.515 0.155 124.685 0.325 ;
      RECT 124.515 2.875 124.685 3.045 ;
      RECT 124.46 2.155 124.63 2.325 ;
      RECT 124.055 0.155 124.225 0.325 ;
      RECT 124.055 2.875 124.225 3.045 ;
      RECT 123.685 1.615 123.855 1.785 ;
      RECT 123.595 0.155 123.765 0.325 ;
      RECT 123.595 2.875 123.765 3.045 ;
      RECT 123.365 0.785 123.535 0.955 ;
      RECT 123.22 1.225 123.39 1.395 ;
      RECT 123.135 0.155 123.305 0.325 ;
      RECT 123.135 2.875 123.305 3.045 ;
      RECT 122.675 0.155 122.845 0.325 ;
      RECT 122.675 2.875 122.845 3.045 ;
      RECT 122.61 1.265 122.78 1.435 ;
      RECT 122.265 0.9 122.435 1.07 ;
      RECT 122.255 2.26 122.425 2.43 ;
      RECT 122.215 0.155 122.385 0.325 ;
      RECT 122.215 2.875 122.385 3.045 ;
      RECT 121.84 1.5 122.01 1.67 ;
      RECT 121.755 0.155 121.925 0.325 ;
      RECT 121.755 2.875 121.925 3.045 ;
      RECT 121.49 0.975 121.66 1.145 ;
      RECT 121.31 2.29 121.48 2.46 ;
      RECT 121.295 0.155 121.465 0.325 ;
      RECT 121.295 2.875 121.465 3.045 ;
      RECT 121.03 1.605 121.2 1.775 ;
      RECT 120.835 0.155 121.005 0.325 ;
      RECT 120.835 2.875 121.005 3.045 ;
      RECT 120.71 1.23 120.88 1.4 ;
      RECT 120.375 0.155 120.545 0.325 ;
      RECT 120.375 2.875 120.545 3.045 ;
      RECT 120.02 0.71 120.19 0.88 ;
      RECT 119.945 1.18 120.115 1.35 ;
      RECT 119.915 0.155 120.085 0.325 ;
      RECT 119.915 2.875 120.085 3.045 ;
      RECT 119.455 0.155 119.625 0.325 ;
      RECT 119.455 2.875 119.625 3.045 ;
      RECT 119.095 0.905 119.265 1.075 ;
      RECT 118.995 0.155 119.165 0.325 ;
      RECT 118.995 2.875 119.165 3.045 ;
      RECT 118.755 2.1 118.925 2.27 ;
      RECT 118.72 1.435 118.89 1.605 ;
      RECT 118.535 0.155 118.705 0.325 ;
      RECT 118.535 2.875 118.705 3.045 ;
      RECT 118.11 1.29 118.28 1.46 ;
      RECT 118.075 0.155 118.245 0.325 ;
      RECT 118.075 2.875 118.245 3.045 ;
      RECT 118.04 1.99 118.21 2.16 ;
      RECT 117.98 0.825 118.15 0.995 ;
      RECT 117.615 0.155 117.785 0.325 ;
      RECT 117.615 2.875 117.785 3.045 ;
      RECT 117.34 1.74 117.51 1.91 ;
      RECT 117.155 0.155 117.325 0.325 ;
      RECT 117.155 2.875 117.325 3.045 ;
      RECT 116.835 1.245 117.005 1.415 ;
      RECT 116.695 0.155 116.865 0.325 ;
      RECT 116.695 2.875 116.865 3.045 ;
      RECT 116.615 1.99 116.785 2.16 ;
      RECT 116.41 0.87 116.58 1.04 ;
      RECT 116.235 0.155 116.405 0.325 ;
      RECT 116.235 2.875 116.405 3.045 ;
      RECT 116.14 1.74 116.31 1.91 ;
      RECT 116.1 1.17 116.27 1.34 ;
      RECT 115.775 0.155 115.945 0.325 ;
      RECT 115.775 2.875 115.945 3.045 ;
      RECT 115.555 2.215 115.725 2.385 ;
      RECT 115.415 0.835 115.585 1.005 ;
      RECT 115.315 0.155 115.485 0.325 ;
      RECT 115.315 2.875 115.485 3.045 ;
      RECT 114.855 0.155 115.025 0.325 ;
      RECT 114.855 2.875 115.025 3.045 ;
      RECT 114.845 1.755 115.015 1.925 ;
      RECT 114.395 0.155 114.565 0.325 ;
      RECT 114.395 2.875 114.565 3.045 ;
      RECT 113.935 0.155 114.105 0.325 ;
      RECT 113.935 2.875 114.105 3.045 ;
      RECT 113.865 1.7 114.035 1.87 ;
      RECT 113.475 0.155 113.645 0.325 ;
      RECT 113.475 2.875 113.645 3.045 ;
      RECT 113.015 0.155 113.185 0.325 ;
      RECT 113.015 2.875 113.185 3.045 ;
      RECT 113.005 0.745 113.175 0.915 ;
      RECT 112.555 0.155 112.725 0.325 ;
      RECT 112.555 2.875 112.725 3.045 ;
      RECT 112.095 0.155 112.265 0.325 ;
      RECT 112.095 2.875 112.265 3.045 ;
      RECT 111.635 0.155 111.805 0.325 ;
      RECT 111.635 2.875 111.805 3.045 ;
      RECT 111.175 0.155 111.345 0.325 ;
      RECT 111.175 2.875 111.345 3.045 ;
      RECT 110.715 0.155 110.885 0.325 ;
      RECT 110.715 2.875 110.885 3.045 ;
      RECT 110.66 1.815 110.83 1.985 ;
      RECT 110.255 0.155 110.425 0.325 ;
      RECT 110.255 2.875 110.425 3.045 ;
      RECT 109.795 0.155 109.965 0.325 ;
      RECT 109.795 2.875 109.965 3.045 ;
      RECT 109.335 0.155 109.505 0.325 ;
      RECT 109.335 2.875 109.505 3.045 ;
      RECT 108.875 0.155 109.045 0.325 ;
      RECT 108.875 2.875 109.045 3.045 ;
      RECT 108.415 0.155 108.585 0.325 ;
      RECT 108.415 2.875 108.585 3.045 ;
      RECT 108.21 1.34 108.38 1.51 ;
      RECT 107.955 0.155 108.125 0.325 ;
      RECT 107.955 2.875 108.125 3.045 ;
      RECT 107.495 0.155 107.665 0.325 ;
      RECT 107.495 2.875 107.665 3.045 ;
      RECT 107.25 1.555 107.42 1.725 ;
      RECT 107.035 0.155 107.205 0.325 ;
      RECT 107.035 2.875 107.205 3.045 ;
      RECT 106.575 0.155 106.745 0.325 ;
      RECT 106.575 2.875 106.745 3.045 ;
      RECT 106.115 0.155 106.285 0.325 ;
      RECT 106.115 2.875 106.285 3.045 ;
      RECT 105.655 0.155 105.825 0.325 ;
      RECT 105.655 2.875 105.825 3.045 ;
      RECT 105.45 1.345 105.62 1.515 ;
      RECT 105.195 0.155 105.365 0.325 ;
      RECT 105.195 2.875 105.365 3.045 ;
      RECT 104.735 0.155 104.905 0.325 ;
      RECT 104.735 2.875 104.905 3.045 ;
      RECT 104.275 0.155 104.445 0.325 ;
      RECT 104.275 2.875 104.445 3.045 ;
      RECT 104.205 1.7 104.375 1.87 ;
      RECT 103.815 0.155 103.985 0.325 ;
      RECT 103.815 2.875 103.985 3.045 ;
      RECT 103.355 0.155 103.525 0.325 ;
      RECT 103.355 2.875 103.525 3.045 ;
      RECT 103.345 0.815 103.515 0.985 ;
      RECT 102.9 0.695 103.07 0.865 ;
      RECT 102.895 0.155 103.065 0.325 ;
      RECT 102.895 2.875 103.065 3.045 ;
      RECT 102.435 0.155 102.605 0.325 ;
      RECT 102.435 2.875 102.605 3.045 ;
      RECT 101.975 0.155 102.145 0.325 ;
      RECT 101.975 2.875 102.145 3.045 ;
      RECT 101.515 0.155 101.685 0.325 ;
      RECT 101.515 2.875 101.685 3.045 ;
      RECT 101.055 0.155 101.225 0.325 ;
      RECT 101.055 2.875 101.225 3.045 ;
      RECT 101 1.315 101.17 1.485 ;
      RECT 100.6 0.155 100.77 0.325 ;
      RECT 100.6 2.875 100.77 3.045 ;
      RECT 100.14 0.155 100.31 0.325 ;
      RECT 100.14 2.875 100.31 3.045 ;
      RECT 100.07 1.7 100.24 1.87 ;
      RECT 99.68 0.155 99.85 0.325 ;
      RECT 99.68 2.875 99.85 3.045 ;
      RECT 99.22 0.155 99.39 0.325 ;
      RECT 99.22 2.875 99.39 3.045 ;
      RECT 98.805 0.755 98.975 0.925 ;
      RECT 98.76 0.155 98.93 0.325 ;
      RECT 98.76 2.875 98.93 3.045 ;
      RECT 98.39 1.48 98.56 1.65 ;
      RECT 98.3 0.155 98.47 0.325 ;
      RECT 98.3 2.875 98.47 3.045 ;
      RECT 97.84 0.155 98.01 0.325 ;
      RECT 97.84 2.875 98.01 3.045 ;
      RECT 97.38 0.155 97.55 0.325 ;
      RECT 97.38 2.875 97.55 3.045 ;
      RECT 96.92 0.155 97.09 0.325 ;
      RECT 96.92 2.875 97.09 3.045 ;
      RECT 96.865 2.155 97.035 2.325 ;
      RECT 96.46 0.155 96.63 0.325 ;
      RECT 96.46 2.875 96.63 3.045 ;
      RECT 96.09 1.615 96.26 1.785 ;
      RECT 96 0.155 96.17 0.325 ;
      RECT 96 2.875 96.17 3.045 ;
      RECT 95.77 0.785 95.94 0.955 ;
      RECT 95.625 1.225 95.795 1.395 ;
      RECT 95.54 0.155 95.71 0.325 ;
      RECT 95.54 2.875 95.71 3.045 ;
      RECT 95.08 0.155 95.25 0.325 ;
      RECT 95.08 2.875 95.25 3.045 ;
      RECT 95.015 1.265 95.185 1.435 ;
      RECT 94.67 0.9 94.84 1.07 ;
      RECT 94.66 2.26 94.83 2.43 ;
      RECT 94.62 0.155 94.79 0.325 ;
      RECT 94.62 2.875 94.79 3.045 ;
      RECT 94.245 1.5 94.415 1.67 ;
      RECT 94.16 0.155 94.33 0.325 ;
      RECT 94.16 2.875 94.33 3.045 ;
      RECT 93.895 0.975 94.065 1.145 ;
      RECT 93.715 2.29 93.885 2.46 ;
      RECT 93.7 0.155 93.87 0.325 ;
      RECT 93.7 2.875 93.87 3.045 ;
      RECT 93.435 1.605 93.605 1.775 ;
      RECT 93.24 0.155 93.41 0.325 ;
      RECT 93.24 2.875 93.41 3.045 ;
      RECT 93.115 1.23 93.285 1.4 ;
      RECT 92.78 0.155 92.95 0.325 ;
      RECT 92.78 2.875 92.95 3.045 ;
      RECT 92.425 0.71 92.595 0.88 ;
      RECT 92.35 1.18 92.52 1.35 ;
      RECT 92.32 0.155 92.49 0.325 ;
      RECT 92.32 2.875 92.49 3.045 ;
      RECT 91.86 0.155 92.03 0.325 ;
      RECT 91.86 2.875 92.03 3.045 ;
      RECT 91.5 0.905 91.67 1.075 ;
      RECT 91.4 0.155 91.57 0.325 ;
      RECT 91.4 2.875 91.57 3.045 ;
      RECT 91.16 2.1 91.33 2.27 ;
      RECT 91.125 1.435 91.295 1.605 ;
      RECT 90.94 0.155 91.11 0.325 ;
      RECT 90.94 2.875 91.11 3.045 ;
      RECT 90.515 1.29 90.685 1.46 ;
      RECT 90.48 0.155 90.65 0.325 ;
      RECT 90.48 2.875 90.65 3.045 ;
      RECT 90.445 1.99 90.615 2.16 ;
      RECT 90.385 0.825 90.555 0.995 ;
      RECT 90.02 0.155 90.19 0.325 ;
      RECT 90.02 2.875 90.19 3.045 ;
      RECT 89.745 1.74 89.915 1.91 ;
      RECT 89.56 0.155 89.73 0.325 ;
      RECT 89.56 2.875 89.73 3.045 ;
      RECT 89.24 1.245 89.41 1.415 ;
      RECT 89.1 0.155 89.27 0.325 ;
      RECT 89.1 2.875 89.27 3.045 ;
      RECT 89.02 1.99 89.19 2.16 ;
      RECT 88.815 0.87 88.985 1.04 ;
      RECT 88.64 0.155 88.81 0.325 ;
      RECT 88.64 2.875 88.81 3.045 ;
      RECT 88.545 1.74 88.715 1.91 ;
      RECT 88.505 1.17 88.675 1.34 ;
      RECT 88.18 0.155 88.35 0.325 ;
      RECT 88.18 2.875 88.35 3.045 ;
      RECT 87.96 2.215 88.13 2.385 ;
      RECT 87.82 0.835 87.99 1.005 ;
      RECT 87.72 0.155 87.89 0.325 ;
      RECT 87.72 2.875 87.89 3.045 ;
      RECT 87.26 0.155 87.43 0.325 ;
      RECT 87.26 2.875 87.43 3.045 ;
      RECT 87.25 1.755 87.42 1.925 ;
      RECT 86.8 0.155 86.97 0.325 ;
      RECT 86.8 2.875 86.97 3.045 ;
      RECT 86.34 0.155 86.51 0.325 ;
      RECT 86.34 2.875 86.51 3.045 ;
      RECT 86.27 1.7 86.44 1.87 ;
      RECT 85.88 0.155 86.05 0.325 ;
      RECT 85.88 2.875 86.05 3.045 ;
      RECT 85.42 0.155 85.59 0.325 ;
      RECT 85.42 2.875 85.59 3.045 ;
      RECT 85.41 0.745 85.58 0.915 ;
      RECT 84.96 0.155 85.13 0.325 ;
      RECT 84.96 2.875 85.13 3.045 ;
      RECT 84.5 0.155 84.67 0.325 ;
      RECT 84.5 2.875 84.67 3.045 ;
      RECT 84.04 0.155 84.21 0.325 ;
      RECT 84.04 2.875 84.21 3.045 ;
      RECT 83.58 0.155 83.75 0.325 ;
      RECT 83.58 2.875 83.75 3.045 ;
      RECT 83.12 0.155 83.29 0.325 ;
      RECT 83.12 2.875 83.29 3.045 ;
      RECT 83.065 1.815 83.235 1.985 ;
      RECT 82.66 0.155 82.83 0.325 ;
      RECT 82.66 2.875 82.83 3.045 ;
      RECT 82.2 0.155 82.37 0.325 ;
      RECT 82.2 2.875 82.37 3.045 ;
      RECT 81.74 0.155 81.91 0.325 ;
      RECT 81.74 2.875 81.91 3.045 ;
      RECT 81.28 0.155 81.45 0.325 ;
      RECT 81.28 2.875 81.45 3.045 ;
      RECT 80.82 0.155 80.99 0.325 ;
      RECT 80.82 2.875 80.99 3.045 ;
      RECT 80.615 1.34 80.785 1.51 ;
      RECT 80.36 0.155 80.53 0.325 ;
      RECT 80.36 2.875 80.53 3.045 ;
      RECT 79.9 0.155 80.07 0.325 ;
      RECT 79.9 2.875 80.07 3.045 ;
      RECT 79.655 1.555 79.825 1.725 ;
      RECT 79.44 0.155 79.61 0.325 ;
      RECT 79.44 2.875 79.61 3.045 ;
      RECT 78.98 0.155 79.15 0.325 ;
      RECT 78.98 2.875 79.15 3.045 ;
      RECT 78.52 0.155 78.69 0.325 ;
      RECT 78.52 2.875 78.69 3.045 ;
      RECT 78.06 0.155 78.23 0.325 ;
      RECT 78.06 2.875 78.23 3.045 ;
      RECT 77.855 1.345 78.025 1.515 ;
      RECT 77.6 0.155 77.77 0.325 ;
      RECT 77.6 2.875 77.77 3.045 ;
      RECT 77.14 0.155 77.31 0.325 ;
      RECT 77.14 2.875 77.31 3.045 ;
      RECT 76.68 0.155 76.85 0.325 ;
      RECT 76.68 2.875 76.85 3.045 ;
      RECT 76.61 1.7 76.78 1.87 ;
      RECT 76.22 0.155 76.39 0.325 ;
      RECT 76.22 2.875 76.39 3.045 ;
      RECT 75.76 0.155 75.93 0.325 ;
      RECT 75.76 2.875 75.93 3.045 ;
      RECT 75.75 0.815 75.92 0.985 ;
      RECT 75.305 0.695 75.475 0.865 ;
      RECT 75.3 0.155 75.47 0.325 ;
      RECT 75.3 2.875 75.47 3.045 ;
      RECT 74.84 0.155 75.01 0.325 ;
      RECT 74.84 2.875 75.01 3.045 ;
      RECT 74.38 0.155 74.55 0.325 ;
      RECT 74.38 2.875 74.55 3.045 ;
      RECT 73.92 0.155 74.09 0.325 ;
      RECT 73.92 2.875 74.09 3.045 ;
      RECT 73.46 0.155 73.63 0.325 ;
      RECT 73.46 2.875 73.63 3.045 ;
      RECT 73.405 1.315 73.575 1.485 ;
      RECT 73.005 0.155 73.175 0.325 ;
      RECT 73.005 2.875 73.175 3.045 ;
      RECT 72.545 0.155 72.715 0.325 ;
      RECT 72.545 2.875 72.715 3.045 ;
      RECT 72.475 1.7 72.645 1.87 ;
      RECT 72.085 0.155 72.255 0.325 ;
      RECT 72.085 2.875 72.255 3.045 ;
      RECT 71.625 0.155 71.795 0.325 ;
      RECT 71.625 2.875 71.795 3.045 ;
      RECT 71.21 0.755 71.38 0.925 ;
      RECT 71.165 0.155 71.335 0.325 ;
      RECT 71.165 2.875 71.335 3.045 ;
      RECT 70.795 1.48 70.965 1.65 ;
      RECT 70.705 0.155 70.875 0.325 ;
      RECT 70.705 2.875 70.875 3.045 ;
      RECT 70.245 0.155 70.415 0.325 ;
      RECT 70.245 2.875 70.415 3.045 ;
      RECT 69.785 0.155 69.955 0.325 ;
      RECT 69.785 2.875 69.955 3.045 ;
      RECT 69.325 0.155 69.495 0.325 ;
      RECT 69.325 2.875 69.495 3.045 ;
      RECT 69.27 2.155 69.44 2.325 ;
      RECT 68.865 0.155 69.035 0.325 ;
      RECT 68.865 2.875 69.035 3.045 ;
      RECT 68.495 1.615 68.665 1.785 ;
      RECT 68.405 0.155 68.575 0.325 ;
      RECT 68.405 2.875 68.575 3.045 ;
      RECT 68.175 0.785 68.345 0.955 ;
      RECT 68.03 1.225 68.2 1.395 ;
      RECT 67.945 0.155 68.115 0.325 ;
      RECT 67.945 2.875 68.115 3.045 ;
      RECT 67.485 0.155 67.655 0.325 ;
      RECT 67.485 2.875 67.655 3.045 ;
      RECT 67.42 1.265 67.59 1.435 ;
      RECT 67.075 0.9 67.245 1.07 ;
      RECT 67.065 2.26 67.235 2.43 ;
      RECT 67.025 0.155 67.195 0.325 ;
      RECT 67.025 2.875 67.195 3.045 ;
      RECT 66.65 1.5 66.82 1.67 ;
      RECT 66.565 0.155 66.735 0.325 ;
      RECT 66.565 2.875 66.735 3.045 ;
      RECT 66.3 0.975 66.47 1.145 ;
      RECT 66.12 2.29 66.29 2.46 ;
      RECT 66.105 0.155 66.275 0.325 ;
      RECT 66.105 2.875 66.275 3.045 ;
      RECT 65.84 1.605 66.01 1.775 ;
      RECT 65.645 0.155 65.815 0.325 ;
      RECT 65.645 2.875 65.815 3.045 ;
      RECT 65.52 1.23 65.69 1.4 ;
      RECT 65.185 0.155 65.355 0.325 ;
      RECT 65.185 2.875 65.355 3.045 ;
      RECT 64.83 0.71 65 0.88 ;
      RECT 64.755 1.18 64.925 1.35 ;
      RECT 64.725 0.155 64.895 0.325 ;
      RECT 64.725 2.875 64.895 3.045 ;
      RECT 64.265 0.155 64.435 0.325 ;
      RECT 64.265 2.875 64.435 3.045 ;
      RECT 63.905 0.905 64.075 1.075 ;
      RECT 63.805 0.155 63.975 0.325 ;
      RECT 63.805 2.875 63.975 3.045 ;
      RECT 63.565 2.1 63.735 2.27 ;
      RECT 63.53 1.435 63.7 1.605 ;
      RECT 63.345 0.155 63.515 0.325 ;
      RECT 63.345 2.875 63.515 3.045 ;
      RECT 62.92 1.29 63.09 1.46 ;
      RECT 62.885 0.155 63.055 0.325 ;
      RECT 62.885 2.875 63.055 3.045 ;
      RECT 62.85 1.99 63.02 2.16 ;
      RECT 62.79 0.825 62.96 0.995 ;
      RECT 62.425 0.155 62.595 0.325 ;
      RECT 62.425 2.875 62.595 3.045 ;
      RECT 62.15 1.74 62.32 1.91 ;
      RECT 61.965 0.155 62.135 0.325 ;
      RECT 61.965 2.875 62.135 3.045 ;
      RECT 61.645 1.245 61.815 1.415 ;
      RECT 61.505 0.155 61.675 0.325 ;
      RECT 61.505 2.875 61.675 3.045 ;
      RECT 61.425 1.99 61.595 2.16 ;
      RECT 61.22 0.87 61.39 1.04 ;
      RECT 61.045 0.155 61.215 0.325 ;
      RECT 61.045 2.875 61.215 3.045 ;
      RECT 60.95 1.74 61.12 1.91 ;
      RECT 60.91 1.17 61.08 1.34 ;
      RECT 60.585 0.155 60.755 0.325 ;
      RECT 60.585 2.875 60.755 3.045 ;
      RECT 60.365 2.215 60.535 2.385 ;
      RECT 60.225 0.835 60.395 1.005 ;
      RECT 60.125 0.155 60.295 0.325 ;
      RECT 60.125 2.875 60.295 3.045 ;
      RECT 59.665 0.155 59.835 0.325 ;
      RECT 59.665 2.875 59.835 3.045 ;
      RECT 59.655 1.755 59.825 1.925 ;
      RECT 59.205 0.155 59.375 0.325 ;
      RECT 59.205 2.875 59.375 3.045 ;
      RECT 58.745 0.155 58.915 0.325 ;
      RECT 58.745 2.875 58.915 3.045 ;
      RECT 58.675 1.7 58.845 1.87 ;
      RECT 58.285 0.155 58.455 0.325 ;
      RECT 58.285 2.875 58.455 3.045 ;
      RECT 57.825 0.155 57.995 0.325 ;
      RECT 57.825 2.875 57.995 3.045 ;
      RECT 57.815 0.745 57.985 0.915 ;
      RECT 57.365 0.155 57.535 0.325 ;
      RECT 57.365 2.875 57.535 3.045 ;
      RECT 56.905 0.155 57.075 0.325 ;
      RECT 56.905 2.875 57.075 3.045 ;
      RECT 56.445 0.155 56.615 0.325 ;
      RECT 56.445 2.875 56.615 3.045 ;
      RECT 55.985 0.155 56.155 0.325 ;
      RECT 55.985 2.875 56.155 3.045 ;
      RECT 55.525 0.155 55.695 0.325 ;
      RECT 55.525 2.875 55.695 3.045 ;
      RECT 55.47 1.815 55.64 1.985 ;
      RECT 55.065 0.155 55.235 0.325 ;
      RECT 55.065 2.875 55.235 3.045 ;
      RECT 54.605 0.155 54.775 0.325 ;
      RECT 54.605 2.875 54.775 3.045 ;
      RECT 54.145 0.155 54.315 0.325 ;
      RECT 54.145 2.875 54.315 3.045 ;
      RECT 53.685 0.155 53.855 0.325 ;
      RECT 53.685 2.875 53.855 3.045 ;
      RECT 53.225 0.155 53.395 0.325 ;
      RECT 53.225 2.875 53.395 3.045 ;
      RECT 53.02 1.34 53.19 1.51 ;
      RECT 52.765 0.155 52.935 0.325 ;
      RECT 52.765 2.875 52.935 3.045 ;
      RECT 52.305 0.155 52.475 0.325 ;
      RECT 52.305 2.875 52.475 3.045 ;
      RECT 52.06 1.555 52.23 1.725 ;
      RECT 51.845 0.155 52.015 0.325 ;
      RECT 51.845 2.875 52.015 3.045 ;
      RECT 51.385 0.155 51.555 0.325 ;
      RECT 51.385 2.875 51.555 3.045 ;
      RECT 50.925 0.155 51.095 0.325 ;
      RECT 50.925 2.875 51.095 3.045 ;
      RECT 50.465 0.155 50.635 0.325 ;
      RECT 50.465 2.875 50.635 3.045 ;
      RECT 50.26 1.345 50.43 1.515 ;
      RECT 50.005 0.155 50.175 0.325 ;
      RECT 50.005 2.875 50.175 3.045 ;
      RECT 49.545 0.155 49.715 0.325 ;
      RECT 49.545 2.875 49.715 3.045 ;
      RECT 49.085 0.155 49.255 0.325 ;
      RECT 49.085 2.875 49.255 3.045 ;
      RECT 49.015 1.7 49.185 1.87 ;
      RECT 48.625 0.155 48.795 0.325 ;
      RECT 48.625 2.875 48.795 3.045 ;
      RECT 48.165 0.155 48.335 0.325 ;
      RECT 48.165 2.875 48.335 3.045 ;
      RECT 48.155 0.815 48.325 0.985 ;
      RECT 47.71 0.695 47.88 0.865 ;
      RECT 47.705 0.155 47.875 0.325 ;
      RECT 47.705 2.875 47.875 3.045 ;
      RECT 47.245 0.155 47.415 0.325 ;
      RECT 47.245 2.875 47.415 3.045 ;
      RECT 46.785 0.155 46.955 0.325 ;
      RECT 46.785 2.875 46.955 3.045 ;
      RECT 46.325 0.155 46.495 0.325 ;
      RECT 46.325 2.875 46.495 3.045 ;
      RECT 45.865 0.155 46.035 0.325 ;
      RECT 45.865 2.875 46.035 3.045 ;
      RECT 45.81 1.315 45.98 1.485 ;
      RECT 45.41 0.155 45.58 0.325 ;
      RECT 45.41 2.875 45.58 3.045 ;
      RECT 44.95 0.155 45.12 0.325 ;
      RECT 44.95 2.875 45.12 3.045 ;
      RECT 44.88 1.7 45.05 1.87 ;
      RECT 44.49 0.155 44.66 0.325 ;
      RECT 44.49 2.875 44.66 3.045 ;
      RECT 44.03 0.155 44.2 0.325 ;
      RECT 44.03 2.875 44.2 3.045 ;
      RECT 43.615 0.755 43.785 0.925 ;
      RECT 43.57 0.155 43.74 0.325 ;
      RECT 43.57 2.875 43.74 3.045 ;
      RECT 43.2 1.48 43.37 1.65 ;
      RECT 43.11 0.155 43.28 0.325 ;
      RECT 43.11 2.875 43.28 3.045 ;
      RECT 42.65 0.155 42.82 0.325 ;
      RECT 42.65 2.875 42.82 3.045 ;
      RECT 42.19 0.155 42.36 0.325 ;
      RECT 42.19 2.875 42.36 3.045 ;
      RECT 41.73 0.155 41.9 0.325 ;
      RECT 41.73 2.875 41.9 3.045 ;
      RECT 41.675 2.155 41.845 2.325 ;
      RECT 41.27 0.155 41.44 0.325 ;
      RECT 41.27 2.875 41.44 3.045 ;
      RECT 40.9 1.615 41.07 1.785 ;
      RECT 40.81 0.155 40.98 0.325 ;
      RECT 40.81 2.875 40.98 3.045 ;
      RECT 40.58 0.785 40.75 0.955 ;
      RECT 40.435 1.225 40.605 1.395 ;
      RECT 40.35 0.155 40.52 0.325 ;
      RECT 40.35 2.875 40.52 3.045 ;
      RECT 39.89 0.155 40.06 0.325 ;
      RECT 39.89 2.875 40.06 3.045 ;
      RECT 39.825 1.265 39.995 1.435 ;
      RECT 39.48 0.9 39.65 1.07 ;
      RECT 39.47 2.26 39.64 2.43 ;
      RECT 39.43 0.155 39.6 0.325 ;
      RECT 39.43 2.875 39.6 3.045 ;
      RECT 39.055 1.5 39.225 1.67 ;
      RECT 38.97 0.155 39.14 0.325 ;
      RECT 38.97 2.875 39.14 3.045 ;
      RECT 38.705 0.975 38.875 1.145 ;
      RECT 38.525 2.29 38.695 2.46 ;
      RECT 38.51 0.155 38.68 0.325 ;
      RECT 38.51 2.875 38.68 3.045 ;
      RECT 38.245 1.605 38.415 1.775 ;
      RECT 38.05 0.155 38.22 0.325 ;
      RECT 38.05 2.875 38.22 3.045 ;
      RECT 37.925 1.23 38.095 1.4 ;
      RECT 37.59 0.155 37.76 0.325 ;
      RECT 37.59 2.875 37.76 3.045 ;
      RECT 37.235 0.71 37.405 0.88 ;
      RECT 37.16 1.18 37.33 1.35 ;
      RECT 37.13 0.155 37.3 0.325 ;
      RECT 37.13 2.875 37.3 3.045 ;
      RECT 36.67 0.155 36.84 0.325 ;
      RECT 36.67 2.875 36.84 3.045 ;
      RECT 36.31 0.905 36.48 1.075 ;
      RECT 36.21 0.155 36.38 0.325 ;
      RECT 36.21 2.875 36.38 3.045 ;
      RECT 35.97 2.1 36.14 2.27 ;
      RECT 35.935 1.435 36.105 1.605 ;
      RECT 35.75 0.155 35.92 0.325 ;
      RECT 35.75 2.875 35.92 3.045 ;
      RECT 35.325 1.29 35.495 1.46 ;
      RECT 35.29 0.155 35.46 0.325 ;
      RECT 35.29 2.875 35.46 3.045 ;
      RECT 35.255 1.99 35.425 2.16 ;
      RECT 35.195 0.825 35.365 0.995 ;
      RECT 34.83 0.155 35 0.325 ;
      RECT 34.83 2.875 35 3.045 ;
      RECT 34.555 1.74 34.725 1.91 ;
      RECT 34.37 0.155 34.54 0.325 ;
      RECT 34.37 2.875 34.54 3.045 ;
      RECT 34.05 1.245 34.22 1.415 ;
      RECT 33.91 0.155 34.08 0.325 ;
      RECT 33.91 2.875 34.08 3.045 ;
      RECT 33.83 1.99 34 2.16 ;
      RECT 33.625 0.87 33.795 1.04 ;
      RECT 33.45 0.155 33.62 0.325 ;
      RECT 33.45 2.875 33.62 3.045 ;
      RECT 33.355 1.74 33.525 1.91 ;
      RECT 33.315 1.17 33.485 1.34 ;
      RECT 32.99 0.155 33.16 0.325 ;
      RECT 32.99 2.875 33.16 3.045 ;
      RECT 32.77 2.215 32.94 2.385 ;
      RECT 32.63 0.835 32.8 1.005 ;
      RECT 32.53 0.155 32.7 0.325 ;
      RECT 32.53 2.875 32.7 3.045 ;
      RECT 32.07 0.155 32.24 0.325 ;
      RECT 32.07 2.875 32.24 3.045 ;
      RECT 32.06 1.755 32.23 1.925 ;
      RECT 31.61 0.155 31.78 0.325 ;
      RECT 31.61 2.875 31.78 3.045 ;
      RECT 31.15 0.155 31.32 0.325 ;
      RECT 31.15 2.875 31.32 3.045 ;
      RECT 31.08 1.7 31.25 1.87 ;
      RECT 30.69 0.155 30.86 0.325 ;
      RECT 30.69 2.875 30.86 3.045 ;
      RECT 30.23 0.155 30.4 0.325 ;
      RECT 30.23 2.875 30.4 3.045 ;
      RECT 30.22 0.745 30.39 0.915 ;
      RECT 29.77 0.155 29.94 0.325 ;
      RECT 29.77 2.875 29.94 3.045 ;
      RECT 29.31 0.155 29.48 0.325 ;
      RECT 29.31 2.875 29.48 3.045 ;
      RECT 28.85 0.155 29.02 0.325 ;
      RECT 28.85 2.875 29.02 3.045 ;
      RECT 28.39 0.155 28.56 0.325 ;
      RECT 28.39 2.875 28.56 3.045 ;
      RECT 27.93 0.155 28.1 0.325 ;
      RECT 27.93 2.875 28.1 3.045 ;
      RECT 27.875 1.815 28.045 1.985 ;
      RECT 27.47 0.155 27.64 0.325 ;
      RECT 27.47 2.875 27.64 3.045 ;
      RECT 27.01 0.155 27.18 0.325 ;
      RECT 27.01 2.875 27.18 3.045 ;
      RECT 26.55 0.155 26.72 0.325 ;
      RECT 26.55 2.875 26.72 3.045 ;
      RECT 26.09 0.155 26.26 0.325 ;
      RECT 26.09 2.875 26.26 3.045 ;
      RECT 25.63 0.155 25.8 0.325 ;
      RECT 25.63 2.875 25.8 3.045 ;
      RECT 25.425 1.34 25.595 1.51 ;
      RECT 25.17 0.155 25.34 0.325 ;
      RECT 25.17 2.875 25.34 3.045 ;
      RECT 24.71 0.155 24.88 0.325 ;
      RECT 24.71 2.875 24.88 3.045 ;
      RECT 24.465 1.515 24.635 1.685 ;
      RECT 24.25 0.155 24.42 0.325 ;
      RECT 24.25 2.875 24.42 3.045 ;
      RECT 23.79 0.155 23.96 0.325 ;
      RECT 23.79 2.875 23.96 3.045 ;
      RECT 23.33 0.155 23.5 0.325 ;
      RECT 23.33 2.875 23.5 3.045 ;
      RECT 22.87 0.155 23.04 0.325 ;
      RECT 22.87 2.875 23.04 3.045 ;
      RECT 22.665 1.345 22.835 1.515 ;
      RECT 22.41 0.155 22.58 0.325 ;
      RECT 22.41 2.875 22.58 3.045 ;
      RECT 21.95 0.155 22.12 0.325 ;
      RECT 21.95 2.875 22.12 3.045 ;
      RECT 21.49 0.155 21.66 0.325 ;
      RECT 21.49 2.875 21.66 3.045 ;
      RECT 21.42 1.7 21.59 1.87 ;
      RECT 21.03 0.155 21.2 0.325 ;
      RECT 21.03 2.875 21.2 3.045 ;
      RECT 20.57 0.155 20.74 0.325 ;
      RECT 20.57 2.875 20.74 3.045 ;
      RECT 20.56 0.815 20.73 0.985 ;
      RECT 20.115 0.695 20.285 0.865 ;
      RECT 20.11 0.155 20.28 0.325 ;
      RECT 20.11 2.875 20.28 3.045 ;
      RECT 19.65 0.155 19.82 0.325 ;
      RECT 19.65 2.875 19.82 3.045 ;
      RECT 19.19 0.155 19.36 0.325 ;
      RECT 19.19 2.875 19.36 3.045 ;
      RECT 18.73 0.155 18.9 0.325 ;
      RECT 18.73 2.875 18.9 3.045 ;
      RECT 18.27 0.155 18.44 0.325 ;
      RECT 18.27 2.875 18.44 3.045 ;
      RECT 18.215 1.315 18.385 1.485 ;
      RECT 17.815 0.155 17.985 0.325 ;
      RECT 17.815 2.875 17.985 3.045 ;
      RECT 17.355 0.155 17.525 0.325 ;
      RECT 17.355 2.875 17.525 3.045 ;
      RECT 17.285 1.7 17.455 1.87 ;
      RECT 16.895 0.155 17.065 0.325 ;
      RECT 16.895 2.875 17.065 3.045 ;
      RECT 16.435 0.155 16.605 0.325 ;
      RECT 16.435 2.875 16.605 3.045 ;
      RECT 16.02 0.755 16.19 0.925 ;
      RECT 15.975 0.155 16.145 0.325 ;
      RECT 15.975 2.875 16.145 3.045 ;
      RECT 15.605 1.48 15.775 1.65 ;
      RECT 15.515 0.155 15.685 0.325 ;
      RECT 15.515 2.875 15.685 3.045 ;
      RECT 15.055 0.155 15.225 0.325 ;
      RECT 15.055 2.875 15.225 3.045 ;
      RECT 14.595 0.155 14.765 0.325 ;
      RECT 14.595 2.875 14.765 3.045 ;
      RECT 14.135 0.155 14.305 0.325 ;
      RECT 14.135 2.875 14.305 3.045 ;
      RECT 14.08 2.155 14.25 2.325 ;
      RECT 13.675 0.155 13.845 0.325 ;
      RECT 13.675 2.875 13.845 3.045 ;
      RECT 13.305 1.615 13.475 1.785 ;
      RECT 13.215 0.155 13.385 0.325 ;
      RECT 13.215 2.875 13.385 3.045 ;
      RECT 12.985 0.785 13.155 0.955 ;
      RECT 12.84 1.225 13.01 1.395 ;
      RECT 12.755 0.155 12.925 0.325 ;
      RECT 12.755 2.875 12.925 3.045 ;
      RECT 12.295 0.155 12.465 0.325 ;
      RECT 12.295 2.875 12.465 3.045 ;
      RECT 12.23 1.265 12.4 1.435 ;
      RECT 11.885 0.9 12.055 1.07 ;
      RECT 11.875 2.26 12.045 2.43 ;
      RECT 11.835 0.155 12.005 0.325 ;
      RECT 11.835 2.875 12.005 3.045 ;
      RECT 11.46 1.5 11.63 1.67 ;
      RECT 11.375 0.155 11.545 0.325 ;
      RECT 11.375 2.875 11.545 3.045 ;
      RECT 11.11 0.975 11.28 1.145 ;
      RECT 10.93 2.29 11.1 2.46 ;
      RECT 10.915 0.155 11.085 0.325 ;
      RECT 10.915 2.875 11.085 3.045 ;
      RECT 10.65 1.605 10.82 1.775 ;
      RECT 10.455 0.155 10.625 0.325 ;
      RECT 10.455 2.875 10.625 3.045 ;
      RECT 10.33 1.23 10.5 1.4 ;
      RECT 9.995 0.155 10.165 0.325 ;
      RECT 9.995 2.875 10.165 3.045 ;
      RECT 9.64 0.71 9.81 0.88 ;
      RECT 9.565 1.18 9.735 1.35 ;
      RECT 9.535 0.155 9.705 0.325 ;
      RECT 9.535 2.875 9.705 3.045 ;
      RECT 9.075 0.155 9.245 0.325 ;
      RECT 9.075 2.875 9.245 3.045 ;
      RECT 8.715 0.905 8.885 1.075 ;
      RECT 8.615 0.155 8.785 0.325 ;
      RECT 8.615 2.875 8.785 3.045 ;
      RECT 8.375 2.1 8.545 2.27 ;
      RECT 8.34 1.435 8.51 1.605 ;
      RECT 8.155 0.155 8.325 0.325 ;
      RECT 8.155 2.875 8.325 3.045 ;
      RECT 7.73 1.29 7.9 1.46 ;
      RECT 7.695 0.155 7.865 0.325 ;
      RECT 7.695 2.875 7.865 3.045 ;
      RECT 7.66 1.99 7.83 2.16 ;
      RECT 7.6 0.825 7.77 0.995 ;
      RECT 7.235 0.155 7.405 0.325 ;
      RECT 7.235 2.875 7.405 3.045 ;
      RECT 6.96 1.74 7.13 1.91 ;
      RECT 6.775 0.155 6.945 0.325 ;
      RECT 6.775 2.875 6.945 3.045 ;
      RECT 6.455 1.245 6.625 1.415 ;
      RECT 6.315 0.155 6.485 0.325 ;
      RECT 6.315 2.875 6.485 3.045 ;
      RECT 6.235 1.99 6.405 2.16 ;
      RECT 6.03 0.87 6.2 1.04 ;
      RECT 5.855 0.155 6.025 0.325 ;
      RECT 5.855 2.875 6.025 3.045 ;
      RECT 5.76 1.74 5.93 1.91 ;
      RECT 5.72 1.17 5.89 1.34 ;
      RECT 5.395 0.155 5.565 0.325 ;
      RECT 5.395 2.875 5.565 3.045 ;
      RECT 5.175 2.215 5.345 2.385 ;
      RECT 5.035 0.835 5.205 1.005 ;
      RECT 4.935 0.155 5.105 0.325 ;
      RECT 4.935 2.875 5.105 3.045 ;
      RECT 4.475 0.155 4.645 0.325 ;
      RECT 4.475 2.875 4.645 3.045 ;
      RECT 4.465 1.755 4.635 1.925 ;
      RECT 4.015 0.155 4.185 0.325 ;
      RECT 4.015 2.875 4.185 3.045 ;
      RECT 3.555 0.155 3.725 0.325 ;
      RECT 3.555 2.875 3.725 3.045 ;
      RECT 3.485 1.7 3.655 1.87 ;
      RECT 3.095 0.155 3.265 0.325 ;
      RECT 3.095 2.875 3.265 3.045 ;
      RECT 2.635 0.155 2.805 0.325 ;
      RECT 2.635 2.875 2.805 3.045 ;
      RECT 2.625 0.745 2.795 0.915 ;
      RECT 2.175 0.155 2.345 0.325 ;
      RECT 2.175 2.875 2.345 3.045 ;
      RECT 1.715 0.155 1.885 0.325 ;
      RECT 1.715 2.875 1.885 3.045 ;
      RECT 1.255 0.155 1.425 0.325 ;
      RECT 1.255 2.875 1.425 3.045 ;
      RECT 0.795 0.155 0.965 0.325 ;
      RECT 0.795 2.875 0.965 3.045 ;
      RECT 0.335 0.155 0.505 0.325 ;
      RECT 0.335 2.875 0.505 3.045 ;
      RECT 0.28 1.815 0.45 1.985 ;
      RECT -0.125 0.155 0.045 0.325 ;
      RECT -0.125 2.875 0.045 3.045 ;
      RECT -0.585 0.155 -0.415 0.325 ;
      RECT -0.585 2.875 -0.415 3.045 ;
      RECT -1.045 0.155 -0.875 0.325 ;
      RECT -1.045 2.875 -0.875 3.045 ;
      RECT -1.495 1.7 -1.325 1.87 ;
      RECT -1.505 0.155 -1.335 0.325 ;
      RECT -1.505 2.875 -1.335 3.045 ;
      RECT -1.925 0.695 -1.755 0.865 ;
      RECT -1.965 0.155 -1.795 0.325 ;
      RECT -1.965 2.875 -1.795 3.045 ;
      RECT -2.425 0.155 -2.255 0.325 ;
      RECT -2.425 2.875 -2.255 3.045 ;
      RECT -2.885 0.155 -2.715 0.325 ;
      RECT -2.885 2.875 -2.715 3.045 ;
      RECT -3.345 0.155 -3.175 0.325 ;
      RECT -3.345 2.875 -3.175 3.045 ;
      RECT -3.775 1.815 -3.605 1.985 ;
      RECT -3.805 0.155 -3.635 0.325 ;
      RECT -3.805 2.875 -3.635 3.045 ;
    LAYER li ;
      RECT 112.56 0.155 112.835 1.655 ;
      RECT 84.965 0.155 85.24 1.655 ;
      RECT 57.37 0.155 57.645 1.655 ;
      RECT 29.775 0.155 30.05 1.655 ;
      RECT 2.18 0.155 2.455 1.655 ;
      RECT 137.105 0.155 137.335 1.145 ;
      RECT 135.725 0.155 135.955 1.145 ;
      RECT 134.345 0.155 134.575 1.145 ;
      RECT 132.965 0.155 133.195 1.145 ;
      RECT 109.51 0.155 109.74 1.145 ;
      RECT 108.13 0.155 108.36 1.145 ;
      RECT 106.75 0.155 106.98 1.145 ;
      RECT 105.37 0.155 105.6 1.145 ;
      RECT 81.915 0.155 82.145 1.145 ;
      RECT 80.535 0.155 80.765 1.145 ;
      RECT 79.155 0.155 79.385 1.145 ;
      RECT 77.775 0.155 78.005 1.145 ;
      RECT 54.32 0.155 54.55 1.145 ;
      RECT 52.94 0.155 53.17 1.145 ;
      RECT 51.56 0.155 51.79 1.145 ;
      RECT 50.18 0.155 50.41 1.145 ;
      RECT 26.725 0.155 26.955 1.145 ;
      RECT 25.345 0.155 25.575 1.145 ;
      RECT 23.965 0.155 24.195 1.145 ;
      RECT 22.585 0.155 22.815 1.145 ;
      RECT 131.31 0.155 131.82 0.86 ;
      RECT 127.175 0.155 127.685 0.86 ;
      RECT 113.375 0.155 113.885 0.86 ;
      RECT 103.715 0.155 104.225 0.86 ;
      RECT 99.58 0.155 100.09 0.86 ;
      RECT 85.78 0.155 86.29 0.86 ;
      RECT 76.12 0.155 76.63 0.86 ;
      RECT 71.985 0.155 72.495 0.86 ;
      RECT 58.185 0.155 58.695 0.86 ;
      RECT 48.525 0.155 49.035 0.86 ;
      RECT 44.39 0.155 44.9 0.86 ;
      RECT 30.59 0.155 31.1 0.86 ;
      RECT 20.93 0.155 21.44 0.86 ;
      RECT 16.795 0.155 17.305 0.86 ;
      RECT 2.995 0.155 3.505 0.86 ;
      RECT -1.145 0.155 -0.635 0.86 ;
      RECT 122.84 0.155 123.01 0.825 ;
      RECT 120.88 0.155 121.05 0.825 ;
      RECT 118.44 0.155 118.61 0.825 ;
      RECT 117.48 0.155 117.65 0.825 ;
      RECT 116.96 0.155 117.13 0.825 ;
      RECT 116 0.155 116.17 0.825 ;
      RECT 115.04 0.155 115.21 0.825 ;
      RECT 95.245 0.155 95.415 0.825 ;
      RECT 93.285 0.155 93.455 0.825 ;
      RECT 90.845 0.155 91.015 0.825 ;
      RECT 89.885 0.155 90.055 0.825 ;
      RECT 89.365 0.155 89.535 0.825 ;
      RECT 88.405 0.155 88.575 0.825 ;
      RECT 87.445 0.155 87.615 0.825 ;
      RECT 67.65 0.155 67.82 0.825 ;
      RECT 65.69 0.155 65.86 0.825 ;
      RECT 63.25 0.155 63.42 0.825 ;
      RECT 62.29 0.155 62.46 0.825 ;
      RECT 61.77 0.155 61.94 0.825 ;
      RECT 60.81 0.155 60.98 0.825 ;
      RECT 59.85 0.155 60.02 0.825 ;
      RECT 40.055 0.155 40.225 0.825 ;
      RECT 38.095 0.155 38.265 0.825 ;
      RECT 35.655 0.155 35.825 0.825 ;
      RECT 34.695 0.155 34.865 0.825 ;
      RECT 34.175 0.155 34.345 0.825 ;
      RECT 33.215 0.155 33.385 0.825 ;
      RECT 32.255 0.155 32.425 0.825 ;
      RECT 12.46 0.155 12.63 0.825 ;
      RECT 10.5 0.155 10.67 0.825 ;
      RECT 8.06 0.155 8.23 0.825 ;
      RECT 7.1 0.155 7.27 0.825 ;
      RECT 6.58 0.155 6.75 0.825 ;
      RECT 5.62 0.155 5.79 0.825 ;
      RECT 4.66 0.155 4.83 0.825 ;
      RECT 129.02 0.155 129.35 0.725 ;
      RECT 124.885 0.155 125.215 0.725 ;
      RECT 111.085 0.155 111.415 0.725 ;
      RECT 101.425 0.155 101.755 0.725 ;
      RECT 97.29 0.155 97.62 0.725 ;
      RECT 83.49 0.155 83.82 0.725 ;
      RECT 73.83 0.155 74.16 0.725 ;
      RECT 69.695 0.155 70.025 0.725 ;
      RECT 55.895 0.155 56.225 0.725 ;
      RECT 46.235 0.155 46.565 0.725 ;
      RECT 42.1 0.155 42.43 0.725 ;
      RECT 28.3 0.155 28.63 0.725 ;
      RECT 18.64 0.155 18.97 0.725 ;
      RECT 14.505 0.155 14.835 0.725 ;
      RECT 0.705 0.155 1.035 0.725 ;
      RECT -3.435 0.155 -3.105 0.725 ;
      RECT -3.95 0.155 138.165 0.325 ;
      RECT -3.95 2.875 138.165 3.045 ;
      RECT 137.125 1.735 137.335 3.045 ;
      RECT 135.745 1.735 135.955 3.045 ;
      RECT 134.365 1.735 134.575 3.045 ;
      RECT 132.985 1.735 133.195 3.045 ;
      RECT 131.64 2.115 131.81 3.045 ;
      RECT 129.1 1.735 129.27 3.045 ;
      RECT 127.505 2.115 127.675 3.045 ;
      RECT 124.965 1.735 125.135 3.045 ;
      RECT 123.8 2.285 123.97 3.045 ;
      RECT 122.84 2.375 123.01 3.045 ;
      RECT 120.4 2.375 120.57 3.045 ;
      RECT 119.4 2.375 119.57 3.045 ;
      RECT 118.44 2.375 118.61 3.045 ;
      RECT 116 2.375 116.17 3.045 ;
      RECT 113.705 2.115 113.875 3.045 ;
      RECT 111.165 1.735 111.335 3.045 ;
      RECT 109.53 1.735 109.74 3.045 ;
      RECT 108.15 1.735 108.36 3.045 ;
      RECT 106.77 1.735 106.98 3.045 ;
      RECT 105.39 1.735 105.6 3.045 ;
      RECT 104.045 2.115 104.215 3.045 ;
      RECT 101.505 1.735 101.675 3.045 ;
      RECT 99.91 2.115 100.08 3.045 ;
      RECT 97.37 1.735 97.54 3.045 ;
      RECT 96.205 2.285 96.375 3.045 ;
      RECT 95.245 2.375 95.415 3.045 ;
      RECT 92.805 2.375 92.975 3.045 ;
      RECT 91.805 2.375 91.975 3.045 ;
      RECT 90.845 2.375 91.015 3.045 ;
      RECT 88.405 2.375 88.575 3.045 ;
      RECT 86.11 2.115 86.28 3.045 ;
      RECT 83.57 1.735 83.74 3.045 ;
      RECT 81.935 1.735 82.145 3.045 ;
      RECT 80.555 1.735 80.765 3.045 ;
      RECT 79.175 1.735 79.385 3.045 ;
      RECT 77.795 1.735 78.005 3.045 ;
      RECT 76.45 2.115 76.62 3.045 ;
      RECT 73.91 1.735 74.08 3.045 ;
      RECT 72.315 2.115 72.485 3.045 ;
      RECT 69.775 1.735 69.945 3.045 ;
      RECT 68.61 2.285 68.78 3.045 ;
      RECT 67.65 2.375 67.82 3.045 ;
      RECT 65.21 2.375 65.38 3.045 ;
      RECT 64.21 2.375 64.38 3.045 ;
      RECT 63.25 2.375 63.42 3.045 ;
      RECT 60.81 2.375 60.98 3.045 ;
      RECT 58.515 2.115 58.685 3.045 ;
      RECT 55.975 1.735 56.145 3.045 ;
      RECT 54.34 1.735 54.55 3.045 ;
      RECT 52.96 1.735 53.17 3.045 ;
      RECT 51.58 1.735 51.79 3.045 ;
      RECT 50.2 1.735 50.41 3.045 ;
      RECT 48.855 2.115 49.025 3.045 ;
      RECT 46.315 1.735 46.485 3.045 ;
      RECT 44.72 2.115 44.89 3.045 ;
      RECT 42.18 1.735 42.35 3.045 ;
      RECT 41.015 2.285 41.185 3.045 ;
      RECT 40.055 2.375 40.225 3.045 ;
      RECT 37.615 2.375 37.785 3.045 ;
      RECT 36.615 2.375 36.785 3.045 ;
      RECT 35.655 2.375 35.825 3.045 ;
      RECT 33.215 2.375 33.385 3.045 ;
      RECT 30.92 2.115 31.09 3.045 ;
      RECT 28.38 1.735 28.55 3.045 ;
      RECT 26.745 1.735 26.955 3.045 ;
      RECT 25.365 1.735 25.575 3.045 ;
      RECT 23.985 1.735 24.195 3.045 ;
      RECT 22.605 1.735 22.815 3.045 ;
      RECT 21.26 2.115 21.43 3.045 ;
      RECT 18.72 1.735 18.89 3.045 ;
      RECT 17.125 2.115 17.295 3.045 ;
      RECT 14.585 1.735 14.755 3.045 ;
      RECT 13.42 2.285 13.59 3.045 ;
      RECT 12.46 2.375 12.63 3.045 ;
      RECT 10.02 2.375 10.19 3.045 ;
      RECT 9.02 2.375 9.19 3.045 ;
      RECT 8.06 2.375 8.23 3.045 ;
      RECT 5.62 2.375 5.79 3.045 ;
      RECT 3.325 2.115 3.495 3.045 ;
      RECT 0.785 1.735 0.955 3.045 ;
      RECT -0.815 2.115 -0.645 3.045 ;
      RECT -3.355 1.735 -3.185 3.045 ;
      RECT 137.505 1.725 137.835 2.705 ;
      RECT 137.605 0.495 137.835 2.705 ;
      RECT 137.505 0.495 137.835 1.125 ;
      RECT 136.125 1.725 136.455 2.705 ;
      RECT 136.225 0.495 136.455 2.705 ;
      RECT 136.225 1.315 137.435 1.555 ;
      RECT 136.125 0.495 136.455 1.125 ;
      RECT 134.745 1.725 135.075 2.705 ;
      RECT 134.845 0.495 135.075 2.705 ;
      RECT 134.745 0.495 135.075 1.125 ;
      RECT 133.365 1.725 133.695 2.705 ;
      RECT 133.465 0.495 133.695 2.705 ;
      RECT 133.465 1.315 134.675 1.555 ;
      RECT 133.365 0.495 133.695 1.125 ;
      RECT 132.045 2.115 132.56 2.525 ;
      RECT 132.22 1.135 132.56 2.525 ;
      RECT 131.33 1.135 132.56 1.305 ;
      RECT 132.04 0.53 132.285 1.305 ;
      RECT 129.44 2.535 131.47 2.705 ;
      RECT 131.3 1.68 131.47 2.705 ;
      RECT 129.44 1.235 129.61 2.705 ;
      RECT 131.3 1.68 132.05 1.87 ;
      RECT 129.415 1.235 129.61 1.565 ;
      RECT 130.12 1.855 131.13 2.025 ;
      RECT 130.94 0.495 131.13 2.025 ;
      RECT 130.12 1.055 130.29 2.025 ;
      RECT 129.78 2.195 130.905 2.365 ;
      RECT 129.78 0.495 129.95 2.365 ;
      RECT 128.935 1.235 129.19 1.565 ;
      RECT 129.02 0.895 129.19 1.565 ;
      RECT 129.02 0.895 129.95 1.065 ;
      RECT 129.775 0.495 129.95 1.065 ;
      RECT 129.775 0.495 130.305 0.86 ;
      RECT 128.595 1.735 128.93 2.705 ;
      RECT 128.595 0.495 128.765 2.705 ;
      RECT 128.595 0.495 128.85 1.065 ;
      RECT 127.91 2.115 128.425 2.525 ;
      RECT 128.085 1.135 128.425 2.525 ;
      RECT 127.195 1.135 128.425 1.305 ;
      RECT 127.905 0.53 128.15 1.305 ;
      RECT 125.305 2.535 127.335 2.705 ;
      RECT 127.165 1.68 127.335 2.705 ;
      RECT 125.305 1.235 125.475 2.705 ;
      RECT 127.165 1.68 127.915 1.87 ;
      RECT 125.28 1.235 125.475 1.565 ;
      RECT 125.985 1.855 126.995 2.025 ;
      RECT 126.805 0.495 126.995 2.025 ;
      RECT 125.985 1.055 126.155 2.025 ;
      RECT 125.645 2.195 126.77 2.365 ;
      RECT 125.645 0.495 125.815 2.365 ;
      RECT 124.8 1.235 125.055 1.565 ;
      RECT 124.885 0.895 125.055 1.565 ;
      RECT 124.885 0.895 125.815 1.065 ;
      RECT 125.64 0.495 125.815 1.065 ;
      RECT 125.64 0.495 126.17 0.86 ;
      RECT 124.46 1.735 124.795 2.705 ;
      RECT 124.46 0.495 124.63 2.705 ;
      RECT 124.46 0.495 124.715 1.065 ;
      RECT 123.365 0.715 124.095 0.955 ;
      RECT 123.907 0.51 124.095 0.955 ;
      RECT 123.735 0.522 124.11 0.949 ;
      RECT 123.65 0.537 124.13 0.934 ;
      RECT 123.65 0.552 124.135 0.924 ;
      RECT 123.605 0.572 124.15 0.916 ;
      RECT 123.582 0.607 124.165 0.87 ;
      RECT 123.496 0.63 124.17 0.83 ;
      RECT 123.496 0.648 124.18 0.8 ;
      RECT 123.365 0.717 124.185 0.763 ;
      RECT 123.41 0.66 124.18 0.8 ;
      RECT 123.496 0.612 124.165 0.87 ;
      RECT 123.582 0.581 124.15 0.916 ;
      RECT 123.605 0.562 124.135 0.924 ;
      RECT 123.65 0.535 124.11 0.949 ;
      RECT 123.735 0.517 124.095 0.955 ;
      RECT 123.821 0.511 124.095 0.955 ;
      RECT 123.907 0.506 124.04 0.955 ;
      RECT 123.993 0.501 124.04 0.955 ;
      RECT 123.685 1.399 123.855 1.785 ;
      RECT 123.68 1.399 123.855 1.78 ;
      RECT 123.655 1.399 123.855 1.745 ;
      RECT 123.655 1.427 123.865 1.735 ;
      RECT 123.635 1.427 123.865 1.695 ;
      RECT 123.63 1.427 123.865 1.668 ;
      RECT 123.63 1.445 123.87 1.66 ;
      RECT 123.575 1.445 123.87 1.595 ;
      RECT 123.575 1.462 123.88 1.578 ;
      RECT 123.565 1.462 123.88 1.518 ;
      RECT 123.565 1.479 123.885 1.515 ;
      RECT 123.56 1.315 123.73 1.493 ;
      RECT 123.56 1.349 123.816 1.493 ;
      RECT 123.555 2.115 123.56 2.128 ;
      RECT 123.55 2.01 123.555 2.133 ;
      RECT 123.525 1.87 123.55 2.148 ;
      RECT 123.49 1.821 123.525 2.18 ;
      RECT 123.485 1.789 123.49 2.2 ;
      RECT 123.48 1.78 123.485 2.2 ;
      RECT 123.4 1.745 123.48 2.2 ;
      RECT 123.337 1.715 123.4 2.2 ;
      RECT 123.251 1.703 123.337 2.2 ;
      RECT 123.165 1.689 123.251 2.2 ;
      RECT 123.085 1.676 123.165 2.186 ;
      RECT 123.05 1.668 123.085 2.166 ;
      RECT 123.04 1.665 123.05 2.157 ;
      RECT 123.01 1.66 123.04 2.144 ;
      RECT 122.96 1.635 123.01 2.12 ;
      RECT 122.946 1.609 122.96 2.102 ;
      RECT 122.86 1.569 122.946 2.078 ;
      RECT 122.815 1.517 122.86 2.047 ;
      RECT 122.805 1.492 122.815 2.034 ;
      RECT 122.8 1.273 122.805 1.295 ;
      RECT 122.795 1.475 122.805 2.03 ;
      RECT 122.795 1.271 122.8 1.385 ;
      RECT 122.785 1.267 122.795 2.026 ;
      RECT 122.741 1.265 122.785 2.014 ;
      RECT 122.655 1.265 122.741 1.985 ;
      RECT 122.625 1.265 122.655 1.958 ;
      RECT 122.61 1.265 122.625 1.946 ;
      RECT 122.57 1.277 122.61 1.931 ;
      RECT 122.55 1.296 122.57 1.91 ;
      RECT 122.54 1.306 122.55 1.894 ;
      RECT 122.53 1.312 122.54 1.883 ;
      RECT 122.51 1.322 122.53 1.866 ;
      RECT 122.505 1.331 122.51 1.853 ;
      RECT 122.5 1.335 122.505 1.803 ;
      RECT 122.49 1.341 122.5 1.72 ;
      RECT 122.485 1.345 122.49 1.634 ;
      RECT 122.48 1.365 122.485 1.571 ;
      RECT 122.475 1.388 122.48 1.518 ;
      RECT 122.47 1.406 122.475 1.463 ;
      RECT 123.08 1.225 123.25 1.485 ;
      RECT 123.25 1.19 123.295 1.471 ;
      RECT 123.211 1.192 123.3 1.454 ;
      RECT 123.1 1.209 123.386 1.425 ;
      RECT 123.1 1.224 123.39 1.397 ;
      RECT 123.1 1.205 123.3 1.454 ;
      RECT 123.125 1.193 123.25 1.485 ;
      RECT 123.211 1.191 123.295 1.471 ;
      RECT 122.265 0.58 122.435 1.07 ;
      RECT 122.265 0.58 122.47 1.05 ;
      RECT 122.4 0.5 122.51 1.01 ;
      RECT 122.381 0.504 122.53 0.98 ;
      RECT 122.295 0.512 122.55 0.963 ;
      RECT 122.295 0.518 122.555 0.953 ;
      RECT 122.295 0.527 122.575 0.941 ;
      RECT 122.27 0.552 122.605 0.919 ;
      RECT 122.27 0.572 122.61 0.899 ;
      RECT 122.265 0.585 122.62 0.879 ;
      RECT 122.265 0.652 122.625 0.86 ;
      RECT 122.265 0.785 122.63 0.847 ;
      RECT 122.26 0.59 122.62 0.68 ;
      RECT 122.27 0.547 122.575 0.941 ;
      RECT 122.381 0.502 122.51 1.01 ;
      RECT 122.255 2.255 122.555 2.51 ;
      RECT 122.34 2.221 122.555 2.51 ;
      RECT 122.34 2.224 122.56 2.37 ;
      RECT 122.275 2.245 122.56 2.37 ;
      RECT 122.31 2.235 122.555 2.51 ;
      RECT 122.305 2.24 122.56 2.37 ;
      RECT 122.34 2.219 122.541 2.51 ;
      RECT 122.426 2.21 122.541 2.51 ;
      RECT 122.426 2.204 122.455 2.51 ;
      RECT 121.915 1.845 121.925 2.335 ;
      RECT 121.575 1.78 121.585 2.08 ;
      RECT 122.09 1.952 122.095 2.171 ;
      RECT 122.08 1.932 122.09 2.188 ;
      RECT 122.07 1.912 122.08 2.218 ;
      RECT 122.065 1.902 122.07 2.233 ;
      RECT 122.06 1.898 122.065 2.238 ;
      RECT 122.045 1.89 122.06 2.245 ;
      RECT 122.005 1.87 122.045 2.27 ;
      RECT 121.98 1.852 122.005 2.303 ;
      RECT 121.975 1.85 121.98 2.316 ;
      RECT 121.955 1.847 121.975 2.32 ;
      RECT 121.925 1.845 121.955 2.33 ;
      RECT 121.855 1.847 121.915 2.331 ;
      RECT 121.835 1.847 121.855 2.325 ;
      RECT 121.81 1.845 121.835 2.322 ;
      RECT 121.775 1.84 121.81 2.318 ;
      RECT 121.755 1.834 121.775 2.305 ;
      RECT 121.745 1.831 121.755 2.293 ;
      RECT 121.725 1.828 121.745 2.278 ;
      RECT 121.705 1.824 121.725 2.26 ;
      RECT 121.7 1.821 121.705 2.25 ;
      RECT 121.695 1.82 121.7 2.248 ;
      RECT 121.685 1.817 121.695 2.24 ;
      RECT 121.675 1.811 121.685 2.223 ;
      RECT 121.665 1.805 121.675 2.205 ;
      RECT 121.655 1.799 121.665 2.193 ;
      RECT 121.645 1.793 121.655 2.173 ;
      RECT 121.64 1.789 121.645 2.158 ;
      RECT 121.635 1.787 121.64 2.15 ;
      RECT 121.63 1.785 121.635 2.143 ;
      RECT 121.625 1.783 121.63 2.133 ;
      RECT 121.62 1.781 121.625 2.127 ;
      RECT 121.61 1.78 121.62 2.117 ;
      RECT 121.6 1.78 121.61 2.108 ;
      RECT 121.585 1.78 121.6 2.093 ;
      RECT 121.545 1.78 121.575 2.077 ;
      RECT 121.525 1.782 121.545 2.072 ;
      RECT 121.52 1.787 121.525 2.07 ;
      RECT 121.49 1.795 121.52 2.068 ;
      RECT 121.46 1.81 121.49 2.067 ;
      RECT 121.415 1.832 121.46 2.072 ;
      RECT 121.41 1.847 121.415 2.076 ;
      RECT 121.395 1.852 121.41 2.078 ;
      RECT 121.39 1.856 121.395 2.08 ;
      RECT 121.33 1.879 121.39 2.089 ;
      RECT 121.31 1.905 121.33 2.102 ;
      RECT 121.3 1.912 121.31 2.106 ;
      RECT 121.285 1.919 121.3 2.109 ;
      RECT 121.265 1.929 121.285 2.112 ;
      RECT 121.26 1.937 121.265 2.115 ;
      RECT 121.215 1.942 121.26 2.122 ;
      RECT 121.205 1.945 121.215 2.129 ;
      RECT 121.195 1.945 121.205 2.133 ;
      RECT 121.16 1.947 121.195 2.145 ;
      RECT 121.14 1.95 121.16 2.158 ;
      RECT 121.1 1.953 121.14 2.169 ;
      RECT 121.085 1.955 121.1 2.182 ;
      RECT 121.075 1.955 121.085 2.187 ;
      RECT 121.05 1.956 121.075 2.195 ;
      RECT 121.04 1.958 121.05 2.2 ;
      RECT 121.035 1.959 121.04 2.203 ;
      RECT 121.01 1.957 121.035 2.206 ;
      RECT 120.995 1.955 121.01 2.207 ;
      RECT 120.975 1.952 120.995 2.209 ;
      RECT 120.955 1.947 120.975 2.209 ;
      RECT 120.895 1.942 120.955 2.206 ;
      RECT 120.86 1.917 120.895 2.202 ;
      RECT 120.85 1.894 120.86 2.2 ;
      RECT 120.82 1.871 120.85 2.2 ;
      RECT 120.81 1.85 120.82 2.2 ;
      RECT 120.785 1.832 120.81 2.198 ;
      RECT 120.77 1.81 120.785 2.195 ;
      RECT 120.755 1.792 120.77 2.193 ;
      RECT 120.735 1.782 120.755 2.191 ;
      RECT 120.72 1.777 120.735 2.19 ;
      RECT 120.705 1.775 120.72 2.189 ;
      RECT 120.675 1.776 120.705 2.187 ;
      RECT 120.655 1.779 120.675 2.185 ;
      RECT 120.598 1.783 120.655 2.185 ;
      RECT 120.512 1.792 120.598 2.185 ;
      RECT 120.426 1.803 120.512 2.185 ;
      RECT 120.34 1.814 120.426 2.185 ;
      RECT 120.32 1.821 120.34 2.193 ;
      RECT 120.31 1.824 120.32 2.2 ;
      RECT 120.245 1.829 120.31 2.218 ;
      RECT 120.215 1.836 120.245 2.243 ;
      RECT 120.205 1.839 120.215 2.25 ;
      RECT 120.16 1.843 120.205 2.255 ;
      RECT 120.13 1.848 120.16 2.26 ;
      RECT 120.129 1.85 120.13 2.26 ;
      RECT 120.043 1.856 120.129 2.26 ;
      RECT 119.957 1.867 120.043 2.26 ;
      RECT 119.871 1.879 119.957 2.26 ;
      RECT 119.785 1.89 119.871 2.26 ;
      RECT 119.77 1.897 119.785 2.255 ;
      RECT 119.765 1.899 119.77 2.249 ;
      RECT 119.745 1.91 119.765 2.244 ;
      RECT 119.735 1.928 119.745 2.238 ;
      RECT 119.73 1.94 119.735 2.038 ;
      RECT 122.025 0.693 122.045 0.78 ;
      RECT 122.02 0.628 122.025 0.812 ;
      RECT 122.01 0.595 122.02 0.817 ;
      RECT 122.005 0.575 122.01 0.823 ;
      RECT 121.975 0.575 122.005 0.84 ;
      RECT 121.926 0.575 121.975 0.876 ;
      RECT 121.84 0.575 121.926 0.934 ;
      RECT 121.811 0.585 121.84 0.983 ;
      RECT 121.725 0.627 121.811 1.036 ;
      RECT 121.705 0.665 121.725 1.083 ;
      RECT 121.68 0.682 121.705 1.103 ;
      RECT 121.67 0.696 121.68 1.123 ;
      RECT 121.665 0.702 121.67 1.133 ;
      RECT 121.66 0.706 121.665 1.14 ;
      RECT 121.61 0.726 121.66 1.145 ;
      RECT 121.545 0.77 121.61 1.145 ;
      RECT 121.52 0.82 121.545 1.145 ;
      RECT 121.51 0.85 121.52 1.145 ;
      RECT 121.505 0.877 121.51 1.145 ;
      RECT 121.5 0.895 121.505 1.145 ;
      RECT 121.49 0.937 121.5 1.145 ;
      RECT 121.84 1.495 122.01 1.67 ;
      RECT 121.78 1.323 121.84 1.658 ;
      RECT 121.77 1.316 121.78 1.641 ;
      RECT 121.725 1.495 122.01 1.621 ;
      RECT 121.706 1.495 122.01 1.599 ;
      RECT 121.62 1.495 122.01 1.564 ;
      RECT 121.6 1.315 121.77 1.52 ;
      RECT 121.6 1.462 122.005 1.52 ;
      RECT 121.6 1.41 121.98 1.52 ;
      RECT 121.6 1.365 121.945 1.52 ;
      RECT 121.6 1.347 121.91 1.52 ;
      RECT 121.6 1.337 121.905 1.52 ;
      RECT 121.32 2.295 121.51 2.52 ;
      RECT 121.31 2.296 121.515 2.515 ;
      RECT 121.31 2.298 121.525 2.495 ;
      RECT 121.31 2.302 121.53 2.48 ;
      RECT 121.31 2.289 121.48 2.515 ;
      RECT 121.31 2.292 121.505 2.515 ;
      RECT 121.32 2.288 121.48 2.52 ;
      RECT 121.406 2.286 121.48 2.52 ;
      RECT 121.03 1.537 121.2 1.775 ;
      RECT 121.03 1.537 121.286 1.689 ;
      RECT 121.03 1.537 121.29 1.599 ;
      RECT 121.08 1.31 121.3 1.578 ;
      RECT 121.075 1.327 121.305 1.551 ;
      RECT 121.04 1.485 121.305 1.551 ;
      RECT 121.06 1.335 121.2 1.775 ;
      RECT 121.05 1.417 121.31 1.534 ;
      RECT 121.045 1.465 121.31 1.534 ;
      RECT 121.05 1.375 121.305 1.551 ;
      RECT 121.075 1.312 121.3 1.578 ;
      RECT 120.64 1.287 120.81 1.485 ;
      RECT 120.64 1.287 120.855 1.46 ;
      RECT 120.71 1.23 120.88 1.418 ;
      RECT 120.685 1.245 120.88 1.418 ;
      RECT 120.3 1.291 120.33 1.485 ;
      RECT 120.295 1.263 120.3 1.485 ;
      RECT 120.265 1.237 120.295 1.487 ;
      RECT 120.24 1.195 120.265 1.49 ;
      RECT 120.23 1.167 120.24 1.492 ;
      RECT 120.195 1.147 120.23 1.494 ;
      RECT 120.13 1.132 120.195 1.5 ;
      RECT 120.08 1.13 120.13 1.506 ;
      RECT 120.057 1.132 120.08 1.511 ;
      RECT 119.971 1.143 120.057 1.517 ;
      RECT 119.885 1.161 119.971 1.527 ;
      RECT 119.87 1.172 119.885 1.533 ;
      RECT 119.8 1.195 119.87 1.539 ;
      RECT 119.745 1.227 119.8 1.547 ;
      RECT 119.705 1.25 119.745 1.553 ;
      RECT 119.691 1.263 119.705 1.556 ;
      RECT 119.605 1.285 119.691 1.562 ;
      RECT 119.59 1.31 119.605 1.568 ;
      RECT 119.55 1.325 119.59 1.572 ;
      RECT 119.5 1.34 119.55 1.577 ;
      RECT 119.475 1.347 119.5 1.581 ;
      RECT 119.415 1.342 119.475 1.585 ;
      RECT 119.4 1.333 119.415 1.589 ;
      RECT 119.33 1.323 119.4 1.585 ;
      RECT 119.305 1.315 119.325 1.575 ;
      RECT 119.246 1.315 119.305 1.553 ;
      RECT 119.16 1.315 119.246 1.51 ;
      RECT 119.325 1.315 119.33 1.58 ;
      RECT 120.02 0.546 120.19 0.88 ;
      RECT 119.99 0.546 120.19 0.875 ;
      RECT 119.93 0.513 119.99 0.863 ;
      RECT 119.93 0.569 120.2 0.858 ;
      RECT 119.905 0.569 120.2 0.852 ;
      RECT 119.9 0.51 119.93 0.849 ;
      RECT 119.885 0.516 120.02 0.847 ;
      RECT 119.88 0.524 120.105 0.835 ;
      RECT 119.88 0.576 120.215 0.788 ;
      RECT 119.865 0.532 120.105 0.783 ;
      RECT 119.865 0.602 120.225 0.724 ;
      RECT 119.835 0.552 120.19 0.685 ;
      RECT 119.835 0.642 120.235 0.681 ;
      RECT 119.885 0.521 120.105 0.847 ;
      RECT 119.225 0.851 119.28 1.115 ;
      RECT 119.225 0.851 119.345 1.114 ;
      RECT 119.225 0.851 119.37 1.113 ;
      RECT 119.225 0.851 119.435 1.112 ;
      RECT 119.37 0.817 119.45 1.111 ;
      RECT 119.185 0.861 119.595 1.11 ;
      RECT 119.225 0.858 119.595 1.11 ;
      RECT 119.185 0.866 119.6 1.103 ;
      RECT 119.17 0.868 119.6 1.102 ;
      RECT 119.17 0.875 119.605 1.098 ;
      RECT 119.15 0.874 119.6 1.094 ;
      RECT 119.15 0.882 119.61 1.093 ;
      RECT 119.145 0.879 119.605 1.089 ;
      RECT 119.145 0.892 119.62 1.088 ;
      RECT 119.13 0.882 119.61 1.087 ;
      RECT 119.095 0.895 119.62 1.08 ;
      RECT 119.28 0.85 119.59 1.11 ;
      RECT 119.28 0.835 119.54 1.11 ;
      RECT 119.345 0.822 119.475 1.11 ;
      RECT 118.89 1.911 118.905 2.304 ;
      RECT 118.855 1.916 118.905 2.303 ;
      RECT 118.89 1.915 118.95 2.302 ;
      RECT 118.835 1.926 118.95 2.301 ;
      RECT 118.85 1.922 118.95 2.301 ;
      RECT 118.815 1.932 119.025 2.298 ;
      RECT 118.815 1.951 119.07 2.296 ;
      RECT 118.815 1.958 119.075 2.293 ;
      RECT 118.8 1.935 119.025 2.29 ;
      RECT 118.78 1.94 119.025 2.283 ;
      RECT 118.775 1.944 119.025 2.279 ;
      RECT 118.775 1.961 119.085 2.278 ;
      RECT 118.755 1.955 119.07 2.274 ;
      RECT 118.755 1.964 119.09 2.268 ;
      RECT 118.75 1.97 119.09 2.04 ;
      RECT 118.815 1.93 118.95 2.298 ;
      RECT 118.69 1.293 118.89 1.605 ;
      RECT 118.765 1.271 118.89 1.605 ;
      RECT 118.705 1.29 118.895 1.59 ;
      RECT 118.675 1.301 118.895 1.588 ;
      RECT 118.69 1.296 118.9 1.554 ;
      RECT 118.675 1.4 118.905 1.521 ;
      RECT 118.705 1.272 118.89 1.605 ;
      RECT 118.765 1.25 118.865 1.605 ;
      RECT 118.79 1.247 118.865 1.605 ;
      RECT 118.79 1.242 118.81 1.605 ;
      RECT 118.195 1.31 118.37 1.485 ;
      RECT 118.19 1.31 118.37 1.483 ;
      RECT 118.165 1.31 118.37 1.478 ;
      RECT 118.11 1.29 118.28 1.468 ;
      RECT 118.11 1.297 118.345 1.468 ;
      RECT 118.195 1.977 118.21 2.16 ;
      RECT 118.185 1.955 118.195 2.16 ;
      RECT 118.17 1.935 118.185 2.16 ;
      RECT 118.16 1.91 118.17 2.16 ;
      RECT 118.13 1.875 118.16 2.16 ;
      RECT 118.095 1.815 118.13 2.16 ;
      RECT 118.09 1.777 118.095 2.16 ;
      RECT 118.04 1.728 118.09 2.16 ;
      RECT 118.03 1.678 118.04 2.148 ;
      RECT 118.015 1.657 118.03 2.108 ;
      RECT 117.995 1.625 118.015 2.058 ;
      RECT 117.97 1.581 117.995 1.998 ;
      RECT 117.965 1.553 117.97 1.953 ;
      RECT 117.96 1.544 117.965 1.939 ;
      RECT 117.955 1.537 117.96 1.926 ;
      RECT 117.95 1.532 117.955 1.915 ;
      RECT 117.945 1.517 117.95 1.905 ;
      RECT 117.94 1.495 117.945 1.892 ;
      RECT 117.93 1.455 117.94 1.867 ;
      RECT 117.905 1.385 117.93 1.823 ;
      RECT 117.9 1.325 117.905 1.788 ;
      RECT 117.885 1.305 117.9 1.755 ;
      RECT 117.88 1.305 117.885 1.73 ;
      RECT 117.85 1.305 117.88 1.685 ;
      RECT 117.805 1.305 117.85 1.625 ;
      RECT 117.73 1.305 117.805 1.573 ;
      RECT 117.725 1.305 117.73 1.538 ;
      RECT 117.72 1.305 117.725 1.528 ;
      RECT 117.715 1.305 117.72 1.508 ;
      RECT 117.98 0.525 118.15 0.995 ;
      RECT 117.925 0.518 118.12 0.979 ;
      RECT 117.925 0.532 118.155 0.978 ;
      RECT 117.91 0.533 118.155 0.959 ;
      RECT 117.905 0.551 118.155 0.945 ;
      RECT 117.91 0.534 118.16 0.943 ;
      RECT 117.895 0.565 118.16 0.928 ;
      RECT 117.91 0.54 118.165 0.913 ;
      RECT 117.89 0.58 118.165 0.91 ;
      RECT 117.905 0.552 118.17 0.895 ;
      RECT 117.905 0.564 118.175 0.875 ;
      RECT 117.89 0.58 118.18 0.858 ;
      RECT 117.89 0.59 118.185 0.713 ;
      RECT 117.885 0.59 118.185 0.67 ;
      RECT 117.885 0.605 118.19 0.648 ;
      RECT 117.98 0.515 118.12 0.995 ;
      RECT 117.98 0.513 118.09 0.995 ;
      RECT 118.066 0.51 118.09 0.995 ;
      RECT 117.725 2.177 117.73 2.223 ;
      RECT 117.715 2.025 117.725 2.247 ;
      RECT 117.71 1.87 117.715 2.272 ;
      RECT 117.695 1.832 117.71 2.283 ;
      RECT 117.69 1.815 117.695 2.29 ;
      RECT 117.68 1.803 117.69 2.297 ;
      RECT 117.675 1.794 117.68 2.299 ;
      RECT 117.67 1.792 117.675 2.303 ;
      RECT 117.625 1.783 117.67 2.318 ;
      RECT 117.62 1.775 117.625 2.332 ;
      RECT 117.615 1.772 117.62 2.336 ;
      RECT 117.6 1.767 117.615 2.344 ;
      RECT 117.545 1.757 117.6 2.355 ;
      RECT 117.51 1.745 117.545 2.356 ;
      RECT 117.501 1.74 117.51 2.35 ;
      RECT 117.415 1.74 117.501 2.34 ;
      RECT 117.385 1.74 117.415 2.318 ;
      RECT 117.375 1.74 117.38 2.298 ;
      RECT 117.37 1.74 117.375 2.26 ;
      RECT 117.365 1.74 117.37 2.218 ;
      RECT 117.36 1.74 117.365 2.178 ;
      RECT 117.355 1.74 117.36 2.108 ;
      RECT 117.345 1.74 117.355 2.03 ;
      RECT 117.34 1.74 117.345 1.93 ;
      RECT 117.38 1.74 117.385 2.3 ;
      RECT 116.875 1.822 116.965 2.3 ;
      RECT 116.86 1.825 116.98 2.298 ;
      RECT 116.875 1.824 116.98 2.298 ;
      RECT 116.84 1.831 117.005 2.288 ;
      RECT 116.86 1.825 117.005 2.288 ;
      RECT 116.825 1.837 117.005 2.276 ;
      RECT 116.86 1.828 117.055 2.269 ;
      RECT 116.811 1.845 117.055 2.267 ;
      RECT 116.84 1.835 117.065 2.255 ;
      RECT 116.811 1.856 117.095 2.246 ;
      RECT 116.725 1.88 117.095 2.24 ;
      RECT 116.725 1.893 117.135 2.223 ;
      RECT 116.72 1.915 117.135 2.216 ;
      RECT 116.69 1.93 117.135 2.206 ;
      RECT 116.685 1.941 117.135 2.196 ;
      RECT 116.655 1.954 117.135 2.187 ;
      RECT 116.64 1.972 117.135 2.176 ;
      RECT 116.615 1.985 117.135 2.166 ;
      RECT 116.875 1.821 116.885 2.3 ;
      RECT 116.921 1.245 116.96 1.49 ;
      RECT 116.835 1.245 116.97 1.488 ;
      RECT 116.72 1.27 116.97 1.485 ;
      RECT 116.72 1.27 116.975 1.483 ;
      RECT 116.72 1.27 116.99 1.478 ;
      RECT 116.826 1.245 117.005 1.458 ;
      RECT 116.74 1.253 117.005 1.458 ;
      RECT 116.41 0.605 116.58 1.04 ;
      RECT 116.4 0.639 116.58 1.023 ;
      RECT 116.48 0.575 116.65 1.01 ;
      RECT 116.385 0.65 116.65 0.988 ;
      RECT 116.48 0.585 116.655 0.978 ;
      RECT 116.41 0.637 116.685 0.963 ;
      RECT 116.37 0.663 116.685 0.948 ;
      RECT 116.37 0.705 116.695 0.928 ;
      RECT 116.365 0.73 116.7 0.91 ;
      RECT 116.365 0.74 116.705 0.895 ;
      RECT 116.36 0.677 116.685 0.893 ;
      RECT 116.36 0.75 116.71 0.878 ;
      RECT 116.355 0.687 116.685 0.875 ;
      RECT 116.35 0.771 116.715 0.858 ;
      RECT 116.35 0.803 116.72 0.838 ;
      RECT 116.345 0.717 116.695 0.83 ;
      RECT 116.35 0.702 116.685 0.858 ;
      RECT 116.365 0.672 116.685 0.91 ;
      RECT 116.21 1.259 116.435 1.515 ;
      RECT 116.21 1.292 116.455 1.505 ;
      RECT 116.175 1.292 116.455 1.503 ;
      RECT 116.175 1.305 116.46 1.493 ;
      RECT 116.175 1.325 116.47 1.485 ;
      RECT 116.175 1.422 116.475 1.478 ;
      RECT 116.155 1.17 116.285 1.468 ;
      RECT 116.11 1.325 116.47 1.41 ;
      RECT 116.1 1.17 116.285 1.355 ;
      RECT 116.1 1.202 116.371 1.355 ;
      RECT 116.065 1.732 116.085 1.91 ;
      RECT 116.03 1.685 116.065 1.91 ;
      RECT 116.015 1.625 116.03 1.91 ;
      RECT 115.99 1.572 116.015 1.91 ;
      RECT 115.975 1.525 115.99 1.91 ;
      RECT 115.955 1.502 115.975 1.91 ;
      RECT 115.93 1.467 115.955 1.91 ;
      RECT 115.92 1.313 115.93 1.91 ;
      RECT 115.89 1.308 115.92 1.901 ;
      RECT 115.885 1.305 115.89 1.891 ;
      RECT 115.87 1.305 115.885 1.865 ;
      RECT 115.865 1.305 115.87 1.828 ;
      RECT 115.84 1.305 115.865 1.78 ;
      RECT 115.82 1.305 115.84 1.705 ;
      RECT 115.81 1.305 115.82 1.665 ;
      RECT 115.805 1.305 115.81 1.64 ;
      RECT 115.8 1.305 115.805 1.623 ;
      RECT 115.795 1.305 115.8 1.605 ;
      RECT 115.79 1.306 115.795 1.595 ;
      RECT 115.78 1.308 115.79 1.563 ;
      RECT 115.77 1.31 115.78 1.53 ;
      RECT 115.76 1.313 115.77 1.503 ;
      RECT 116.085 1.74 116.31 1.91 ;
      RECT 115.415 0.552 115.585 1.005 ;
      RECT 115.415 0.552 115.675 0.971 ;
      RECT 115.415 0.552 115.705 0.955 ;
      RECT 115.415 0.552 115.735 0.928 ;
      RECT 115.671 0.53 115.75 0.91 ;
      RECT 115.45 0.537 115.755 0.895 ;
      RECT 115.45 0.545 115.765 0.858 ;
      RECT 115.41 0.572 115.765 0.83 ;
      RECT 115.395 0.585 115.765 0.795 ;
      RECT 115.415 0.56 115.785 0.785 ;
      RECT 115.39 0.625 115.785 0.755 ;
      RECT 115.39 0.655 115.79 0.738 ;
      RECT 115.385 0.685 115.79 0.725 ;
      RECT 115.45 0.534 115.75 0.91 ;
      RECT 115.585 0.531 115.671 0.989 ;
      RECT 115.536 0.532 115.75 0.91 ;
      RECT 115.68 2.192 115.725 2.385 ;
      RECT 115.67 2.162 115.68 2.385 ;
      RECT 115.665 2.147 115.67 2.385 ;
      RECT 115.625 2.057 115.665 2.385 ;
      RECT 115.62 1.97 115.625 2.385 ;
      RECT 115.61 1.94 115.62 2.385 ;
      RECT 115.605 1.9 115.61 2.385 ;
      RECT 115.595 1.862 115.605 2.385 ;
      RECT 115.59 1.827 115.595 2.385 ;
      RECT 115.57 1.78 115.59 2.385 ;
      RECT 115.555 1.705 115.57 2.385 ;
      RECT 115.55 1.66 115.555 2.38 ;
      RECT 115.545 1.64 115.55 2.353 ;
      RECT 115.54 1.62 115.545 2.338 ;
      RECT 115.535 1.595 115.54 2.318 ;
      RECT 115.53 1.573 115.535 2.303 ;
      RECT 115.525 1.551 115.53 2.285 ;
      RECT 115.52 1.53 115.525 2.275 ;
      RECT 115.51 1.502 115.52 2.245 ;
      RECT 115.5 1.465 115.51 2.213 ;
      RECT 115.49 1.425 115.5 2.18 ;
      RECT 115.48 1.403 115.49 2.15 ;
      RECT 115.45 1.355 115.48 2.082 ;
      RECT 115.435 1.315 115.45 2.009 ;
      RECT 115.425 1.315 115.435 1.975 ;
      RECT 115.42 1.315 115.425 1.95 ;
      RECT 115.415 1.315 115.42 1.935 ;
      RECT 115.41 1.315 115.415 1.913 ;
      RECT 115.405 1.315 115.41 1.9 ;
      RECT 115.39 1.315 115.405 1.865 ;
      RECT 115.37 1.315 115.39 1.805 ;
      RECT 115.36 1.315 115.37 1.755 ;
      RECT 115.34 1.315 115.36 1.703 ;
      RECT 115.32 1.315 115.34 1.66 ;
      RECT 115.31 1.315 115.32 1.648 ;
      RECT 115.28 1.315 115.31 1.635 ;
      RECT 115.25 1.336 115.28 1.615 ;
      RECT 115.24 1.364 115.25 1.595 ;
      RECT 115.225 1.381 115.24 1.563 ;
      RECT 115.22 1.395 115.225 1.53 ;
      RECT 115.215 1.403 115.22 1.503 ;
      RECT 115.21 1.411 115.215 1.465 ;
      RECT 115.215 1.935 115.22 2.27 ;
      RECT 115.18 1.922 115.215 2.269 ;
      RECT 115.11 1.862 115.18 2.268 ;
      RECT 115.03 1.805 115.11 2.267 ;
      RECT 114.895 1.765 115.03 2.266 ;
      RECT 114.895 1.952 115.23 2.255 ;
      RECT 114.855 1.952 115.23 2.245 ;
      RECT 114.855 1.97 115.235 2.24 ;
      RECT 114.855 2.06 115.24 2.23 ;
      RECT 114.85 1.755 115.015 2.21 ;
      RECT 114.845 1.755 115.015 1.953 ;
      RECT 114.845 1.912 115.21 1.953 ;
      RECT 114.845 1.9 115.205 1.953 ;
      RECT 114.11 2.115 114.625 2.525 ;
      RECT 114.285 1.135 114.625 2.525 ;
      RECT 113.395 1.135 114.625 1.305 ;
      RECT 114.105 0.53 114.35 1.305 ;
      RECT 111.505 2.535 113.535 2.705 ;
      RECT 113.365 1.68 113.535 2.705 ;
      RECT 111.505 1.235 111.675 2.705 ;
      RECT 113.365 1.68 114.115 1.87 ;
      RECT 111.48 1.235 111.675 1.565 ;
      RECT 112.185 1.855 113.195 2.025 ;
      RECT 113.005 0.495 113.195 2.025 ;
      RECT 112.185 1.055 112.355 2.025 ;
      RECT 111.845 2.195 112.97 2.365 ;
      RECT 111.845 0.495 112.015 2.365 ;
      RECT 111 1.235 111.255 1.565 ;
      RECT 111.085 0.895 111.255 1.565 ;
      RECT 111.085 0.895 112.015 1.065 ;
      RECT 111.84 0.495 112.015 1.065 ;
      RECT 111.84 0.495 112.37 0.86 ;
      RECT 110.66 1.735 110.995 2.705 ;
      RECT 110.66 0.495 110.83 2.705 ;
      RECT 110.66 0.495 110.915 1.065 ;
      RECT 109.91 1.725 110.24 2.705 ;
      RECT 110.01 0.495 110.24 2.705 ;
      RECT 109.91 0.495 110.24 1.125 ;
      RECT 108.53 1.725 108.86 2.705 ;
      RECT 108.63 0.495 108.86 2.705 ;
      RECT 108.63 1.315 109.84 1.555 ;
      RECT 108.53 0.495 108.86 1.125 ;
      RECT 107.15 1.725 107.48 2.705 ;
      RECT 107.25 0.495 107.48 2.705 ;
      RECT 107.15 0.495 107.48 1.125 ;
      RECT 105.77 1.725 106.1 2.705 ;
      RECT 105.87 0.495 106.1 2.705 ;
      RECT 105.87 1.315 107.08 1.555 ;
      RECT 105.77 0.495 106.1 1.125 ;
      RECT 104.45 2.115 104.965 2.525 ;
      RECT 104.625 1.135 104.965 2.525 ;
      RECT 103.735 1.135 104.965 1.305 ;
      RECT 104.445 0.53 104.69 1.305 ;
      RECT 101.845 2.535 103.875 2.705 ;
      RECT 103.705 1.68 103.875 2.705 ;
      RECT 101.845 1.235 102.015 2.705 ;
      RECT 103.705 1.68 104.455 1.87 ;
      RECT 101.82 1.235 102.015 1.565 ;
      RECT 102.525 1.855 103.535 2.025 ;
      RECT 103.345 0.495 103.535 2.025 ;
      RECT 102.525 1.055 102.695 2.025 ;
      RECT 102.185 2.195 103.31 2.365 ;
      RECT 102.185 0.495 102.355 2.365 ;
      RECT 101.34 1.235 101.595 1.565 ;
      RECT 101.425 0.895 101.595 1.565 ;
      RECT 101.425 0.895 102.355 1.065 ;
      RECT 102.18 0.495 102.355 1.065 ;
      RECT 102.18 0.495 102.71 0.86 ;
      RECT 101 1.735 101.335 2.705 ;
      RECT 101 0.495 101.17 2.705 ;
      RECT 101 0.495 101.255 1.065 ;
      RECT 100.315 2.115 100.83 2.525 ;
      RECT 100.49 1.135 100.83 2.525 ;
      RECT 99.6 1.135 100.83 1.305 ;
      RECT 100.31 0.53 100.555 1.305 ;
      RECT 97.71 2.535 99.74 2.705 ;
      RECT 99.57 1.68 99.74 2.705 ;
      RECT 97.71 1.235 97.88 2.705 ;
      RECT 99.57 1.68 100.32 1.87 ;
      RECT 97.685 1.235 97.88 1.565 ;
      RECT 98.39 1.855 99.4 2.025 ;
      RECT 99.21 0.495 99.4 2.025 ;
      RECT 98.39 1.055 98.56 2.025 ;
      RECT 98.05 2.195 99.175 2.365 ;
      RECT 98.05 0.495 98.22 2.365 ;
      RECT 97.205 1.235 97.46 1.565 ;
      RECT 97.29 0.895 97.46 1.565 ;
      RECT 97.29 0.895 98.22 1.065 ;
      RECT 98.045 0.495 98.22 1.065 ;
      RECT 98.045 0.495 98.575 0.86 ;
      RECT 96.865 1.735 97.2 2.705 ;
      RECT 96.865 0.495 97.035 2.705 ;
      RECT 96.865 0.495 97.12 1.065 ;
      RECT 95.77 0.715 96.5 0.955 ;
      RECT 96.312 0.51 96.5 0.955 ;
      RECT 96.14 0.522 96.515 0.949 ;
      RECT 96.055 0.537 96.535 0.934 ;
      RECT 96.055 0.552 96.54 0.924 ;
      RECT 96.01 0.572 96.555 0.916 ;
      RECT 95.987 0.607 96.57 0.87 ;
      RECT 95.901 0.63 96.575 0.83 ;
      RECT 95.901 0.648 96.585 0.8 ;
      RECT 95.77 0.717 96.59 0.763 ;
      RECT 95.815 0.66 96.585 0.8 ;
      RECT 95.901 0.612 96.57 0.87 ;
      RECT 95.987 0.581 96.555 0.916 ;
      RECT 96.01 0.562 96.54 0.924 ;
      RECT 96.055 0.535 96.515 0.949 ;
      RECT 96.14 0.517 96.5 0.955 ;
      RECT 96.226 0.511 96.5 0.955 ;
      RECT 96.312 0.506 96.445 0.955 ;
      RECT 96.398 0.501 96.445 0.955 ;
      RECT 96.09 1.399 96.26 1.785 ;
      RECT 96.085 1.399 96.26 1.78 ;
      RECT 96.06 1.399 96.26 1.745 ;
      RECT 96.06 1.427 96.27 1.735 ;
      RECT 96.04 1.427 96.27 1.695 ;
      RECT 96.035 1.427 96.27 1.668 ;
      RECT 96.035 1.445 96.275 1.66 ;
      RECT 95.98 1.445 96.275 1.595 ;
      RECT 95.98 1.462 96.285 1.578 ;
      RECT 95.97 1.462 96.285 1.518 ;
      RECT 95.97 1.479 96.29 1.515 ;
      RECT 95.965 1.315 96.135 1.493 ;
      RECT 95.965 1.349 96.221 1.493 ;
      RECT 95.96 2.115 95.965 2.128 ;
      RECT 95.955 2.01 95.96 2.133 ;
      RECT 95.93 1.87 95.955 2.148 ;
      RECT 95.895 1.821 95.93 2.18 ;
      RECT 95.89 1.789 95.895 2.2 ;
      RECT 95.885 1.78 95.89 2.2 ;
      RECT 95.805 1.745 95.885 2.2 ;
      RECT 95.742 1.715 95.805 2.2 ;
      RECT 95.656 1.703 95.742 2.2 ;
      RECT 95.57 1.689 95.656 2.2 ;
      RECT 95.49 1.676 95.57 2.186 ;
      RECT 95.455 1.668 95.49 2.166 ;
      RECT 95.445 1.665 95.455 2.157 ;
      RECT 95.415 1.66 95.445 2.144 ;
      RECT 95.365 1.635 95.415 2.12 ;
      RECT 95.351 1.609 95.365 2.102 ;
      RECT 95.265 1.569 95.351 2.078 ;
      RECT 95.22 1.517 95.265 2.047 ;
      RECT 95.21 1.492 95.22 2.034 ;
      RECT 95.205 1.273 95.21 1.295 ;
      RECT 95.2 1.475 95.21 2.03 ;
      RECT 95.2 1.271 95.205 1.385 ;
      RECT 95.19 1.267 95.2 2.026 ;
      RECT 95.146 1.265 95.19 2.014 ;
      RECT 95.06 1.265 95.146 1.985 ;
      RECT 95.03 1.265 95.06 1.958 ;
      RECT 95.015 1.265 95.03 1.946 ;
      RECT 94.975 1.277 95.015 1.931 ;
      RECT 94.955 1.296 94.975 1.91 ;
      RECT 94.945 1.306 94.955 1.894 ;
      RECT 94.935 1.312 94.945 1.883 ;
      RECT 94.915 1.322 94.935 1.866 ;
      RECT 94.91 1.331 94.915 1.853 ;
      RECT 94.905 1.335 94.91 1.803 ;
      RECT 94.895 1.341 94.905 1.72 ;
      RECT 94.89 1.345 94.895 1.634 ;
      RECT 94.885 1.365 94.89 1.571 ;
      RECT 94.88 1.388 94.885 1.518 ;
      RECT 94.875 1.406 94.88 1.463 ;
      RECT 95.485 1.225 95.655 1.485 ;
      RECT 95.655 1.19 95.7 1.471 ;
      RECT 95.616 1.192 95.705 1.454 ;
      RECT 95.505 1.209 95.791 1.425 ;
      RECT 95.505 1.224 95.795 1.397 ;
      RECT 95.505 1.205 95.705 1.454 ;
      RECT 95.53 1.193 95.655 1.485 ;
      RECT 95.616 1.191 95.7 1.471 ;
      RECT 94.67 0.58 94.84 1.07 ;
      RECT 94.67 0.58 94.875 1.05 ;
      RECT 94.805 0.5 94.915 1.01 ;
      RECT 94.786 0.504 94.935 0.98 ;
      RECT 94.7 0.512 94.955 0.963 ;
      RECT 94.7 0.518 94.96 0.953 ;
      RECT 94.7 0.527 94.98 0.941 ;
      RECT 94.675 0.552 95.01 0.919 ;
      RECT 94.675 0.572 95.015 0.899 ;
      RECT 94.67 0.585 95.025 0.879 ;
      RECT 94.67 0.652 95.03 0.86 ;
      RECT 94.67 0.785 95.035 0.847 ;
      RECT 94.665 0.59 95.025 0.68 ;
      RECT 94.675 0.547 94.98 0.941 ;
      RECT 94.786 0.502 94.915 1.01 ;
      RECT 94.66 2.255 94.96 2.51 ;
      RECT 94.745 2.221 94.96 2.51 ;
      RECT 94.745 2.224 94.965 2.37 ;
      RECT 94.68 2.245 94.965 2.37 ;
      RECT 94.715 2.235 94.96 2.51 ;
      RECT 94.71 2.24 94.965 2.37 ;
      RECT 94.745 2.219 94.946 2.51 ;
      RECT 94.831 2.21 94.946 2.51 ;
      RECT 94.831 2.204 94.86 2.51 ;
      RECT 94.32 1.845 94.33 2.335 ;
      RECT 93.98 1.78 93.99 2.08 ;
      RECT 94.495 1.952 94.5 2.171 ;
      RECT 94.485 1.932 94.495 2.188 ;
      RECT 94.475 1.912 94.485 2.218 ;
      RECT 94.47 1.902 94.475 2.233 ;
      RECT 94.465 1.898 94.47 2.238 ;
      RECT 94.45 1.89 94.465 2.245 ;
      RECT 94.41 1.87 94.45 2.27 ;
      RECT 94.385 1.852 94.41 2.303 ;
      RECT 94.38 1.85 94.385 2.316 ;
      RECT 94.36 1.847 94.38 2.32 ;
      RECT 94.33 1.845 94.36 2.33 ;
      RECT 94.26 1.847 94.32 2.331 ;
      RECT 94.24 1.847 94.26 2.325 ;
      RECT 94.215 1.845 94.24 2.322 ;
      RECT 94.18 1.84 94.215 2.318 ;
      RECT 94.16 1.834 94.18 2.305 ;
      RECT 94.15 1.831 94.16 2.293 ;
      RECT 94.13 1.828 94.15 2.278 ;
      RECT 94.11 1.824 94.13 2.26 ;
      RECT 94.105 1.821 94.11 2.25 ;
      RECT 94.1 1.82 94.105 2.248 ;
      RECT 94.09 1.817 94.1 2.24 ;
      RECT 94.08 1.811 94.09 2.223 ;
      RECT 94.07 1.805 94.08 2.205 ;
      RECT 94.06 1.799 94.07 2.193 ;
      RECT 94.05 1.793 94.06 2.173 ;
      RECT 94.045 1.789 94.05 2.158 ;
      RECT 94.04 1.787 94.045 2.15 ;
      RECT 94.035 1.785 94.04 2.143 ;
      RECT 94.03 1.783 94.035 2.133 ;
      RECT 94.025 1.781 94.03 2.127 ;
      RECT 94.015 1.78 94.025 2.117 ;
      RECT 94.005 1.78 94.015 2.108 ;
      RECT 93.99 1.78 94.005 2.093 ;
      RECT 93.95 1.78 93.98 2.077 ;
      RECT 93.93 1.782 93.95 2.072 ;
      RECT 93.925 1.787 93.93 2.07 ;
      RECT 93.895 1.795 93.925 2.068 ;
      RECT 93.865 1.81 93.895 2.067 ;
      RECT 93.82 1.832 93.865 2.072 ;
      RECT 93.815 1.847 93.82 2.076 ;
      RECT 93.8 1.852 93.815 2.078 ;
      RECT 93.795 1.856 93.8 2.08 ;
      RECT 93.735 1.879 93.795 2.089 ;
      RECT 93.715 1.905 93.735 2.102 ;
      RECT 93.705 1.912 93.715 2.106 ;
      RECT 93.69 1.919 93.705 2.109 ;
      RECT 93.67 1.929 93.69 2.112 ;
      RECT 93.665 1.937 93.67 2.115 ;
      RECT 93.62 1.942 93.665 2.122 ;
      RECT 93.61 1.945 93.62 2.129 ;
      RECT 93.6 1.945 93.61 2.133 ;
      RECT 93.565 1.947 93.6 2.145 ;
      RECT 93.545 1.95 93.565 2.158 ;
      RECT 93.505 1.953 93.545 2.169 ;
      RECT 93.49 1.955 93.505 2.182 ;
      RECT 93.48 1.955 93.49 2.187 ;
      RECT 93.455 1.956 93.48 2.195 ;
      RECT 93.445 1.958 93.455 2.2 ;
      RECT 93.44 1.959 93.445 2.203 ;
      RECT 93.415 1.957 93.44 2.206 ;
      RECT 93.4 1.955 93.415 2.207 ;
      RECT 93.38 1.952 93.4 2.209 ;
      RECT 93.36 1.947 93.38 2.209 ;
      RECT 93.3 1.942 93.36 2.206 ;
      RECT 93.265 1.917 93.3 2.202 ;
      RECT 93.255 1.894 93.265 2.2 ;
      RECT 93.225 1.871 93.255 2.2 ;
      RECT 93.215 1.85 93.225 2.2 ;
      RECT 93.19 1.832 93.215 2.198 ;
      RECT 93.175 1.81 93.19 2.195 ;
      RECT 93.16 1.792 93.175 2.193 ;
      RECT 93.14 1.782 93.16 2.191 ;
      RECT 93.125 1.777 93.14 2.19 ;
      RECT 93.11 1.775 93.125 2.189 ;
      RECT 93.08 1.776 93.11 2.187 ;
      RECT 93.06 1.779 93.08 2.185 ;
      RECT 93.003 1.783 93.06 2.185 ;
      RECT 92.917 1.792 93.003 2.185 ;
      RECT 92.831 1.803 92.917 2.185 ;
      RECT 92.745 1.814 92.831 2.185 ;
      RECT 92.725 1.821 92.745 2.193 ;
      RECT 92.715 1.824 92.725 2.2 ;
      RECT 92.65 1.829 92.715 2.218 ;
      RECT 92.62 1.836 92.65 2.243 ;
      RECT 92.61 1.839 92.62 2.25 ;
      RECT 92.565 1.843 92.61 2.255 ;
      RECT 92.535 1.848 92.565 2.26 ;
      RECT 92.534 1.85 92.535 2.26 ;
      RECT 92.448 1.856 92.534 2.26 ;
      RECT 92.362 1.867 92.448 2.26 ;
      RECT 92.276 1.879 92.362 2.26 ;
      RECT 92.19 1.89 92.276 2.26 ;
      RECT 92.175 1.897 92.19 2.255 ;
      RECT 92.17 1.899 92.175 2.249 ;
      RECT 92.15 1.91 92.17 2.244 ;
      RECT 92.14 1.928 92.15 2.238 ;
      RECT 92.135 1.94 92.14 2.038 ;
      RECT 94.43 0.693 94.45 0.78 ;
      RECT 94.425 0.628 94.43 0.812 ;
      RECT 94.415 0.595 94.425 0.817 ;
      RECT 94.41 0.575 94.415 0.823 ;
      RECT 94.38 0.575 94.41 0.84 ;
      RECT 94.331 0.575 94.38 0.876 ;
      RECT 94.245 0.575 94.331 0.934 ;
      RECT 94.216 0.585 94.245 0.983 ;
      RECT 94.13 0.627 94.216 1.036 ;
      RECT 94.11 0.665 94.13 1.083 ;
      RECT 94.085 0.682 94.11 1.103 ;
      RECT 94.075 0.696 94.085 1.123 ;
      RECT 94.07 0.702 94.075 1.133 ;
      RECT 94.065 0.706 94.07 1.14 ;
      RECT 94.015 0.726 94.065 1.145 ;
      RECT 93.95 0.77 94.015 1.145 ;
      RECT 93.925 0.82 93.95 1.145 ;
      RECT 93.915 0.85 93.925 1.145 ;
      RECT 93.91 0.877 93.915 1.145 ;
      RECT 93.905 0.895 93.91 1.145 ;
      RECT 93.895 0.937 93.905 1.145 ;
      RECT 94.245 1.495 94.415 1.67 ;
      RECT 94.185 1.323 94.245 1.658 ;
      RECT 94.175 1.316 94.185 1.641 ;
      RECT 94.13 1.495 94.415 1.621 ;
      RECT 94.111 1.495 94.415 1.599 ;
      RECT 94.025 1.495 94.415 1.564 ;
      RECT 94.005 1.315 94.175 1.52 ;
      RECT 94.005 1.462 94.41 1.52 ;
      RECT 94.005 1.41 94.385 1.52 ;
      RECT 94.005 1.365 94.35 1.52 ;
      RECT 94.005 1.347 94.315 1.52 ;
      RECT 94.005 1.337 94.31 1.52 ;
      RECT 93.725 2.295 93.915 2.52 ;
      RECT 93.715 2.296 93.92 2.515 ;
      RECT 93.715 2.298 93.93 2.495 ;
      RECT 93.715 2.302 93.935 2.48 ;
      RECT 93.715 2.289 93.885 2.515 ;
      RECT 93.715 2.292 93.91 2.515 ;
      RECT 93.725 2.288 93.885 2.52 ;
      RECT 93.811 2.286 93.885 2.52 ;
      RECT 93.435 1.537 93.605 1.775 ;
      RECT 93.435 1.537 93.691 1.689 ;
      RECT 93.435 1.537 93.695 1.599 ;
      RECT 93.485 1.31 93.705 1.578 ;
      RECT 93.48 1.327 93.71 1.551 ;
      RECT 93.445 1.485 93.71 1.551 ;
      RECT 93.465 1.335 93.605 1.775 ;
      RECT 93.455 1.417 93.715 1.534 ;
      RECT 93.45 1.465 93.715 1.534 ;
      RECT 93.455 1.375 93.71 1.551 ;
      RECT 93.48 1.312 93.705 1.578 ;
      RECT 93.045 1.287 93.215 1.485 ;
      RECT 93.045 1.287 93.26 1.46 ;
      RECT 93.115 1.23 93.285 1.418 ;
      RECT 93.09 1.245 93.285 1.418 ;
      RECT 92.705 1.291 92.735 1.485 ;
      RECT 92.7 1.263 92.705 1.485 ;
      RECT 92.67 1.237 92.7 1.487 ;
      RECT 92.645 1.195 92.67 1.49 ;
      RECT 92.635 1.167 92.645 1.492 ;
      RECT 92.6 1.147 92.635 1.494 ;
      RECT 92.535 1.132 92.6 1.5 ;
      RECT 92.485 1.13 92.535 1.506 ;
      RECT 92.462 1.132 92.485 1.511 ;
      RECT 92.376 1.143 92.462 1.517 ;
      RECT 92.29 1.161 92.376 1.527 ;
      RECT 92.275 1.172 92.29 1.533 ;
      RECT 92.205 1.195 92.275 1.539 ;
      RECT 92.15 1.227 92.205 1.547 ;
      RECT 92.11 1.25 92.15 1.553 ;
      RECT 92.096 1.263 92.11 1.556 ;
      RECT 92.01 1.285 92.096 1.562 ;
      RECT 91.995 1.31 92.01 1.568 ;
      RECT 91.955 1.325 91.995 1.572 ;
      RECT 91.905 1.34 91.955 1.577 ;
      RECT 91.88 1.347 91.905 1.581 ;
      RECT 91.82 1.342 91.88 1.585 ;
      RECT 91.805 1.333 91.82 1.589 ;
      RECT 91.735 1.323 91.805 1.585 ;
      RECT 91.71 1.315 91.73 1.575 ;
      RECT 91.651 1.315 91.71 1.553 ;
      RECT 91.565 1.315 91.651 1.51 ;
      RECT 91.73 1.315 91.735 1.58 ;
      RECT 92.425 0.546 92.595 0.88 ;
      RECT 92.395 0.546 92.595 0.875 ;
      RECT 92.335 0.513 92.395 0.863 ;
      RECT 92.335 0.569 92.605 0.858 ;
      RECT 92.31 0.569 92.605 0.852 ;
      RECT 92.305 0.51 92.335 0.849 ;
      RECT 92.29 0.516 92.425 0.847 ;
      RECT 92.285 0.524 92.51 0.835 ;
      RECT 92.285 0.576 92.62 0.788 ;
      RECT 92.27 0.532 92.51 0.783 ;
      RECT 92.27 0.602 92.63 0.724 ;
      RECT 92.24 0.552 92.595 0.685 ;
      RECT 92.24 0.642 92.64 0.681 ;
      RECT 92.29 0.521 92.51 0.847 ;
      RECT 91.63 0.851 91.685 1.115 ;
      RECT 91.63 0.851 91.75 1.114 ;
      RECT 91.63 0.851 91.775 1.113 ;
      RECT 91.63 0.851 91.84 1.112 ;
      RECT 91.775 0.817 91.855 1.111 ;
      RECT 91.59 0.861 92 1.11 ;
      RECT 91.63 0.858 92 1.11 ;
      RECT 91.59 0.866 92.005 1.103 ;
      RECT 91.575 0.868 92.005 1.102 ;
      RECT 91.575 0.875 92.01 1.098 ;
      RECT 91.555 0.874 92.005 1.094 ;
      RECT 91.555 0.882 92.015 1.093 ;
      RECT 91.55 0.879 92.01 1.089 ;
      RECT 91.55 0.892 92.025 1.088 ;
      RECT 91.535 0.882 92.015 1.087 ;
      RECT 91.5 0.895 92.025 1.08 ;
      RECT 91.685 0.85 91.995 1.11 ;
      RECT 91.685 0.835 91.945 1.11 ;
      RECT 91.75 0.822 91.88 1.11 ;
      RECT 91.295 1.911 91.31 2.304 ;
      RECT 91.26 1.916 91.31 2.303 ;
      RECT 91.295 1.915 91.355 2.302 ;
      RECT 91.24 1.926 91.355 2.301 ;
      RECT 91.255 1.922 91.355 2.301 ;
      RECT 91.22 1.932 91.43 2.298 ;
      RECT 91.22 1.951 91.475 2.296 ;
      RECT 91.22 1.958 91.48 2.293 ;
      RECT 91.205 1.935 91.43 2.29 ;
      RECT 91.185 1.94 91.43 2.283 ;
      RECT 91.18 1.944 91.43 2.279 ;
      RECT 91.18 1.961 91.49 2.278 ;
      RECT 91.16 1.955 91.475 2.274 ;
      RECT 91.16 1.964 91.495 2.268 ;
      RECT 91.155 1.97 91.495 2.04 ;
      RECT 91.22 1.93 91.355 2.298 ;
      RECT 91.095 1.293 91.295 1.605 ;
      RECT 91.17 1.271 91.295 1.605 ;
      RECT 91.11 1.29 91.3 1.59 ;
      RECT 91.08 1.301 91.3 1.588 ;
      RECT 91.095 1.296 91.305 1.554 ;
      RECT 91.08 1.4 91.31 1.521 ;
      RECT 91.11 1.272 91.295 1.605 ;
      RECT 91.17 1.25 91.27 1.605 ;
      RECT 91.195 1.247 91.27 1.605 ;
      RECT 91.195 1.242 91.215 1.605 ;
      RECT 90.6 1.31 90.775 1.485 ;
      RECT 90.595 1.31 90.775 1.483 ;
      RECT 90.57 1.31 90.775 1.478 ;
      RECT 90.515 1.29 90.685 1.468 ;
      RECT 90.515 1.297 90.75 1.468 ;
      RECT 90.6 1.977 90.615 2.16 ;
      RECT 90.59 1.955 90.6 2.16 ;
      RECT 90.575 1.935 90.59 2.16 ;
      RECT 90.565 1.91 90.575 2.16 ;
      RECT 90.535 1.875 90.565 2.16 ;
      RECT 90.5 1.815 90.535 2.16 ;
      RECT 90.495 1.777 90.5 2.16 ;
      RECT 90.445 1.728 90.495 2.16 ;
      RECT 90.435 1.678 90.445 2.148 ;
      RECT 90.42 1.657 90.435 2.108 ;
      RECT 90.4 1.625 90.42 2.058 ;
      RECT 90.375 1.581 90.4 1.998 ;
      RECT 90.37 1.553 90.375 1.953 ;
      RECT 90.365 1.544 90.37 1.939 ;
      RECT 90.36 1.537 90.365 1.926 ;
      RECT 90.355 1.532 90.36 1.915 ;
      RECT 90.35 1.517 90.355 1.905 ;
      RECT 90.345 1.495 90.35 1.892 ;
      RECT 90.335 1.455 90.345 1.867 ;
      RECT 90.31 1.385 90.335 1.823 ;
      RECT 90.305 1.325 90.31 1.788 ;
      RECT 90.29 1.305 90.305 1.755 ;
      RECT 90.285 1.305 90.29 1.73 ;
      RECT 90.255 1.305 90.285 1.685 ;
      RECT 90.21 1.305 90.255 1.625 ;
      RECT 90.135 1.305 90.21 1.573 ;
      RECT 90.13 1.305 90.135 1.538 ;
      RECT 90.125 1.305 90.13 1.528 ;
      RECT 90.12 1.305 90.125 1.508 ;
      RECT 90.385 0.525 90.555 0.995 ;
      RECT 90.33 0.518 90.525 0.979 ;
      RECT 90.33 0.532 90.56 0.978 ;
      RECT 90.315 0.533 90.56 0.959 ;
      RECT 90.31 0.551 90.56 0.945 ;
      RECT 90.315 0.534 90.565 0.943 ;
      RECT 90.3 0.565 90.565 0.928 ;
      RECT 90.315 0.54 90.57 0.913 ;
      RECT 90.295 0.58 90.57 0.91 ;
      RECT 90.31 0.552 90.575 0.895 ;
      RECT 90.31 0.564 90.58 0.875 ;
      RECT 90.295 0.58 90.585 0.858 ;
      RECT 90.295 0.59 90.59 0.713 ;
      RECT 90.29 0.59 90.59 0.67 ;
      RECT 90.29 0.605 90.595 0.648 ;
      RECT 90.385 0.515 90.525 0.995 ;
      RECT 90.385 0.513 90.495 0.995 ;
      RECT 90.471 0.51 90.495 0.995 ;
      RECT 90.13 2.177 90.135 2.223 ;
      RECT 90.12 2.025 90.13 2.247 ;
      RECT 90.115 1.87 90.12 2.272 ;
      RECT 90.1 1.832 90.115 2.283 ;
      RECT 90.095 1.815 90.1 2.29 ;
      RECT 90.085 1.803 90.095 2.297 ;
      RECT 90.08 1.794 90.085 2.299 ;
      RECT 90.075 1.792 90.08 2.303 ;
      RECT 90.03 1.783 90.075 2.318 ;
      RECT 90.025 1.775 90.03 2.332 ;
      RECT 90.02 1.772 90.025 2.336 ;
      RECT 90.005 1.767 90.02 2.344 ;
      RECT 89.95 1.757 90.005 2.355 ;
      RECT 89.915 1.745 89.95 2.356 ;
      RECT 89.906 1.74 89.915 2.35 ;
      RECT 89.82 1.74 89.906 2.34 ;
      RECT 89.79 1.74 89.82 2.318 ;
      RECT 89.78 1.74 89.785 2.298 ;
      RECT 89.775 1.74 89.78 2.26 ;
      RECT 89.77 1.74 89.775 2.218 ;
      RECT 89.765 1.74 89.77 2.178 ;
      RECT 89.76 1.74 89.765 2.108 ;
      RECT 89.75 1.74 89.76 2.03 ;
      RECT 89.745 1.74 89.75 1.93 ;
      RECT 89.785 1.74 89.79 2.3 ;
      RECT 89.28 1.822 89.37 2.3 ;
      RECT 89.265 1.825 89.385 2.298 ;
      RECT 89.28 1.824 89.385 2.298 ;
      RECT 89.245 1.831 89.41 2.288 ;
      RECT 89.265 1.825 89.41 2.288 ;
      RECT 89.23 1.837 89.41 2.276 ;
      RECT 89.265 1.828 89.46 2.269 ;
      RECT 89.216 1.845 89.46 2.267 ;
      RECT 89.245 1.835 89.47 2.255 ;
      RECT 89.216 1.856 89.5 2.246 ;
      RECT 89.13 1.88 89.5 2.24 ;
      RECT 89.13 1.893 89.54 2.223 ;
      RECT 89.125 1.915 89.54 2.216 ;
      RECT 89.095 1.93 89.54 2.206 ;
      RECT 89.09 1.941 89.54 2.196 ;
      RECT 89.06 1.954 89.54 2.187 ;
      RECT 89.045 1.972 89.54 2.176 ;
      RECT 89.02 1.985 89.54 2.166 ;
      RECT 89.28 1.821 89.29 2.3 ;
      RECT 89.326 1.245 89.365 1.49 ;
      RECT 89.24 1.245 89.375 1.488 ;
      RECT 89.125 1.27 89.375 1.485 ;
      RECT 89.125 1.27 89.38 1.483 ;
      RECT 89.125 1.27 89.395 1.478 ;
      RECT 89.231 1.245 89.41 1.458 ;
      RECT 89.145 1.253 89.41 1.458 ;
      RECT 88.815 0.605 88.985 1.04 ;
      RECT 88.805 0.639 88.985 1.023 ;
      RECT 88.885 0.575 89.055 1.01 ;
      RECT 88.79 0.65 89.055 0.988 ;
      RECT 88.885 0.585 89.06 0.978 ;
      RECT 88.815 0.637 89.09 0.963 ;
      RECT 88.775 0.663 89.09 0.948 ;
      RECT 88.775 0.705 89.1 0.928 ;
      RECT 88.77 0.73 89.105 0.91 ;
      RECT 88.77 0.74 89.11 0.895 ;
      RECT 88.765 0.677 89.09 0.893 ;
      RECT 88.765 0.75 89.115 0.878 ;
      RECT 88.76 0.687 89.09 0.875 ;
      RECT 88.755 0.771 89.12 0.858 ;
      RECT 88.755 0.803 89.125 0.838 ;
      RECT 88.75 0.717 89.1 0.83 ;
      RECT 88.755 0.702 89.09 0.858 ;
      RECT 88.77 0.672 89.09 0.91 ;
      RECT 88.615 1.259 88.84 1.515 ;
      RECT 88.615 1.292 88.86 1.505 ;
      RECT 88.58 1.292 88.86 1.503 ;
      RECT 88.58 1.305 88.865 1.493 ;
      RECT 88.58 1.325 88.875 1.485 ;
      RECT 88.58 1.422 88.88 1.478 ;
      RECT 88.56 1.17 88.69 1.468 ;
      RECT 88.515 1.325 88.875 1.41 ;
      RECT 88.505 1.17 88.69 1.355 ;
      RECT 88.505 1.202 88.776 1.355 ;
      RECT 88.47 1.732 88.49 1.91 ;
      RECT 88.435 1.685 88.47 1.91 ;
      RECT 88.42 1.625 88.435 1.91 ;
      RECT 88.395 1.572 88.42 1.91 ;
      RECT 88.38 1.525 88.395 1.91 ;
      RECT 88.36 1.502 88.38 1.91 ;
      RECT 88.335 1.467 88.36 1.91 ;
      RECT 88.325 1.313 88.335 1.91 ;
      RECT 88.295 1.308 88.325 1.901 ;
      RECT 88.29 1.305 88.295 1.891 ;
      RECT 88.275 1.305 88.29 1.865 ;
      RECT 88.27 1.305 88.275 1.828 ;
      RECT 88.245 1.305 88.27 1.78 ;
      RECT 88.225 1.305 88.245 1.705 ;
      RECT 88.215 1.305 88.225 1.665 ;
      RECT 88.21 1.305 88.215 1.64 ;
      RECT 88.205 1.305 88.21 1.623 ;
      RECT 88.2 1.305 88.205 1.605 ;
      RECT 88.195 1.306 88.2 1.595 ;
      RECT 88.185 1.308 88.195 1.563 ;
      RECT 88.175 1.31 88.185 1.53 ;
      RECT 88.165 1.313 88.175 1.503 ;
      RECT 88.49 1.74 88.715 1.91 ;
      RECT 87.82 0.552 87.99 1.005 ;
      RECT 87.82 0.552 88.08 0.971 ;
      RECT 87.82 0.552 88.11 0.955 ;
      RECT 87.82 0.552 88.14 0.928 ;
      RECT 88.076 0.53 88.155 0.91 ;
      RECT 87.855 0.537 88.16 0.895 ;
      RECT 87.855 0.545 88.17 0.858 ;
      RECT 87.815 0.572 88.17 0.83 ;
      RECT 87.8 0.585 88.17 0.795 ;
      RECT 87.82 0.56 88.19 0.785 ;
      RECT 87.795 0.625 88.19 0.755 ;
      RECT 87.795 0.655 88.195 0.738 ;
      RECT 87.79 0.685 88.195 0.725 ;
      RECT 87.855 0.534 88.155 0.91 ;
      RECT 87.99 0.531 88.076 0.989 ;
      RECT 87.941 0.532 88.155 0.91 ;
      RECT 88.085 2.192 88.13 2.385 ;
      RECT 88.075 2.162 88.085 2.385 ;
      RECT 88.07 2.147 88.075 2.385 ;
      RECT 88.03 2.057 88.07 2.385 ;
      RECT 88.025 1.97 88.03 2.385 ;
      RECT 88.015 1.94 88.025 2.385 ;
      RECT 88.01 1.9 88.015 2.385 ;
      RECT 88 1.862 88.01 2.385 ;
      RECT 87.995 1.827 88 2.385 ;
      RECT 87.975 1.78 87.995 2.385 ;
      RECT 87.96 1.705 87.975 2.385 ;
      RECT 87.955 1.66 87.96 2.38 ;
      RECT 87.95 1.64 87.955 2.353 ;
      RECT 87.945 1.62 87.95 2.338 ;
      RECT 87.94 1.595 87.945 2.318 ;
      RECT 87.935 1.573 87.94 2.303 ;
      RECT 87.93 1.551 87.935 2.285 ;
      RECT 87.925 1.53 87.93 2.275 ;
      RECT 87.915 1.502 87.925 2.245 ;
      RECT 87.905 1.465 87.915 2.213 ;
      RECT 87.895 1.425 87.905 2.18 ;
      RECT 87.885 1.403 87.895 2.15 ;
      RECT 87.855 1.355 87.885 2.082 ;
      RECT 87.84 1.315 87.855 2.009 ;
      RECT 87.83 1.315 87.84 1.975 ;
      RECT 87.825 1.315 87.83 1.95 ;
      RECT 87.82 1.315 87.825 1.935 ;
      RECT 87.815 1.315 87.82 1.913 ;
      RECT 87.81 1.315 87.815 1.9 ;
      RECT 87.795 1.315 87.81 1.865 ;
      RECT 87.775 1.315 87.795 1.805 ;
      RECT 87.765 1.315 87.775 1.755 ;
      RECT 87.745 1.315 87.765 1.703 ;
      RECT 87.725 1.315 87.745 1.66 ;
      RECT 87.715 1.315 87.725 1.648 ;
      RECT 87.685 1.315 87.715 1.635 ;
      RECT 87.655 1.336 87.685 1.615 ;
      RECT 87.645 1.364 87.655 1.595 ;
      RECT 87.63 1.381 87.645 1.563 ;
      RECT 87.625 1.395 87.63 1.53 ;
      RECT 87.62 1.403 87.625 1.503 ;
      RECT 87.615 1.411 87.62 1.465 ;
      RECT 87.62 1.935 87.625 2.27 ;
      RECT 87.585 1.922 87.62 2.269 ;
      RECT 87.515 1.862 87.585 2.268 ;
      RECT 87.435 1.805 87.515 2.267 ;
      RECT 87.3 1.765 87.435 2.266 ;
      RECT 87.3 1.952 87.635 2.255 ;
      RECT 87.26 1.952 87.635 2.245 ;
      RECT 87.26 1.97 87.64 2.24 ;
      RECT 87.26 2.06 87.645 2.23 ;
      RECT 87.255 1.755 87.42 2.21 ;
      RECT 87.25 1.755 87.42 1.953 ;
      RECT 87.25 1.912 87.615 1.953 ;
      RECT 87.25 1.9 87.61 1.953 ;
      RECT 86.515 2.115 87.03 2.525 ;
      RECT 86.69 1.135 87.03 2.525 ;
      RECT 85.8 1.135 87.03 1.305 ;
      RECT 86.51 0.53 86.755 1.305 ;
      RECT 83.91 2.535 85.94 2.705 ;
      RECT 85.77 1.68 85.94 2.705 ;
      RECT 83.91 1.235 84.08 2.705 ;
      RECT 85.77 1.68 86.52 1.87 ;
      RECT 83.885 1.235 84.08 1.565 ;
      RECT 84.59 1.855 85.6 2.025 ;
      RECT 85.41 0.495 85.6 2.025 ;
      RECT 84.59 1.055 84.76 2.025 ;
      RECT 84.25 2.195 85.375 2.365 ;
      RECT 84.25 0.495 84.42 2.365 ;
      RECT 83.405 1.235 83.66 1.565 ;
      RECT 83.49 0.895 83.66 1.565 ;
      RECT 83.49 0.895 84.42 1.065 ;
      RECT 84.245 0.495 84.42 1.065 ;
      RECT 84.245 0.495 84.775 0.86 ;
      RECT 83.065 1.735 83.4 2.705 ;
      RECT 83.065 0.495 83.235 2.705 ;
      RECT 83.065 0.495 83.32 1.065 ;
      RECT 82.315 1.725 82.645 2.705 ;
      RECT 82.415 0.495 82.645 2.705 ;
      RECT 82.315 0.495 82.645 1.125 ;
      RECT 80.935 1.725 81.265 2.705 ;
      RECT 81.035 0.495 81.265 2.705 ;
      RECT 81.035 1.315 82.245 1.555 ;
      RECT 80.935 0.495 81.265 1.125 ;
      RECT 79.555 1.725 79.885 2.705 ;
      RECT 79.655 0.495 79.885 2.705 ;
      RECT 79.555 0.495 79.885 1.125 ;
      RECT 78.175 1.725 78.505 2.705 ;
      RECT 78.275 0.495 78.505 2.705 ;
      RECT 78.275 1.315 79.485 1.555 ;
      RECT 78.175 0.495 78.505 1.125 ;
      RECT 76.855 2.115 77.37 2.525 ;
      RECT 77.03 1.135 77.37 2.525 ;
      RECT 76.14 1.135 77.37 1.305 ;
      RECT 76.85 0.53 77.095 1.305 ;
      RECT 74.25 2.535 76.28 2.705 ;
      RECT 76.11 1.68 76.28 2.705 ;
      RECT 74.25 1.235 74.42 2.705 ;
      RECT 76.11 1.68 76.86 1.87 ;
      RECT 74.225 1.235 74.42 1.565 ;
      RECT 74.93 1.855 75.94 2.025 ;
      RECT 75.75 0.495 75.94 2.025 ;
      RECT 74.93 1.055 75.1 2.025 ;
      RECT 74.59 2.195 75.715 2.365 ;
      RECT 74.59 0.495 74.76 2.365 ;
      RECT 73.745 1.235 74 1.565 ;
      RECT 73.83 0.895 74 1.565 ;
      RECT 73.83 0.895 74.76 1.065 ;
      RECT 74.585 0.495 74.76 1.065 ;
      RECT 74.585 0.495 75.115 0.86 ;
      RECT 73.405 1.735 73.74 2.705 ;
      RECT 73.405 0.495 73.575 2.705 ;
      RECT 73.405 0.495 73.66 1.065 ;
      RECT 72.72 2.115 73.235 2.525 ;
      RECT 72.895 1.135 73.235 2.525 ;
      RECT 72.005 1.135 73.235 1.305 ;
      RECT 72.715 0.53 72.96 1.305 ;
      RECT 70.115 2.535 72.145 2.705 ;
      RECT 71.975 1.68 72.145 2.705 ;
      RECT 70.115 1.235 70.285 2.705 ;
      RECT 71.975 1.68 72.725 1.87 ;
      RECT 70.09 1.235 70.285 1.565 ;
      RECT 70.795 1.855 71.805 2.025 ;
      RECT 71.615 0.495 71.805 2.025 ;
      RECT 70.795 1.055 70.965 2.025 ;
      RECT 70.455 2.195 71.58 2.365 ;
      RECT 70.455 0.495 70.625 2.365 ;
      RECT 69.61 1.235 69.865 1.565 ;
      RECT 69.695 0.895 69.865 1.565 ;
      RECT 69.695 0.895 70.625 1.065 ;
      RECT 70.45 0.495 70.625 1.065 ;
      RECT 70.45 0.495 70.98 0.86 ;
      RECT 69.27 1.735 69.605 2.705 ;
      RECT 69.27 0.495 69.44 2.705 ;
      RECT 69.27 0.495 69.525 1.065 ;
      RECT 68.175 0.715 68.905 0.955 ;
      RECT 68.717 0.51 68.905 0.955 ;
      RECT 68.545 0.522 68.92 0.949 ;
      RECT 68.46 0.537 68.94 0.934 ;
      RECT 68.46 0.552 68.945 0.924 ;
      RECT 68.415 0.572 68.96 0.916 ;
      RECT 68.392 0.607 68.975 0.87 ;
      RECT 68.306 0.63 68.98 0.83 ;
      RECT 68.306 0.648 68.99 0.8 ;
      RECT 68.175 0.717 68.995 0.763 ;
      RECT 68.22 0.66 68.99 0.8 ;
      RECT 68.306 0.612 68.975 0.87 ;
      RECT 68.392 0.581 68.96 0.916 ;
      RECT 68.415 0.562 68.945 0.924 ;
      RECT 68.46 0.535 68.92 0.949 ;
      RECT 68.545 0.517 68.905 0.955 ;
      RECT 68.631 0.511 68.905 0.955 ;
      RECT 68.717 0.506 68.85 0.955 ;
      RECT 68.803 0.501 68.85 0.955 ;
      RECT 68.495 1.399 68.665 1.785 ;
      RECT 68.49 1.399 68.665 1.78 ;
      RECT 68.465 1.399 68.665 1.745 ;
      RECT 68.465 1.427 68.675 1.735 ;
      RECT 68.445 1.427 68.675 1.695 ;
      RECT 68.44 1.427 68.675 1.668 ;
      RECT 68.44 1.445 68.68 1.66 ;
      RECT 68.385 1.445 68.68 1.595 ;
      RECT 68.385 1.462 68.69 1.578 ;
      RECT 68.375 1.462 68.69 1.518 ;
      RECT 68.375 1.479 68.695 1.515 ;
      RECT 68.37 1.315 68.54 1.493 ;
      RECT 68.37 1.349 68.626 1.493 ;
      RECT 68.365 2.115 68.37 2.128 ;
      RECT 68.36 2.01 68.365 2.133 ;
      RECT 68.335 1.87 68.36 2.148 ;
      RECT 68.3 1.821 68.335 2.18 ;
      RECT 68.295 1.789 68.3 2.2 ;
      RECT 68.29 1.78 68.295 2.2 ;
      RECT 68.21 1.745 68.29 2.2 ;
      RECT 68.147 1.715 68.21 2.2 ;
      RECT 68.061 1.703 68.147 2.2 ;
      RECT 67.975 1.689 68.061 2.2 ;
      RECT 67.895 1.676 67.975 2.186 ;
      RECT 67.86 1.668 67.895 2.166 ;
      RECT 67.85 1.665 67.86 2.157 ;
      RECT 67.82 1.66 67.85 2.144 ;
      RECT 67.77 1.635 67.82 2.12 ;
      RECT 67.756 1.609 67.77 2.102 ;
      RECT 67.67 1.569 67.756 2.078 ;
      RECT 67.625 1.517 67.67 2.047 ;
      RECT 67.615 1.492 67.625 2.034 ;
      RECT 67.61 1.273 67.615 1.295 ;
      RECT 67.605 1.475 67.615 2.03 ;
      RECT 67.605 1.271 67.61 1.385 ;
      RECT 67.595 1.267 67.605 2.026 ;
      RECT 67.551 1.265 67.595 2.014 ;
      RECT 67.465 1.265 67.551 1.985 ;
      RECT 67.435 1.265 67.465 1.958 ;
      RECT 67.42 1.265 67.435 1.946 ;
      RECT 67.38 1.277 67.42 1.931 ;
      RECT 67.36 1.296 67.38 1.91 ;
      RECT 67.35 1.306 67.36 1.894 ;
      RECT 67.34 1.312 67.35 1.883 ;
      RECT 67.32 1.322 67.34 1.866 ;
      RECT 67.315 1.331 67.32 1.853 ;
      RECT 67.31 1.335 67.315 1.803 ;
      RECT 67.3 1.341 67.31 1.72 ;
      RECT 67.295 1.345 67.3 1.634 ;
      RECT 67.29 1.365 67.295 1.571 ;
      RECT 67.285 1.388 67.29 1.518 ;
      RECT 67.28 1.406 67.285 1.463 ;
      RECT 67.89 1.225 68.06 1.485 ;
      RECT 68.06 1.19 68.105 1.471 ;
      RECT 68.021 1.192 68.11 1.454 ;
      RECT 67.91 1.209 68.196 1.425 ;
      RECT 67.91 1.224 68.2 1.397 ;
      RECT 67.91 1.205 68.11 1.454 ;
      RECT 67.935 1.193 68.06 1.485 ;
      RECT 68.021 1.191 68.105 1.471 ;
      RECT 67.075 0.58 67.245 1.07 ;
      RECT 67.075 0.58 67.28 1.05 ;
      RECT 67.21 0.5 67.32 1.01 ;
      RECT 67.191 0.504 67.34 0.98 ;
      RECT 67.105 0.512 67.36 0.963 ;
      RECT 67.105 0.518 67.365 0.953 ;
      RECT 67.105 0.527 67.385 0.941 ;
      RECT 67.08 0.552 67.415 0.919 ;
      RECT 67.08 0.572 67.42 0.899 ;
      RECT 67.075 0.585 67.43 0.879 ;
      RECT 67.075 0.652 67.435 0.86 ;
      RECT 67.075 0.785 67.44 0.847 ;
      RECT 67.07 0.59 67.43 0.68 ;
      RECT 67.08 0.547 67.385 0.941 ;
      RECT 67.191 0.502 67.32 1.01 ;
      RECT 67.065 2.255 67.365 2.51 ;
      RECT 67.15 2.221 67.365 2.51 ;
      RECT 67.15 2.224 67.37 2.37 ;
      RECT 67.085 2.245 67.37 2.37 ;
      RECT 67.12 2.235 67.365 2.51 ;
      RECT 67.115 2.24 67.37 2.37 ;
      RECT 67.15 2.219 67.351 2.51 ;
      RECT 67.236 2.21 67.351 2.51 ;
      RECT 67.236 2.204 67.265 2.51 ;
      RECT 66.725 1.845 66.735 2.335 ;
      RECT 66.385 1.78 66.395 2.08 ;
      RECT 66.9 1.952 66.905 2.171 ;
      RECT 66.89 1.932 66.9 2.188 ;
      RECT 66.88 1.912 66.89 2.218 ;
      RECT 66.875 1.902 66.88 2.233 ;
      RECT 66.87 1.898 66.875 2.238 ;
      RECT 66.855 1.89 66.87 2.245 ;
      RECT 66.815 1.87 66.855 2.27 ;
      RECT 66.79 1.852 66.815 2.303 ;
      RECT 66.785 1.85 66.79 2.316 ;
      RECT 66.765 1.847 66.785 2.32 ;
      RECT 66.735 1.845 66.765 2.33 ;
      RECT 66.665 1.847 66.725 2.331 ;
      RECT 66.645 1.847 66.665 2.325 ;
      RECT 66.62 1.845 66.645 2.322 ;
      RECT 66.585 1.84 66.62 2.318 ;
      RECT 66.565 1.834 66.585 2.305 ;
      RECT 66.555 1.831 66.565 2.293 ;
      RECT 66.535 1.828 66.555 2.278 ;
      RECT 66.515 1.824 66.535 2.26 ;
      RECT 66.51 1.821 66.515 2.25 ;
      RECT 66.505 1.82 66.51 2.248 ;
      RECT 66.495 1.817 66.505 2.24 ;
      RECT 66.485 1.811 66.495 2.223 ;
      RECT 66.475 1.805 66.485 2.205 ;
      RECT 66.465 1.799 66.475 2.193 ;
      RECT 66.455 1.793 66.465 2.173 ;
      RECT 66.45 1.789 66.455 2.158 ;
      RECT 66.445 1.787 66.45 2.15 ;
      RECT 66.44 1.785 66.445 2.143 ;
      RECT 66.435 1.783 66.44 2.133 ;
      RECT 66.43 1.781 66.435 2.127 ;
      RECT 66.42 1.78 66.43 2.117 ;
      RECT 66.41 1.78 66.42 2.108 ;
      RECT 66.395 1.78 66.41 2.093 ;
      RECT 66.355 1.78 66.385 2.077 ;
      RECT 66.335 1.782 66.355 2.072 ;
      RECT 66.33 1.787 66.335 2.07 ;
      RECT 66.3 1.795 66.33 2.068 ;
      RECT 66.27 1.81 66.3 2.067 ;
      RECT 66.225 1.832 66.27 2.072 ;
      RECT 66.22 1.847 66.225 2.076 ;
      RECT 66.205 1.852 66.22 2.078 ;
      RECT 66.2 1.856 66.205 2.08 ;
      RECT 66.14 1.879 66.2 2.089 ;
      RECT 66.12 1.905 66.14 2.102 ;
      RECT 66.11 1.912 66.12 2.106 ;
      RECT 66.095 1.919 66.11 2.109 ;
      RECT 66.075 1.929 66.095 2.112 ;
      RECT 66.07 1.937 66.075 2.115 ;
      RECT 66.025 1.942 66.07 2.122 ;
      RECT 66.015 1.945 66.025 2.129 ;
      RECT 66.005 1.945 66.015 2.133 ;
      RECT 65.97 1.947 66.005 2.145 ;
      RECT 65.95 1.95 65.97 2.158 ;
      RECT 65.91 1.953 65.95 2.169 ;
      RECT 65.895 1.955 65.91 2.182 ;
      RECT 65.885 1.955 65.895 2.187 ;
      RECT 65.86 1.956 65.885 2.195 ;
      RECT 65.85 1.958 65.86 2.2 ;
      RECT 65.845 1.959 65.85 2.203 ;
      RECT 65.82 1.957 65.845 2.206 ;
      RECT 65.805 1.955 65.82 2.207 ;
      RECT 65.785 1.952 65.805 2.209 ;
      RECT 65.765 1.947 65.785 2.209 ;
      RECT 65.705 1.942 65.765 2.206 ;
      RECT 65.67 1.917 65.705 2.202 ;
      RECT 65.66 1.894 65.67 2.2 ;
      RECT 65.63 1.871 65.66 2.2 ;
      RECT 65.62 1.85 65.63 2.2 ;
      RECT 65.595 1.832 65.62 2.198 ;
      RECT 65.58 1.81 65.595 2.195 ;
      RECT 65.565 1.792 65.58 2.193 ;
      RECT 65.545 1.782 65.565 2.191 ;
      RECT 65.53 1.777 65.545 2.19 ;
      RECT 65.515 1.775 65.53 2.189 ;
      RECT 65.485 1.776 65.515 2.187 ;
      RECT 65.465 1.779 65.485 2.185 ;
      RECT 65.408 1.783 65.465 2.185 ;
      RECT 65.322 1.792 65.408 2.185 ;
      RECT 65.236 1.803 65.322 2.185 ;
      RECT 65.15 1.814 65.236 2.185 ;
      RECT 65.13 1.821 65.15 2.193 ;
      RECT 65.12 1.824 65.13 2.2 ;
      RECT 65.055 1.829 65.12 2.218 ;
      RECT 65.025 1.836 65.055 2.243 ;
      RECT 65.015 1.839 65.025 2.25 ;
      RECT 64.97 1.843 65.015 2.255 ;
      RECT 64.94 1.848 64.97 2.26 ;
      RECT 64.939 1.85 64.94 2.26 ;
      RECT 64.853 1.856 64.939 2.26 ;
      RECT 64.767 1.867 64.853 2.26 ;
      RECT 64.681 1.879 64.767 2.26 ;
      RECT 64.595 1.89 64.681 2.26 ;
      RECT 64.58 1.897 64.595 2.255 ;
      RECT 64.575 1.899 64.58 2.249 ;
      RECT 64.555 1.91 64.575 2.244 ;
      RECT 64.545 1.928 64.555 2.238 ;
      RECT 64.54 1.94 64.545 2.038 ;
      RECT 66.835 0.693 66.855 0.78 ;
      RECT 66.83 0.628 66.835 0.812 ;
      RECT 66.82 0.595 66.83 0.817 ;
      RECT 66.815 0.575 66.82 0.823 ;
      RECT 66.785 0.575 66.815 0.84 ;
      RECT 66.736 0.575 66.785 0.876 ;
      RECT 66.65 0.575 66.736 0.934 ;
      RECT 66.621 0.585 66.65 0.983 ;
      RECT 66.535 0.627 66.621 1.036 ;
      RECT 66.515 0.665 66.535 1.083 ;
      RECT 66.49 0.682 66.515 1.103 ;
      RECT 66.48 0.696 66.49 1.123 ;
      RECT 66.475 0.702 66.48 1.133 ;
      RECT 66.47 0.706 66.475 1.14 ;
      RECT 66.42 0.726 66.47 1.145 ;
      RECT 66.355 0.77 66.42 1.145 ;
      RECT 66.33 0.82 66.355 1.145 ;
      RECT 66.32 0.85 66.33 1.145 ;
      RECT 66.315 0.877 66.32 1.145 ;
      RECT 66.31 0.895 66.315 1.145 ;
      RECT 66.3 0.937 66.31 1.145 ;
      RECT 66.65 1.495 66.82 1.67 ;
      RECT 66.59 1.323 66.65 1.658 ;
      RECT 66.58 1.316 66.59 1.641 ;
      RECT 66.535 1.495 66.82 1.621 ;
      RECT 66.516 1.495 66.82 1.599 ;
      RECT 66.43 1.495 66.82 1.564 ;
      RECT 66.41 1.315 66.58 1.52 ;
      RECT 66.41 1.462 66.815 1.52 ;
      RECT 66.41 1.41 66.79 1.52 ;
      RECT 66.41 1.365 66.755 1.52 ;
      RECT 66.41 1.347 66.72 1.52 ;
      RECT 66.41 1.337 66.715 1.52 ;
      RECT 66.13 2.295 66.32 2.52 ;
      RECT 66.12 2.296 66.325 2.515 ;
      RECT 66.12 2.298 66.335 2.495 ;
      RECT 66.12 2.302 66.34 2.48 ;
      RECT 66.12 2.289 66.29 2.515 ;
      RECT 66.12 2.292 66.315 2.515 ;
      RECT 66.13 2.288 66.29 2.52 ;
      RECT 66.216 2.286 66.29 2.52 ;
      RECT 65.84 1.537 66.01 1.775 ;
      RECT 65.84 1.537 66.096 1.689 ;
      RECT 65.84 1.537 66.1 1.599 ;
      RECT 65.89 1.31 66.11 1.578 ;
      RECT 65.885 1.327 66.115 1.551 ;
      RECT 65.85 1.485 66.115 1.551 ;
      RECT 65.87 1.335 66.01 1.775 ;
      RECT 65.86 1.417 66.12 1.534 ;
      RECT 65.855 1.465 66.12 1.534 ;
      RECT 65.86 1.375 66.115 1.551 ;
      RECT 65.885 1.312 66.11 1.578 ;
      RECT 65.45 1.287 65.62 1.485 ;
      RECT 65.45 1.287 65.665 1.46 ;
      RECT 65.52 1.23 65.69 1.418 ;
      RECT 65.495 1.245 65.69 1.418 ;
      RECT 65.11 1.291 65.14 1.485 ;
      RECT 65.105 1.263 65.11 1.485 ;
      RECT 65.075 1.237 65.105 1.487 ;
      RECT 65.05 1.195 65.075 1.49 ;
      RECT 65.04 1.167 65.05 1.492 ;
      RECT 65.005 1.147 65.04 1.494 ;
      RECT 64.94 1.132 65.005 1.5 ;
      RECT 64.89 1.13 64.94 1.506 ;
      RECT 64.867 1.132 64.89 1.511 ;
      RECT 64.781 1.143 64.867 1.517 ;
      RECT 64.695 1.161 64.781 1.527 ;
      RECT 64.68 1.172 64.695 1.533 ;
      RECT 64.61 1.195 64.68 1.539 ;
      RECT 64.555 1.227 64.61 1.547 ;
      RECT 64.515 1.25 64.555 1.553 ;
      RECT 64.501 1.263 64.515 1.556 ;
      RECT 64.415 1.285 64.501 1.562 ;
      RECT 64.4 1.31 64.415 1.568 ;
      RECT 64.36 1.325 64.4 1.572 ;
      RECT 64.31 1.34 64.36 1.577 ;
      RECT 64.285 1.347 64.31 1.581 ;
      RECT 64.225 1.342 64.285 1.585 ;
      RECT 64.21 1.333 64.225 1.589 ;
      RECT 64.14 1.323 64.21 1.585 ;
      RECT 64.115 1.315 64.135 1.575 ;
      RECT 64.056 1.315 64.115 1.553 ;
      RECT 63.97 1.315 64.056 1.51 ;
      RECT 64.135 1.315 64.14 1.58 ;
      RECT 64.83 0.546 65 0.88 ;
      RECT 64.8 0.546 65 0.875 ;
      RECT 64.74 0.513 64.8 0.863 ;
      RECT 64.74 0.569 65.01 0.858 ;
      RECT 64.715 0.569 65.01 0.852 ;
      RECT 64.71 0.51 64.74 0.849 ;
      RECT 64.695 0.516 64.83 0.847 ;
      RECT 64.69 0.524 64.915 0.835 ;
      RECT 64.69 0.576 65.025 0.788 ;
      RECT 64.675 0.532 64.915 0.783 ;
      RECT 64.675 0.602 65.035 0.724 ;
      RECT 64.645 0.552 65 0.685 ;
      RECT 64.645 0.642 65.045 0.681 ;
      RECT 64.695 0.521 64.915 0.847 ;
      RECT 64.035 0.851 64.09 1.115 ;
      RECT 64.035 0.851 64.155 1.114 ;
      RECT 64.035 0.851 64.18 1.113 ;
      RECT 64.035 0.851 64.245 1.112 ;
      RECT 64.18 0.817 64.26 1.111 ;
      RECT 63.995 0.861 64.405 1.11 ;
      RECT 64.035 0.858 64.405 1.11 ;
      RECT 63.995 0.866 64.41 1.103 ;
      RECT 63.98 0.868 64.41 1.102 ;
      RECT 63.98 0.875 64.415 1.098 ;
      RECT 63.96 0.874 64.41 1.094 ;
      RECT 63.96 0.882 64.42 1.093 ;
      RECT 63.955 0.879 64.415 1.089 ;
      RECT 63.955 0.892 64.43 1.088 ;
      RECT 63.94 0.882 64.42 1.087 ;
      RECT 63.905 0.895 64.43 1.08 ;
      RECT 64.09 0.85 64.4 1.11 ;
      RECT 64.09 0.835 64.35 1.11 ;
      RECT 64.155 0.822 64.285 1.11 ;
      RECT 63.7 1.911 63.715 2.304 ;
      RECT 63.665 1.916 63.715 2.303 ;
      RECT 63.7 1.915 63.76 2.302 ;
      RECT 63.645 1.926 63.76 2.301 ;
      RECT 63.66 1.922 63.76 2.301 ;
      RECT 63.625 1.932 63.835 2.298 ;
      RECT 63.625 1.951 63.88 2.296 ;
      RECT 63.625 1.958 63.885 2.293 ;
      RECT 63.61 1.935 63.835 2.29 ;
      RECT 63.59 1.94 63.835 2.283 ;
      RECT 63.585 1.944 63.835 2.279 ;
      RECT 63.585 1.961 63.895 2.278 ;
      RECT 63.565 1.955 63.88 2.274 ;
      RECT 63.565 1.964 63.9 2.268 ;
      RECT 63.56 1.97 63.9 2.04 ;
      RECT 63.625 1.93 63.76 2.298 ;
      RECT 63.5 1.293 63.7 1.605 ;
      RECT 63.575 1.271 63.7 1.605 ;
      RECT 63.515 1.29 63.705 1.59 ;
      RECT 63.485 1.301 63.705 1.588 ;
      RECT 63.5 1.296 63.71 1.554 ;
      RECT 63.485 1.4 63.715 1.521 ;
      RECT 63.515 1.272 63.7 1.605 ;
      RECT 63.575 1.25 63.675 1.605 ;
      RECT 63.6 1.247 63.675 1.605 ;
      RECT 63.6 1.242 63.62 1.605 ;
      RECT 63.005 1.31 63.18 1.485 ;
      RECT 63 1.31 63.18 1.483 ;
      RECT 62.975 1.31 63.18 1.478 ;
      RECT 62.92 1.29 63.09 1.468 ;
      RECT 62.92 1.297 63.155 1.468 ;
      RECT 63.005 1.977 63.02 2.16 ;
      RECT 62.995 1.955 63.005 2.16 ;
      RECT 62.98 1.935 62.995 2.16 ;
      RECT 62.97 1.91 62.98 2.16 ;
      RECT 62.94 1.875 62.97 2.16 ;
      RECT 62.905 1.815 62.94 2.16 ;
      RECT 62.9 1.777 62.905 2.16 ;
      RECT 62.85 1.728 62.9 2.16 ;
      RECT 62.84 1.678 62.85 2.148 ;
      RECT 62.825 1.657 62.84 2.108 ;
      RECT 62.805 1.625 62.825 2.058 ;
      RECT 62.78 1.581 62.805 1.998 ;
      RECT 62.775 1.553 62.78 1.953 ;
      RECT 62.77 1.544 62.775 1.939 ;
      RECT 62.765 1.537 62.77 1.926 ;
      RECT 62.76 1.532 62.765 1.915 ;
      RECT 62.755 1.517 62.76 1.905 ;
      RECT 62.75 1.495 62.755 1.892 ;
      RECT 62.74 1.455 62.75 1.867 ;
      RECT 62.715 1.385 62.74 1.823 ;
      RECT 62.71 1.325 62.715 1.788 ;
      RECT 62.695 1.305 62.71 1.755 ;
      RECT 62.69 1.305 62.695 1.73 ;
      RECT 62.66 1.305 62.69 1.685 ;
      RECT 62.615 1.305 62.66 1.625 ;
      RECT 62.54 1.305 62.615 1.573 ;
      RECT 62.535 1.305 62.54 1.538 ;
      RECT 62.53 1.305 62.535 1.528 ;
      RECT 62.525 1.305 62.53 1.508 ;
      RECT 62.79 0.525 62.96 0.995 ;
      RECT 62.735 0.518 62.93 0.979 ;
      RECT 62.735 0.532 62.965 0.978 ;
      RECT 62.72 0.533 62.965 0.959 ;
      RECT 62.715 0.551 62.965 0.945 ;
      RECT 62.72 0.534 62.97 0.943 ;
      RECT 62.705 0.565 62.97 0.928 ;
      RECT 62.72 0.54 62.975 0.913 ;
      RECT 62.7 0.58 62.975 0.91 ;
      RECT 62.715 0.552 62.98 0.895 ;
      RECT 62.715 0.564 62.985 0.875 ;
      RECT 62.7 0.58 62.99 0.858 ;
      RECT 62.7 0.59 62.995 0.713 ;
      RECT 62.695 0.59 62.995 0.67 ;
      RECT 62.695 0.605 63 0.648 ;
      RECT 62.79 0.515 62.93 0.995 ;
      RECT 62.79 0.513 62.9 0.995 ;
      RECT 62.876 0.51 62.9 0.995 ;
      RECT 62.535 2.177 62.54 2.223 ;
      RECT 62.525 2.025 62.535 2.247 ;
      RECT 62.52 1.87 62.525 2.272 ;
      RECT 62.505 1.832 62.52 2.283 ;
      RECT 62.5 1.815 62.505 2.29 ;
      RECT 62.49 1.803 62.5 2.297 ;
      RECT 62.485 1.794 62.49 2.299 ;
      RECT 62.48 1.792 62.485 2.303 ;
      RECT 62.435 1.783 62.48 2.318 ;
      RECT 62.43 1.775 62.435 2.332 ;
      RECT 62.425 1.772 62.43 2.336 ;
      RECT 62.41 1.767 62.425 2.344 ;
      RECT 62.355 1.757 62.41 2.355 ;
      RECT 62.32 1.745 62.355 2.356 ;
      RECT 62.311 1.74 62.32 2.35 ;
      RECT 62.225 1.74 62.311 2.34 ;
      RECT 62.195 1.74 62.225 2.318 ;
      RECT 62.185 1.74 62.19 2.298 ;
      RECT 62.18 1.74 62.185 2.26 ;
      RECT 62.175 1.74 62.18 2.218 ;
      RECT 62.17 1.74 62.175 2.178 ;
      RECT 62.165 1.74 62.17 2.108 ;
      RECT 62.155 1.74 62.165 2.03 ;
      RECT 62.15 1.74 62.155 1.93 ;
      RECT 62.19 1.74 62.195 2.3 ;
      RECT 61.685 1.822 61.775 2.3 ;
      RECT 61.67 1.825 61.79 2.298 ;
      RECT 61.685 1.824 61.79 2.298 ;
      RECT 61.65 1.831 61.815 2.288 ;
      RECT 61.67 1.825 61.815 2.288 ;
      RECT 61.635 1.837 61.815 2.276 ;
      RECT 61.67 1.828 61.865 2.269 ;
      RECT 61.621 1.845 61.865 2.267 ;
      RECT 61.65 1.835 61.875 2.255 ;
      RECT 61.621 1.856 61.905 2.246 ;
      RECT 61.535 1.88 61.905 2.24 ;
      RECT 61.535 1.893 61.945 2.223 ;
      RECT 61.53 1.915 61.945 2.216 ;
      RECT 61.5 1.93 61.945 2.206 ;
      RECT 61.495 1.941 61.945 2.196 ;
      RECT 61.465 1.954 61.945 2.187 ;
      RECT 61.45 1.972 61.945 2.176 ;
      RECT 61.425 1.985 61.945 2.166 ;
      RECT 61.685 1.821 61.695 2.3 ;
      RECT 61.731 1.245 61.77 1.49 ;
      RECT 61.645 1.245 61.78 1.488 ;
      RECT 61.53 1.27 61.78 1.485 ;
      RECT 61.53 1.27 61.785 1.483 ;
      RECT 61.53 1.27 61.8 1.478 ;
      RECT 61.636 1.245 61.815 1.458 ;
      RECT 61.55 1.253 61.815 1.458 ;
      RECT 61.22 0.605 61.39 1.04 ;
      RECT 61.21 0.639 61.39 1.023 ;
      RECT 61.29 0.575 61.46 1.01 ;
      RECT 61.195 0.65 61.46 0.988 ;
      RECT 61.29 0.585 61.465 0.978 ;
      RECT 61.22 0.637 61.495 0.963 ;
      RECT 61.18 0.663 61.495 0.948 ;
      RECT 61.18 0.705 61.505 0.928 ;
      RECT 61.175 0.73 61.51 0.91 ;
      RECT 61.175 0.74 61.515 0.895 ;
      RECT 61.17 0.677 61.495 0.893 ;
      RECT 61.17 0.75 61.52 0.878 ;
      RECT 61.165 0.687 61.495 0.875 ;
      RECT 61.16 0.771 61.525 0.858 ;
      RECT 61.16 0.803 61.53 0.838 ;
      RECT 61.155 0.717 61.505 0.83 ;
      RECT 61.16 0.702 61.495 0.858 ;
      RECT 61.175 0.672 61.495 0.91 ;
      RECT 61.02 1.259 61.245 1.515 ;
      RECT 61.02 1.292 61.265 1.505 ;
      RECT 60.985 1.292 61.265 1.503 ;
      RECT 60.985 1.305 61.27 1.493 ;
      RECT 60.985 1.325 61.28 1.485 ;
      RECT 60.985 1.422 61.285 1.478 ;
      RECT 60.965 1.17 61.095 1.468 ;
      RECT 60.92 1.325 61.28 1.41 ;
      RECT 60.91 1.17 61.095 1.355 ;
      RECT 60.91 1.202 61.181 1.355 ;
      RECT 60.875 1.732 60.895 1.91 ;
      RECT 60.84 1.685 60.875 1.91 ;
      RECT 60.825 1.625 60.84 1.91 ;
      RECT 60.8 1.572 60.825 1.91 ;
      RECT 60.785 1.525 60.8 1.91 ;
      RECT 60.765 1.502 60.785 1.91 ;
      RECT 60.74 1.467 60.765 1.91 ;
      RECT 60.73 1.313 60.74 1.91 ;
      RECT 60.7 1.308 60.73 1.901 ;
      RECT 60.695 1.305 60.7 1.891 ;
      RECT 60.68 1.305 60.695 1.865 ;
      RECT 60.675 1.305 60.68 1.828 ;
      RECT 60.65 1.305 60.675 1.78 ;
      RECT 60.63 1.305 60.65 1.705 ;
      RECT 60.62 1.305 60.63 1.665 ;
      RECT 60.615 1.305 60.62 1.64 ;
      RECT 60.61 1.305 60.615 1.623 ;
      RECT 60.605 1.305 60.61 1.605 ;
      RECT 60.6 1.306 60.605 1.595 ;
      RECT 60.59 1.308 60.6 1.563 ;
      RECT 60.58 1.31 60.59 1.53 ;
      RECT 60.57 1.313 60.58 1.503 ;
      RECT 60.895 1.74 61.12 1.91 ;
      RECT 60.225 0.552 60.395 1.005 ;
      RECT 60.225 0.552 60.485 0.971 ;
      RECT 60.225 0.552 60.515 0.955 ;
      RECT 60.225 0.552 60.545 0.928 ;
      RECT 60.481 0.53 60.56 0.91 ;
      RECT 60.26 0.537 60.565 0.895 ;
      RECT 60.26 0.545 60.575 0.858 ;
      RECT 60.22 0.572 60.575 0.83 ;
      RECT 60.205 0.585 60.575 0.795 ;
      RECT 60.225 0.56 60.595 0.785 ;
      RECT 60.2 0.625 60.595 0.755 ;
      RECT 60.2 0.655 60.6 0.738 ;
      RECT 60.195 0.685 60.6 0.725 ;
      RECT 60.26 0.534 60.56 0.91 ;
      RECT 60.395 0.531 60.481 0.989 ;
      RECT 60.346 0.532 60.56 0.91 ;
      RECT 60.49 2.192 60.535 2.385 ;
      RECT 60.48 2.162 60.49 2.385 ;
      RECT 60.475 2.147 60.48 2.385 ;
      RECT 60.435 2.057 60.475 2.385 ;
      RECT 60.43 1.97 60.435 2.385 ;
      RECT 60.42 1.94 60.43 2.385 ;
      RECT 60.415 1.9 60.42 2.385 ;
      RECT 60.405 1.862 60.415 2.385 ;
      RECT 60.4 1.827 60.405 2.385 ;
      RECT 60.38 1.78 60.4 2.385 ;
      RECT 60.365 1.705 60.38 2.385 ;
      RECT 60.36 1.66 60.365 2.38 ;
      RECT 60.355 1.64 60.36 2.353 ;
      RECT 60.35 1.62 60.355 2.338 ;
      RECT 60.345 1.595 60.35 2.318 ;
      RECT 60.34 1.573 60.345 2.303 ;
      RECT 60.335 1.551 60.34 2.285 ;
      RECT 60.33 1.53 60.335 2.275 ;
      RECT 60.32 1.502 60.33 2.245 ;
      RECT 60.31 1.465 60.32 2.213 ;
      RECT 60.3 1.425 60.31 2.18 ;
      RECT 60.29 1.403 60.3 2.15 ;
      RECT 60.26 1.355 60.29 2.082 ;
      RECT 60.245 1.315 60.26 2.009 ;
      RECT 60.235 1.315 60.245 1.975 ;
      RECT 60.23 1.315 60.235 1.95 ;
      RECT 60.225 1.315 60.23 1.935 ;
      RECT 60.22 1.315 60.225 1.913 ;
      RECT 60.215 1.315 60.22 1.9 ;
      RECT 60.2 1.315 60.215 1.865 ;
      RECT 60.18 1.315 60.2 1.805 ;
      RECT 60.17 1.315 60.18 1.755 ;
      RECT 60.15 1.315 60.17 1.703 ;
      RECT 60.13 1.315 60.15 1.66 ;
      RECT 60.12 1.315 60.13 1.648 ;
      RECT 60.09 1.315 60.12 1.635 ;
      RECT 60.06 1.336 60.09 1.615 ;
      RECT 60.05 1.364 60.06 1.595 ;
      RECT 60.035 1.381 60.05 1.563 ;
      RECT 60.03 1.395 60.035 1.53 ;
      RECT 60.025 1.403 60.03 1.503 ;
      RECT 60.02 1.411 60.025 1.465 ;
      RECT 60.025 1.935 60.03 2.27 ;
      RECT 59.99 1.922 60.025 2.269 ;
      RECT 59.92 1.862 59.99 2.268 ;
      RECT 59.84 1.805 59.92 2.267 ;
      RECT 59.705 1.765 59.84 2.266 ;
      RECT 59.705 1.952 60.04 2.255 ;
      RECT 59.665 1.952 60.04 2.245 ;
      RECT 59.665 1.97 60.045 2.24 ;
      RECT 59.665 2.06 60.05 2.23 ;
      RECT 59.66 1.755 59.825 2.21 ;
      RECT 59.655 1.755 59.825 1.953 ;
      RECT 59.655 1.912 60.02 1.953 ;
      RECT 59.655 1.9 60.015 1.953 ;
      RECT 58.92 2.115 59.435 2.525 ;
      RECT 59.095 1.135 59.435 2.525 ;
      RECT 58.205 1.135 59.435 1.305 ;
      RECT 58.915 0.53 59.16 1.305 ;
      RECT 56.315 2.535 58.345 2.705 ;
      RECT 58.175 1.68 58.345 2.705 ;
      RECT 56.315 1.235 56.485 2.705 ;
      RECT 58.175 1.68 58.925 1.87 ;
      RECT 56.29 1.235 56.485 1.565 ;
      RECT 56.995 1.855 58.005 2.025 ;
      RECT 57.815 0.495 58.005 2.025 ;
      RECT 56.995 1.055 57.165 2.025 ;
      RECT 56.655 2.195 57.78 2.365 ;
      RECT 56.655 0.495 56.825 2.365 ;
      RECT 55.81 1.235 56.065 1.565 ;
      RECT 55.895 0.895 56.065 1.565 ;
      RECT 55.895 0.895 56.825 1.065 ;
      RECT 56.65 0.495 56.825 1.065 ;
      RECT 56.65 0.495 57.18 0.86 ;
      RECT 55.47 1.735 55.805 2.705 ;
      RECT 55.47 0.495 55.64 2.705 ;
      RECT 55.47 0.495 55.725 1.065 ;
      RECT 54.72 1.725 55.05 2.705 ;
      RECT 54.82 0.495 55.05 2.705 ;
      RECT 54.72 0.495 55.05 1.125 ;
      RECT 53.34 1.725 53.67 2.705 ;
      RECT 53.44 0.495 53.67 2.705 ;
      RECT 53.44 1.315 54.65 1.555 ;
      RECT 53.34 0.495 53.67 1.125 ;
      RECT 51.96 1.725 52.29 2.705 ;
      RECT 52.06 0.495 52.29 2.705 ;
      RECT 51.96 0.495 52.29 1.125 ;
      RECT 50.58 1.725 50.91 2.705 ;
      RECT 50.68 0.495 50.91 2.705 ;
      RECT 50.68 1.315 51.89 1.555 ;
      RECT 50.58 0.495 50.91 1.125 ;
      RECT 49.26 2.115 49.775 2.525 ;
      RECT 49.435 1.135 49.775 2.525 ;
      RECT 48.545 1.135 49.775 1.305 ;
      RECT 49.255 0.53 49.5 1.305 ;
      RECT 46.655 2.535 48.685 2.705 ;
      RECT 48.515 1.68 48.685 2.705 ;
      RECT 46.655 1.235 46.825 2.705 ;
      RECT 48.515 1.68 49.265 1.87 ;
      RECT 46.63 1.235 46.825 1.565 ;
      RECT 47.335 1.855 48.345 2.025 ;
      RECT 48.155 0.495 48.345 2.025 ;
      RECT 47.335 1.055 47.505 2.025 ;
      RECT 46.995 2.195 48.12 2.365 ;
      RECT 46.995 0.495 47.165 2.365 ;
      RECT 46.15 1.235 46.405 1.565 ;
      RECT 46.235 0.895 46.405 1.565 ;
      RECT 46.235 0.895 47.165 1.065 ;
      RECT 46.99 0.495 47.165 1.065 ;
      RECT 46.99 0.495 47.52 0.86 ;
      RECT 45.81 1.735 46.145 2.705 ;
      RECT 45.81 0.495 45.98 2.705 ;
      RECT 45.81 0.495 46.065 1.065 ;
      RECT 45.125 2.115 45.64 2.525 ;
      RECT 45.3 1.135 45.64 2.525 ;
      RECT 44.41 1.135 45.64 1.305 ;
      RECT 45.12 0.53 45.365 1.305 ;
      RECT 42.52 2.535 44.55 2.705 ;
      RECT 44.38 1.68 44.55 2.705 ;
      RECT 42.52 1.235 42.69 2.705 ;
      RECT 44.38 1.68 45.13 1.87 ;
      RECT 42.495 1.235 42.69 1.565 ;
      RECT 43.2 1.855 44.21 2.025 ;
      RECT 44.02 0.495 44.21 2.025 ;
      RECT 43.2 1.055 43.37 2.025 ;
      RECT 42.86 2.195 43.985 2.365 ;
      RECT 42.86 0.495 43.03 2.365 ;
      RECT 42.015 1.235 42.27 1.565 ;
      RECT 42.1 0.895 42.27 1.565 ;
      RECT 42.1 0.895 43.03 1.065 ;
      RECT 42.855 0.495 43.03 1.065 ;
      RECT 42.855 0.495 43.385 0.86 ;
      RECT 41.675 1.735 42.01 2.705 ;
      RECT 41.675 0.495 41.845 2.705 ;
      RECT 41.675 0.495 41.93 1.065 ;
      RECT 40.58 0.715 41.31 0.955 ;
      RECT 41.122 0.51 41.31 0.955 ;
      RECT 40.95 0.522 41.325 0.949 ;
      RECT 40.865 0.537 41.345 0.934 ;
      RECT 40.865 0.552 41.35 0.924 ;
      RECT 40.82 0.572 41.365 0.916 ;
      RECT 40.797 0.607 41.38 0.87 ;
      RECT 40.711 0.63 41.385 0.83 ;
      RECT 40.711 0.648 41.395 0.8 ;
      RECT 40.58 0.717 41.4 0.763 ;
      RECT 40.625 0.66 41.395 0.8 ;
      RECT 40.711 0.612 41.38 0.87 ;
      RECT 40.797 0.581 41.365 0.916 ;
      RECT 40.82 0.562 41.35 0.924 ;
      RECT 40.865 0.535 41.325 0.949 ;
      RECT 40.95 0.517 41.31 0.955 ;
      RECT 41.036 0.511 41.31 0.955 ;
      RECT 41.122 0.506 41.255 0.955 ;
      RECT 41.208 0.501 41.255 0.955 ;
      RECT 40.9 1.399 41.07 1.785 ;
      RECT 40.895 1.399 41.07 1.78 ;
      RECT 40.87 1.399 41.07 1.745 ;
      RECT 40.87 1.427 41.08 1.735 ;
      RECT 40.85 1.427 41.08 1.695 ;
      RECT 40.845 1.427 41.08 1.668 ;
      RECT 40.845 1.445 41.085 1.66 ;
      RECT 40.79 1.445 41.085 1.595 ;
      RECT 40.79 1.462 41.095 1.578 ;
      RECT 40.78 1.462 41.095 1.518 ;
      RECT 40.78 1.479 41.1 1.515 ;
      RECT 40.775 1.315 40.945 1.493 ;
      RECT 40.775 1.349 41.031 1.493 ;
      RECT 40.77 2.115 40.775 2.128 ;
      RECT 40.765 2.01 40.77 2.133 ;
      RECT 40.74 1.87 40.765 2.148 ;
      RECT 40.705 1.821 40.74 2.18 ;
      RECT 40.7 1.789 40.705 2.2 ;
      RECT 40.695 1.78 40.7 2.2 ;
      RECT 40.615 1.745 40.695 2.2 ;
      RECT 40.552 1.715 40.615 2.2 ;
      RECT 40.466 1.703 40.552 2.2 ;
      RECT 40.38 1.689 40.466 2.2 ;
      RECT 40.3 1.676 40.38 2.186 ;
      RECT 40.265 1.668 40.3 2.166 ;
      RECT 40.255 1.665 40.265 2.157 ;
      RECT 40.225 1.66 40.255 2.144 ;
      RECT 40.175 1.635 40.225 2.12 ;
      RECT 40.161 1.609 40.175 2.102 ;
      RECT 40.075 1.569 40.161 2.078 ;
      RECT 40.03 1.517 40.075 2.047 ;
      RECT 40.02 1.492 40.03 2.034 ;
      RECT 40.015 1.273 40.02 1.295 ;
      RECT 40.01 1.475 40.02 2.03 ;
      RECT 40.01 1.271 40.015 1.385 ;
      RECT 40 1.267 40.01 2.026 ;
      RECT 39.956 1.265 40 2.014 ;
      RECT 39.87 1.265 39.956 1.985 ;
      RECT 39.84 1.265 39.87 1.958 ;
      RECT 39.825 1.265 39.84 1.946 ;
      RECT 39.785 1.277 39.825 1.931 ;
      RECT 39.765 1.296 39.785 1.91 ;
      RECT 39.755 1.306 39.765 1.894 ;
      RECT 39.745 1.312 39.755 1.883 ;
      RECT 39.725 1.322 39.745 1.866 ;
      RECT 39.72 1.331 39.725 1.853 ;
      RECT 39.715 1.335 39.72 1.803 ;
      RECT 39.705 1.341 39.715 1.72 ;
      RECT 39.7 1.345 39.705 1.634 ;
      RECT 39.695 1.365 39.7 1.571 ;
      RECT 39.69 1.388 39.695 1.518 ;
      RECT 39.685 1.406 39.69 1.463 ;
      RECT 40.295 1.225 40.465 1.485 ;
      RECT 40.465 1.19 40.51 1.471 ;
      RECT 40.426 1.192 40.515 1.454 ;
      RECT 40.315 1.209 40.601 1.425 ;
      RECT 40.315 1.224 40.605 1.397 ;
      RECT 40.315 1.205 40.515 1.454 ;
      RECT 40.34 1.193 40.465 1.485 ;
      RECT 40.426 1.191 40.51 1.471 ;
      RECT 39.48 0.58 39.65 1.07 ;
      RECT 39.48 0.58 39.685 1.05 ;
      RECT 39.615 0.5 39.725 1.01 ;
      RECT 39.596 0.504 39.745 0.98 ;
      RECT 39.51 0.512 39.765 0.963 ;
      RECT 39.51 0.518 39.77 0.953 ;
      RECT 39.51 0.527 39.79 0.941 ;
      RECT 39.485 0.552 39.82 0.919 ;
      RECT 39.485 0.572 39.825 0.899 ;
      RECT 39.48 0.585 39.835 0.879 ;
      RECT 39.48 0.652 39.84 0.86 ;
      RECT 39.48 0.785 39.845 0.847 ;
      RECT 39.475 0.59 39.835 0.68 ;
      RECT 39.485 0.547 39.79 0.941 ;
      RECT 39.596 0.502 39.725 1.01 ;
      RECT 39.47 2.255 39.77 2.51 ;
      RECT 39.555 2.221 39.77 2.51 ;
      RECT 39.555 2.224 39.775 2.37 ;
      RECT 39.49 2.245 39.775 2.37 ;
      RECT 39.525 2.235 39.77 2.51 ;
      RECT 39.52 2.24 39.775 2.37 ;
      RECT 39.555 2.219 39.756 2.51 ;
      RECT 39.641 2.21 39.756 2.51 ;
      RECT 39.641 2.204 39.67 2.51 ;
      RECT 39.13 1.845 39.14 2.335 ;
      RECT 38.79 1.78 38.8 2.08 ;
      RECT 39.305 1.952 39.31 2.171 ;
      RECT 39.295 1.932 39.305 2.188 ;
      RECT 39.285 1.912 39.295 2.218 ;
      RECT 39.28 1.902 39.285 2.233 ;
      RECT 39.275 1.898 39.28 2.238 ;
      RECT 39.26 1.89 39.275 2.245 ;
      RECT 39.22 1.87 39.26 2.27 ;
      RECT 39.195 1.852 39.22 2.303 ;
      RECT 39.19 1.85 39.195 2.316 ;
      RECT 39.17 1.847 39.19 2.32 ;
      RECT 39.14 1.845 39.17 2.33 ;
      RECT 39.07 1.847 39.13 2.331 ;
      RECT 39.05 1.847 39.07 2.325 ;
      RECT 39.025 1.845 39.05 2.322 ;
      RECT 38.99 1.84 39.025 2.318 ;
      RECT 38.97 1.834 38.99 2.305 ;
      RECT 38.96 1.831 38.97 2.293 ;
      RECT 38.94 1.828 38.96 2.278 ;
      RECT 38.92 1.824 38.94 2.26 ;
      RECT 38.915 1.821 38.92 2.25 ;
      RECT 38.91 1.82 38.915 2.248 ;
      RECT 38.9 1.817 38.91 2.24 ;
      RECT 38.89 1.811 38.9 2.223 ;
      RECT 38.88 1.805 38.89 2.205 ;
      RECT 38.87 1.799 38.88 2.193 ;
      RECT 38.86 1.793 38.87 2.173 ;
      RECT 38.855 1.789 38.86 2.158 ;
      RECT 38.85 1.787 38.855 2.15 ;
      RECT 38.845 1.785 38.85 2.143 ;
      RECT 38.84 1.783 38.845 2.133 ;
      RECT 38.835 1.781 38.84 2.127 ;
      RECT 38.825 1.78 38.835 2.117 ;
      RECT 38.815 1.78 38.825 2.108 ;
      RECT 38.8 1.78 38.815 2.093 ;
      RECT 38.76 1.78 38.79 2.077 ;
      RECT 38.74 1.782 38.76 2.072 ;
      RECT 38.735 1.787 38.74 2.07 ;
      RECT 38.705 1.795 38.735 2.068 ;
      RECT 38.675 1.81 38.705 2.067 ;
      RECT 38.63 1.832 38.675 2.072 ;
      RECT 38.625 1.847 38.63 2.076 ;
      RECT 38.61 1.852 38.625 2.078 ;
      RECT 38.605 1.856 38.61 2.08 ;
      RECT 38.545 1.879 38.605 2.089 ;
      RECT 38.525 1.905 38.545 2.102 ;
      RECT 38.515 1.912 38.525 2.106 ;
      RECT 38.5 1.919 38.515 2.109 ;
      RECT 38.48 1.929 38.5 2.112 ;
      RECT 38.475 1.937 38.48 2.115 ;
      RECT 38.43 1.942 38.475 2.122 ;
      RECT 38.42 1.945 38.43 2.129 ;
      RECT 38.41 1.945 38.42 2.133 ;
      RECT 38.375 1.947 38.41 2.145 ;
      RECT 38.355 1.95 38.375 2.158 ;
      RECT 38.315 1.953 38.355 2.169 ;
      RECT 38.3 1.955 38.315 2.182 ;
      RECT 38.29 1.955 38.3 2.187 ;
      RECT 38.265 1.956 38.29 2.195 ;
      RECT 38.255 1.958 38.265 2.2 ;
      RECT 38.25 1.959 38.255 2.203 ;
      RECT 38.225 1.957 38.25 2.206 ;
      RECT 38.21 1.955 38.225 2.207 ;
      RECT 38.19 1.952 38.21 2.209 ;
      RECT 38.17 1.947 38.19 2.209 ;
      RECT 38.11 1.942 38.17 2.206 ;
      RECT 38.075 1.917 38.11 2.202 ;
      RECT 38.065 1.894 38.075 2.2 ;
      RECT 38.035 1.871 38.065 2.2 ;
      RECT 38.025 1.85 38.035 2.2 ;
      RECT 38 1.832 38.025 2.198 ;
      RECT 37.985 1.81 38 2.195 ;
      RECT 37.97 1.792 37.985 2.193 ;
      RECT 37.95 1.782 37.97 2.191 ;
      RECT 37.935 1.777 37.95 2.19 ;
      RECT 37.92 1.775 37.935 2.189 ;
      RECT 37.89 1.776 37.92 2.187 ;
      RECT 37.87 1.779 37.89 2.185 ;
      RECT 37.813 1.783 37.87 2.185 ;
      RECT 37.727 1.792 37.813 2.185 ;
      RECT 37.641 1.803 37.727 2.185 ;
      RECT 37.555 1.814 37.641 2.185 ;
      RECT 37.535 1.821 37.555 2.193 ;
      RECT 37.525 1.824 37.535 2.2 ;
      RECT 37.46 1.829 37.525 2.218 ;
      RECT 37.43 1.836 37.46 2.243 ;
      RECT 37.42 1.839 37.43 2.25 ;
      RECT 37.375 1.843 37.42 2.255 ;
      RECT 37.345 1.848 37.375 2.26 ;
      RECT 37.344 1.85 37.345 2.26 ;
      RECT 37.258 1.856 37.344 2.26 ;
      RECT 37.172 1.867 37.258 2.26 ;
      RECT 37.086 1.879 37.172 2.26 ;
      RECT 37 1.89 37.086 2.26 ;
      RECT 36.985 1.897 37 2.255 ;
      RECT 36.98 1.899 36.985 2.249 ;
      RECT 36.96 1.91 36.98 2.244 ;
      RECT 36.95 1.928 36.96 2.238 ;
      RECT 36.945 1.94 36.95 2.038 ;
      RECT 39.24 0.693 39.26 0.78 ;
      RECT 39.235 0.628 39.24 0.812 ;
      RECT 39.225 0.595 39.235 0.817 ;
      RECT 39.22 0.575 39.225 0.823 ;
      RECT 39.19 0.575 39.22 0.84 ;
      RECT 39.141 0.575 39.19 0.876 ;
      RECT 39.055 0.575 39.141 0.934 ;
      RECT 39.026 0.585 39.055 0.983 ;
      RECT 38.94 0.627 39.026 1.036 ;
      RECT 38.92 0.665 38.94 1.083 ;
      RECT 38.895 0.682 38.92 1.103 ;
      RECT 38.885 0.696 38.895 1.123 ;
      RECT 38.88 0.702 38.885 1.133 ;
      RECT 38.875 0.706 38.88 1.14 ;
      RECT 38.825 0.726 38.875 1.145 ;
      RECT 38.76 0.77 38.825 1.145 ;
      RECT 38.735 0.82 38.76 1.145 ;
      RECT 38.725 0.85 38.735 1.145 ;
      RECT 38.72 0.877 38.725 1.145 ;
      RECT 38.715 0.895 38.72 1.145 ;
      RECT 38.705 0.937 38.715 1.145 ;
      RECT 39.055 1.495 39.225 1.67 ;
      RECT 38.995 1.323 39.055 1.658 ;
      RECT 38.985 1.316 38.995 1.641 ;
      RECT 38.94 1.495 39.225 1.621 ;
      RECT 38.921 1.495 39.225 1.599 ;
      RECT 38.835 1.495 39.225 1.564 ;
      RECT 38.815 1.315 38.985 1.52 ;
      RECT 38.815 1.462 39.22 1.52 ;
      RECT 38.815 1.41 39.195 1.52 ;
      RECT 38.815 1.365 39.16 1.52 ;
      RECT 38.815 1.347 39.125 1.52 ;
      RECT 38.815 1.337 39.12 1.52 ;
      RECT 38.535 2.295 38.725 2.52 ;
      RECT 38.525 2.296 38.73 2.515 ;
      RECT 38.525 2.298 38.74 2.495 ;
      RECT 38.525 2.302 38.745 2.48 ;
      RECT 38.525 2.289 38.695 2.515 ;
      RECT 38.525 2.292 38.72 2.515 ;
      RECT 38.535 2.288 38.695 2.52 ;
      RECT 38.621 2.286 38.695 2.52 ;
      RECT 38.245 1.537 38.415 1.775 ;
      RECT 38.245 1.537 38.501 1.689 ;
      RECT 38.245 1.537 38.505 1.599 ;
      RECT 38.295 1.31 38.515 1.578 ;
      RECT 38.29 1.327 38.52 1.551 ;
      RECT 38.255 1.485 38.52 1.551 ;
      RECT 38.275 1.335 38.415 1.775 ;
      RECT 38.265 1.417 38.525 1.534 ;
      RECT 38.26 1.465 38.525 1.534 ;
      RECT 38.265 1.375 38.52 1.551 ;
      RECT 38.29 1.312 38.515 1.578 ;
      RECT 37.855 1.287 38.025 1.485 ;
      RECT 37.855 1.287 38.07 1.46 ;
      RECT 37.925 1.23 38.095 1.418 ;
      RECT 37.9 1.245 38.095 1.418 ;
      RECT 37.515 1.291 37.545 1.485 ;
      RECT 37.51 1.263 37.515 1.485 ;
      RECT 37.48 1.237 37.51 1.487 ;
      RECT 37.455 1.195 37.48 1.49 ;
      RECT 37.445 1.167 37.455 1.492 ;
      RECT 37.41 1.147 37.445 1.494 ;
      RECT 37.345 1.132 37.41 1.5 ;
      RECT 37.295 1.13 37.345 1.506 ;
      RECT 37.272 1.132 37.295 1.511 ;
      RECT 37.186 1.143 37.272 1.517 ;
      RECT 37.1 1.161 37.186 1.527 ;
      RECT 37.085 1.172 37.1 1.533 ;
      RECT 37.015 1.195 37.085 1.539 ;
      RECT 36.96 1.227 37.015 1.547 ;
      RECT 36.92 1.25 36.96 1.553 ;
      RECT 36.906 1.263 36.92 1.556 ;
      RECT 36.82 1.285 36.906 1.562 ;
      RECT 36.805 1.31 36.82 1.568 ;
      RECT 36.765 1.325 36.805 1.572 ;
      RECT 36.715 1.34 36.765 1.577 ;
      RECT 36.69 1.347 36.715 1.581 ;
      RECT 36.63 1.342 36.69 1.585 ;
      RECT 36.615 1.333 36.63 1.589 ;
      RECT 36.545 1.323 36.615 1.585 ;
      RECT 36.52 1.315 36.54 1.575 ;
      RECT 36.461 1.315 36.52 1.553 ;
      RECT 36.375 1.315 36.461 1.51 ;
      RECT 36.54 1.315 36.545 1.58 ;
      RECT 37.235 0.546 37.405 0.88 ;
      RECT 37.205 0.546 37.405 0.875 ;
      RECT 37.145 0.513 37.205 0.863 ;
      RECT 37.145 0.569 37.415 0.858 ;
      RECT 37.12 0.569 37.415 0.852 ;
      RECT 37.115 0.51 37.145 0.849 ;
      RECT 37.1 0.516 37.235 0.847 ;
      RECT 37.095 0.524 37.32 0.835 ;
      RECT 37.095 0.576 37.43 0.788 ;
      RECT 37.08 0.532 37.32 0.783 ;
      RECT 37.08 0.602 37.44 0.724 ;
      RECT 37.05 0.552 37.405 0.685 ;
      RECT 37.05 0.642 37.45 0.681 ;
      RECT 37.1 0.521 37.32 0.847 ;
      RECT 36.44 0.851 36.495 1.115 ;
      RECT 36.44 0.851 36.56 1.114 ;
      RECT 36.44 0.851 36.585 1.113 ;
      RECT 36.44 0.851 36.65 1.112 ;
      RECT 36.585 0.817 36.665 1.111 ;
      RECT 36.4 0.861 36.81 1.11 ;
      RECT 36.44 0.858 36.81 1.11 ;
      RECT 36.4 0.866 36.815 1.103 ;
      RECT 36.385 0.868 36.815 1.102 ;
      RECT 36.385 0.875 36.82 1.098 ;
      RECT 36.365 0.874 36.815 1.094 ;
      RECT 36.365 0.882 36.825 1.093 ;
      RECT 36.36 0.879 36.82 1.089 ;
      RECT 36.36 0.892 36.835 1.088 ;
      RECT 36.345 0.882 36.825 1.087 ;
      RECT 36.31 0.895 36.835 1.08 ;
      RECT 36.495 0.85 36.805 1.11 ;
      RECT 36.495 0.835 36.755 1.11 ;
      RECT 36.56 0.822 36.69 1.11 ;
      RECT 36.105 1.911 36.12 2.304 ;
      RECT 36.07 1.916 36.12 2.303 ;
      RECT 36.105 1.915 36.165 2.302 ;
      RECT 36.05 1.926 36.165 2.301 ;
      RECT 36.065 1.922 36.165 2.301 ;
      RECT 36.03 1.932 36.24 2.298 ;
      RECT 36.03 1.951 36.285 2.296 ;
      RECT 36.03 1.958 36.29 2.293 ;
      RECT 36.015 1.935 36.24 2.29 ;
      RECT 35.995 1.94 36.24 2.283 ;
      RECT 35.99 1.944 36.24 2.279 ;
      RECT 35.99 1.961 36.3 2.278 ;
      RECT 35.97 1.955 36.285 2.274 ;
      RECT 35.97 1.964 36.305 2.268 ;
      RECT 35.965 1.97 36.305 2.04 ;
      RECT 36.03 1.93 36.165 2.298 ;
      RECT 35.905 1.293 36.105 1.605 ;
      RECT 35.98 1.271 36.105 1.605 ;
      RECT 35.92 1.29 36.11 1.59 ;
      RECT 35.89 1.301 36.11 1.588 ;
      RECT 35.905 1.296 36.115 1.554 ;
      RECT 35.89 1.4 36.12 1.521 ;
      RECT 35.92 1.272 36.105 1.605 ;
      RECT 35.98 1.25 36.08 1.605 ;
      RECT 36.005 1.247 36.08 1.605 ;
      RECT 36.005 1.242 36.025 1.605 ;
      RECT 35.41 1.31 35.585 1.485 ;
      RECT 35.405 1.31 35.585 1.483 ;
      RECT 35.38 1.31 35.585 1.478 ;
      RECT 35.325 1.29 35.495 1.468 ;
      RECT 35.325 1.297 35.56 1.468 ;
      RECT 35.41 1.977 35.425 2.16 ;
      RECT 35.4 1.955 35.41 2.16 ;
      RECT 35.385 1.935 35.4 2.16 ;
      RECT 35.375 1.91 35.385 2.16 ;
      RECT 35.345 1.875 35.375 2.16 ;
      RECT 35.31 1.815 35.345 2.16 ;
      RECT 35.305 1.777 35.31 2.16 ;
      RECT 35.255 1.728 35.305 2.16 ;
      RECT 35.245 1.678 35.255 2.148 ;
      RECT 35.23 1.657 35.245 2.108 ;
      RECT 35.21 1.625 35.23 2.058 ;
      RECT 35.185 1.581 35.21 1.998 ;
      RECT 35.18 1.553 35.185 1.953 ;
      RECT 35.175 1.544 35.18 1.939 ;
      RECT 35.17 1.537 35.175 1.926 ;
      RECT 35.165 1.532 35.17 1.915 ;
      RECT 35.16 1.517 35.165 1.905 ;
      RECT 35.155 1.495 35.16 1.892 ;
      RECT 35.145 1.455 35.155 1.867 ;
      RECT 35.12 1.385 35.145 1.823 ;
      RECT 35.115 1.325 35.12 1.788 ;
      RECT 35.1 1.305 35.115 1.755 ;
      RECT 35.095 1.305 35.1 1.73 ;
      RECT 35.065 1.305 35.095 1.685 ;
      RECT 35.02 1.305 35.065 1.625 ;
      RECT 34.945 1.305 35.02 1.573 ;
      RECT 34.94 1.305 34.945 1.538 ;
      RECT 34.935 1.305 34.94 1.528 ;
      RECT 34.93 1.305 34.935 1.508 ;
      RECT 35.195 0.525 35.365 0.995 ;
      RECT 35.14 0.518 35.335 0.979 ;
      RECT 35.14 0.532 35.37 0.978 ;
      RECT 35.125 0.533 35.37 0.959 ;
      RECT 35.12 0.551 35.37 0.945 ;
      RECT 35.125 0.534 35.375 0.943 ;
      RECT 35.11 0.565 35.375 0.928 ;
      RECT 35.125 0.54 35.38 0.913 ;
      RECT 35.105 0.58 35.38 0.91 ;
      RECT 35.12 0.552 35.385 0.895 ;
      RECT 35.12 0.564 35.39 0.875 ;
      RECT 35.105 0.58 35.395 0.858 ;
      RECT 35.105 0.59 35.4 0.713 ;
      RECT 35.1 0.59 35.4 0.67 ;
      RECT 35.1 0.605 35.405 0.648 ;
      RECT 35.195 0.515 35.335 0.995 ;
      RECT 35.195 0.513 35.305 0.995 ;
      RECT 35.281 0.51 35.305 0.995 ;
      RECT 34.94 2.177 34.945 2.223 ;
      RECT 34.93 2.025 34.94 2.247 ;
      RECT 34.925 1.87 34.93 2.272 ;
      RECT 34.91 1.832 34.925 2.283 ;
      RECT 34.905 1.815 34.91 2.29 ;
      RECT 34.895 1.803 34.905 2.297 ;
      RECT 34.89 1.794 34.895 2.299 ;
      RECT 34.885 1.792 34.89 2.303 ;
      RECT 34.84 1.783 34.885 2.318 ;
      RECT 34.835 1.775 34.84 2.332 ;
      RECT 34.83 1.772 34.835 2.336 ;
      RECT 34.815 1.767 34.83 2.344 ;
      RECT 34.76 1.757 34.815 2.355 ;
      RECT 34.725 1.745 34.76 2.356 ;
      RECT 34.716 1.74 34.725 2.35 ;
      RECT 34.63 1.74 34.716 2.34 ;
      RECT 34.6 1.74 34.63 2.318 ;
      RECT 34.59 1.74 34.595 2.298 ;
      RECT 34.585 1.74 34.59 2.26 ;
      RECT 34.58 1.74 34.585 2.218 ;
      RECT 34.575 1.74 34.58 2.178 ;
      RECT 34.57 1.74 34.575 2.108 ;
      RECT 34.56 1.74 34.57 2.03 ;
      RECT 34.555 1.74 34.56 1.93 ;
      RECT 34.595 1.74 34.6 2.3 ;
      RECT 34.09 1.822 34.18 2.3 ;
      RECT 34.075 1.825 34.195 2.298 ;
      RECT 34.09 1.824 34.195 2.298 ;
      RECT 34.055 1.831 34.22 2.288 ;
      RECT 34.075 1.825 34.22 2.288 ;
      RECT 34.04 1.837 34.22 2.276 ;
      RECT 34.075 1.828 34.27 2.269 ;
      RECT 34.026 1.845 34.27 2.267 ;
      RECT 34.055 1.835 34.28 2.255 ;
      RECT 34.026 1.856 34.31 2.246 ;
      RECT 33.94 1.88 34.31 2.24 ;
      RECT 33.94 1.893 34.35 2.223 ;
      RECT 33.935 1.915 34.35 2.216 ;
      RECT 33.905 1.93 34.35 2.206 ;
      RECT 33.9 1.941 34.35 2.196 ;
      RECT 33.87 1.954 34.35 2.187 ;
      RECT 33.855 1.972 34.35 2.176 ;
      RECT 33.83 1.985 34.35 2.166 ;
      RECT 34.09 1.821 34.1 2.3 ;
      RECT 34.136 1.245 34.175 1.49 ;
      RECT 34.05 1.245 34.185 1.488 ;
      RECT 33.935 1.27 34.185 1.485 ;
      RECT 33.935 1.27 34.19 1.483 ;
      RECT 33.935 1.27 34.205 1.478 ;
      RECT 34.041 1.245 34.22 1.458 ;
      RECT 33.955 1.253 34.22 1.458 ;
      RECT 33.625 0.605 33.795 1.04 ;
      RECT 33.615 0.639 33.795 1.023 ;
      RECT 33.695 0.575 33.865 1.01 ;
      RECT 33.6 0.65 33.865 0.988 ;
      RECT 33.695 0.585 33.87 0.978 ;
      RECT 33.625 0.637 33.9 0.963 ;
      RECT 33.585 0.663 33.9 0.948 ;
      RECT 33.585 0.705 33.91 0.928 ;
      RECT 33.58 0.73 33.915 0.91 ;
      RECT 33.58 0.74 33.92 0.895 ;
      RECT 33.575 0.677 33.9 0.893 ;
      RECT 33.575 0.75 33.925 0.878 ;
      RECT 33.57 0.687 33.9 0.875 ;
      RECT 33.565 0.771 33.93 0.858 ;
      RECT 33.565 0.803 33.935 0.838 ;
      RECT 33.56 0.717 33.91 0.83 ;
      RECT 33.565 0.702 33.9 0.858 ;
      RECT 33.58 0.672 33.9 0.91 ;
      RECT 33.425 1.259 33.65 1.515 ;
      RECT 33.425 1.292 33.67 1.505 ;
      RECT 33.39 1.292 33.67 1.503 ;
      RECT 33.39 1.305 33.675 1.493 ;
      RECT 33.39 1.325 33.685 1.485 ;
      RECT 33.39 1.422 33.69 1.478 ;
      RECT 33.37 1.17 33.5 1.468 ;
      RECT 33.325 1.325 33.685 1.41 ;
      RECT 33.315 1.17 33.5 1.355 ;
      RECT 33.315 1.202 33.586 1.355 ;
      RECT 33.28 1.732 33.3 1.91 ;
      RECT 33.245 1.685 33.28 1.91 ;
      RECT 33.23 1.625 33.245 1.91 ;
      RECT 33.205 1.572 33.23 1.91 ;
      RECT 33.19 1.525 33.205 1.91 ;
      RECT 33.17 1.502 33.19 1.91 ;
      RECT 33.145 1.467 33.17 1.91 ;
      RECT 33.135 1.313 33.145 1.91 ;
      RECT 33.105 1.308 33.135 1.901 ;
      RECT 33.1 1.305 33.105 1.891 ;
      RECT 33.085 1.305 33.1 1.865 ;
      RECT 33.08 1.305 33.085 1.828 ;
      RECT 33.055 1.305 33.08 1.78 ;
      RECT 33.035 1.305 33.055 1.705 ;
      RECT 33.025 1.305 33.035 1.665 ;
      RECT 33.02 1.305 33.025 1.64 ;
      RECT 33.015 1.305 33.02 1.623 ;
      RECT 33.01 1.305 33.015 1.605 ;
      RECT 33.005 1.306 33.01 1.595 ;
      RECT 32.995 1.308 33.005 1.563 ;
      RECT 32.985 1.31 32.995 1.53 ;
      RECT 32.975 1.313 32.985 1.503 ;
      RECT 33.3 1.74 33.525 1.91 ;
      RECT 32.63 0.552 32.8 1.005 ;
      RECT 32.63 0.552 32.89 0.971 ;
      RECT 32.63 0.552 32.92 0.955 ;
      RECT 32.63 0.552 32.95 0.928 ;
      RECT 32.886 0.53 32.965 0.91 ;
      RECT 32.665 0.537 32.97 0.895 ;
      RECT 32.665 0.545 32.98 0.858 ;
      RECT 32.625 0.572 32.98 0.83 ;
      RECT 32.61 0.585 32.98 0.795 ;
      RECT 32.63 0.56 33 0.785 ;
      RECT 32.605 0.625 33 0.755 ;
      RECT 32.605 0.655 33.005 0.738 ;
      RECT 32.6 0.685 33.005 0.725 ;
      RECT 32.665 0.534 32.965 0.91 ;
      RECT 32.8 0.531 32.886 0.989 ;
      RECT 32.751 0.532 32.965 0.91 ;
      RECT 32.895 2.192 32.94 2.385 ;
      RECT 32.885 2.162 32.895 2.385 ;
      RECT 32.88 2.147 32.885 2.385 ;
      RECT 32.84 2.057 32.88 2.385 ;
      RECT 32.835 1.97 32.84 2.385 ;
      RECT 32.825 1.94 32.835 2.385 ;
      RECT 32.82 1.9 32.825 2.385 ;
      RECT 32.81 1.862 32.82 2.385 ;
      RECT 32.805 1.827 32.81 2.385 ;
      RECT 32.785 1.78 32.805 2.385 ;
      RECT 32.77 1.705 32.785 2.385 ;
      RECT 32.765 1.66 32.77 2.38 ;
      RECT 32.76 1.64 32.765 2.353 ;
      RECT 32.755 1.62 32.76 2.338 ;
      RECT 32.75 1.595 32.755 2.318 ;
      RECT 32.745 1.573 32.75 2.303 ;
      RECT 32.74 1.551 32.745 2.285 ;
      RECT 32.735 1.53 32.74 2.275 ;
      RECT 32.725 1.502 32.735 2.245 ;
      RECT 32.715 1.465 32.725 2.213 ;
      RECT 32.705 1.425 32.715 2.18 ;
      RECT 32.695 1.403 32.705 2.15 ;
      RECT 32.665 1.355 32.695 2.082 ;
      RECT 32.65 1.315 32.665 2.009 ;
      RECT 32.64 1.315 32.65 1.975 ;
      RECT 32.635 1.315 32.64 1.95 ;
      RECT 32.63 1.315 32.635 1.935 ;
      RECT 32.625 1.315 32.63 1.913 ;
      RECT 32.62 1.315 32.625 1.9 ;
      RECT 32.605 1.315 32.62 1.865 ;
      RECT 32.585 1.315 32.605 1.805 ;
      RECT 32.575 1.315 32.585 1.755 ;
      RECT 32.555 1.315 32.575 1.703 ;
      RECT 32.535 1.315 32.555 1.66 ;
      RECT 32.525 1.315 32.535 1.648 ;
      RECT 32.495 1.315 32.525 1.635 ;
      RECT 32.465 1.336 32.495 1.615 ;
      RECT 32.455 1.364 32.465 1.595 ;
      RECT 32.44 1.381 32.455 1.563 ;
      RECT 32.435 1.395 32.44 1.53 ;
      RECT 32.43 1.403 32.435 1.503 ;
      RECT 32.425 1.411 32.43 1.465 ;
      RECT 32.43 1.935 32.435 2.27 ;
      RECT 32.395 1.922 32.43 2.269 ;
      RECT 32.325 1.862 32.395 2.268 ;
      RECT 32.245 1.805 32.325 2.267 ;
      RECT 32.11 1.765 32.245 2.266 ;
      RECT 32.11 1.952 32.445 2.255 ;
      RECT 32.07 1.952 32.445 2.245 ;
      RECT 32.07 1.97 32.45 2.24 ;
      RECT 32.07 2.06 32.455 2.23 ;
      RECT 32.065 1.755 32.23 2.21 ;
      RECT 32.06 1.755 32.23 1.953 ;
      RECT 32.06 1.912 32.425 1.953 ;
      RECT 32.06 1.9 32.42 1.953 ;
      RECT 31.325 2.115 31.84 2.525 ;
      RECT 31.5 1.135 31.84 2.525 ;
      RECT 30.61 1.135 31.84 1.305 ;
      RECT 31.32 0.53 31.565 1.305 ;
      RECT 28.72 2.535 30.75 2.705 ;
      RECT 30.58 1.68 30.75 2.705 ;
      RECT 28.72 1.235 28.89 2.705 ;
      RECT 30.58 1.68 31.33 1.87 ;
      RECT 28.695 1.235 28.89 1.565 ;
      RECT 29.4 1.855 30.41 2.025 ;
      RECT 30.22 0.495 30.41 2.025 ;
      RECT 29.4 1.055 29.57 2.025 ;
      RECT 29.06 2.195 30.185 2.365 ;
      RECT 29.06 0.495 29.23 2.365 ;
      RECT 28.215 1.235 28.47 1.565 ;
      RECT 28.3 0.895 28.47 1.565 ;
      RECT 28.3 0.895 29.23 1.065 ;
      RECT 29.055 0.495 29.23 1.065 ;
      RECT 29.055 0.495 29.585 0.86 ;
      RECT 27.875 1.735 28.21 2.705 ;
      RECT 27.875 0.495 28.045 2.705 ;
      RECT 27.875 0.495 28.13 1.065 ;
      RECT 27.125 1.725 27.455 2.705 ;
      RECT 27.225 0.495 27.455 2.705 ;
      RECT 27.125 0.495 27.455 1.125 ;
      RECT 25.745 1.725 26.075 2.705 ;
      RECT 25.845 0.495 26.075 2.705 ;
      RECT 25.845 1.315 27.055 1.555 ;
      RECT 25.745 0.495 26.075 1.125 ;
      RECT 24.365 1.725 24.695 2.705 ;
      RECT 24.465 0.495 24.695 2.705 ;
      RECT 24.365 0.495 24.695 1.125 ;
      RECT 22.985 1.725 23.315 2.705 ;
      RECT 23.085 0.495 23.315 2.705 ;
      RECT 23.085 1.315 24.295 1.555 ;
      RECT 22.985 0.495 23.315 1.125 ;
      RECT 21.665 2.115 22.18 2.525 ;
      RECT 21.84 1.135 22.18 2.525 ;
      RECT 20.95 1.135 22.18 1.305 ;
      RECT 21.66 0.53 21.905 1.305 ;
      RECT 19.06 2.535 21.09 2.705 ;
      RECT 20.92 1.68 21.09 2.705 ;
      RECT 19.06 1.235 19.23 2.705 ;
      RECT 20.92 1.68 21.67 1.87 ;
      RECT 19.035 1.235 19.23 1.565 ;
      RECT 19.74 1.855 20.75 2.025 ;
      RECT 20.56 0.495 20.75 2.025 ;
      RECT 19.74 1.055 19.91 2.025 ;
      RECT 19.4 2.195 20.525 2.365 ;
      RECT 19.4 0.495 19.57 2.365 ;
      RECT 18.555 1.235 18.81 1.565 ;
      RECT 18.64 0.895 18.81 1.565 ;
      RECT 18.64 0.895 19.57 1.065 ;
      RECT 19.395 0.495 19.57 1.065 ;
      RECT 19.395 0.495 19.925 0.86 ;
      RECT 18.215 1.735 18.55 2.705 ;
      RECT 18.215 0.495 18.385 2.705 ;
      RECT 18.215 0.495 18.47 1.065 ;
      RECT 17.53 2.115 18.045 2.525 ;
      RECT 17.705 1.135 18.045 2.525 ;
      RECT 16.815 1.135 18.045 1.305 ;
      RECT 17.525 0.53 17.77 1.305 ;
      RECT 14.925 2.535 16.955 2.705 ;
      RECT 16.785 1.68 16.955 2.705 ;
      RECT 14.925 1.235 15.095 2.705 ;
      RECT 16.785 1.68 17.535 1.87 ;
      RECT 14.9 1.235 15.095 1.565 ;
      RECT 15.605 1.855 16.615 2.025 ;
      RECT 16.425 0.495 16.615 2.025 ;
      RECT 15.605 1.055 15.775 2.025 ;
      RECT 15.265 2.195 16.39 2.365 ;
      RECT 15.265 0.495 15.435 2.365 ;
      RECT 14.42 1.235 14.675 1.565 ;
      RECT 14.505 0.895 14.675 1.565 ;
      RECT 14.505 0.895 15.435 1.065 ;
      RECT 15.26 0.495 15.435 1.065 ;
      RECT 15.26 0.495 15.79 0.86 ;
      RECT 14.08 1.735 14.415 2.705 ;
      RECT 14.08 0.495 14.25 2.705 ;
      RECT 14.08 0.495 14.335 1.065 ;
      RECT 12.985 0.715 13.715 0.955 ;
      RECT 13.527 0.51 13.715 0.955 ;
      RECT 13.355 0.522 13.73 0.949 ;
      RECT 13.27 0.537 13.75 0.934 ;
      RECT 13.27 0.552 13.755 0.924 ;
      RECT 13.225 0.572 13.77 0.916 ;
      RECT 13.202 0.607 13.785 0.87 ;
      RECT 13.116 0.63 13.79 0.83 ;
      RECT 13.116 0.648 13.8 0.8 ;
      RECT 12.985 0.717 13.805 0.763 ;
      RECT 13.03 0.66 13.8 0.8 ;
      RECT 13.116 0.612 13.785 0.87 ;
      RECT 13.202 0.581 13.77 0.916 ;
      RECT 13.225 0.562 13.755 0.924 ;
      RECT 13.27 0.535 13.73 0.949 ;
      RECT 13.355 0.517 13.715 0.955 ;
      RECT 13.441 0.511 13.715 0.955 ;
      RECT 13.527 0.506 13.66 0.955 ;
      RECT 13.613 0.501 13.66 0.955 ;
      RECT 13.305 1.399 13.475 1.785 ;
      RECT 13.3 1.399 13.475 1.78 ;
      RECT 13.275 1.399 13.475 1.745 ;
      RECT 13.275 1.427 13.485 1.735 ;
      RECT 13.255 1.427 13.485 1.695 ;
      RECT 13.25 1.427 13.485 1.668 ;
      RECT 13.25 1.445 13.49 1.66 ;
      RECT 13.195 1.445 13.49 1.595 ;
      RECT 13.195 1.462 13.5 1.578 ;
      RECT 13.185 1.462 13.5 1.518 ;
      RECT 13.185 1.479 13.505 1.515 ;
      RECT 13.18 1.315 13.35 1.493 ;
      RECT 13.18 1.349 13.436 1.493 ;
      RECT 13.175 2.115 13.18 2.128 ;
      RECT 13.17 2.01 13.175 2.133 ;
      RECT 13.145 1.87 13.17 2.148 ;
      RECT 13.11 1.821 13.145 2.18 ;
      RECT 13.105 1.789 13.11 2.2 ;
      RECT 13.1 1.78 13.105 2.2 ;
      RECT 13.02 1.745 13.1 2.2 ;
      RECT 12.957 1.715 13.02 2.2 ;
      RECT 12.871 1.703 12.957 2.2 ;
      RECT 12.785 1.689 12.871 2.2 ;
      RECT 12.705 1.676 12.785 2.186 ;
      RECT 12.67 1.668 12.705 2.166 ;
      RECT 12.66 1.665 12.67 2.157 ;
      RECT 12.63 1.66 12.66 2.144 ;
      RECT 12.58 1.635 12.63 2.12 ;
      RECT 12.566 1.609 12.58 2.102 ;
      RECT 12.48 1.569 12.566 2.078 ;
      RECT 12.435 1.517 12.48 2.047 ;
      RECT 12.425 1.492 12.435 2.034 ;
      RECT 12.42 1.273 12.425 1.295 ;
      RECT 12.415 1.475 12.425 2.03 ;
      RECT 12.415 1.271 12.42 1.385 ;
      RECT 12.405 1.267 12.415 2.026 ;
      RECT 12.361 1.265 12.405 2.014 ;
      RECT 12.275 1.265 12.361 1.985 ;
      RECT 12.245 1.265 12.275 1.958 ;
      RECT 12.23 1.265 12.245 1.946 ;
      RECT 12.19 1.277 12.23 1.931 ;
      RECT 12.17 1.296 12.19 1.91 ;
      RECT 12.16 1.306 12.17 1.894 ;
      RECT 12.15 1.312 12.16 1.883 ;
      RECT 12.13 1.322 12.15 1.866 ;
      RECT 12.125 1.331 12.13 1.853 ;
      RECT 12.12 1.335 12.125 1.803 ;
      RECT 12.11 1.341 12.12 1.72 ;
      RECT 12.105 1.345 12.11 1.634 ;
      RECT 12.1 1.365 12.105 1.571 ;
      RECT 12.095 1.388 12.1 1.518 ;
      RECT 12.09 1.406 12.095 1.463 ;
      RECT 12.7 1.225 12.87 1.485 ;
      RECT 12.87 1.19 12.915 1.471 ;
      RECT 12.831 1.192 12.92 1.454 ;
      RECT 12.72 1.209 13.006 1.425 ;
      RECT 12.72 1.224 13.01 1.397 ;
      RECT 12.72 1.205 12.92 1.454 ;
      RECT 12.745 1.193 12.87 1.485 ;
      RECT 12.831 1.191 12.915 1.471 ;
      RECT 11.885 0.58 12.055 1.07 ;
      RECT 11.885 0.58 12.09 1.05 ;
      RECT 12.02 0.5 12.13 1.01 ;
      RECT 12.001 0.504 12.15 0.98 ;
      RECT 11.915 0.512 12.17 0.963 ;
      RECT 11.915 0.518 12.175 0.953 ;
      RECT 11.915 0.527 12.195 0.941 ;
      RECT 11.89 0.552 12.225 0.919 ;
      RECT 11.89 0.572 12.23 0.899 ;
      RECT 11.885 0.585 12.24 0.879 ;
      RECT 11.885 0.652 12.245 0.86 ;
      RECT 11.885 0.785 12.25 0.847 ;
      RECT 11.88 0.59 12.24 0.68 ;
      RECT 11.89 0.547 12.195 0.941 ;
      RECT 12.001 0.502 12.13 1.01 ;
      RECT 11.875 2.255 12.175 2.51 ;
      RECT 11.96 2.221 12.175 2.51 ;
      RECT 11.96 2.224 12.18 2.37 ;
      RECT 11.895 2.245 12.18 2.37 ;
      RECT 11.93 2.235 12.175 2.51 ;
      RECT 11.925 2.24 12.18 2.37 ;
      RECT 11.96 2.219 12.161 2.51 ;
      RECT 12.046 2.21 12.161 2.51 ;
      RECT 12.046 2.204 12.075 2.51 ;
      RECT 11.535 1.845 11.545 2.335 ;
      RECT 11.195 1.78 11.205 2.08 ;
      RECT 11.71 1.952 11.715 2.171 ;
      RECT 11.7 1.932 11.71 2.188 ;
      RECT 11.69 1.912 11.7 2.218 ;
      RECT 11.685 1.902 11.69 2.233 ;
      RECT 11.68 1.898 11.685 2.238 ;
      RECT 11.665 1.89 11.68 2.245 ;
      RECT 11.625 1.87 11.665 2.27 ;
      RECT 11.6 1.852 11.625 2.303 ;
      RECT 11.595 1.85 11.6 2.316 ;
      RECT 11.575 1.847 11.595 2.32 ;
      RECT 11.545 1.845 11.575 2.33 ;
      RECT 11.475 1.847 11.535 2.331 ;
      RECT 11.455 1.847 11.475 2.325 ;
      RECT 11.43 1.845 11.455 2.322 ;
      RECT 11.395 1.84 11.43 2.318 ;
      RECT 11.375 1.834 11.395 2.305 ;
      RECT 11.365 1.831 11.375 2.293 ;
      RECT 11.345 1.828 11.365 2.278 ;
      RECT 11.325 1.824 11.345 2.26 ;
      RECT 11.32 1.821 11.325 2.25 ;
      RECT 11.315 1.82 11.32 2.248 ;
      RECT 11.305 1.817 11.315 2.24 ;
      RECT 11.295 1.811 11.305 2.223 ;
      RECT 11.285 1.805 11.295 2.205 ;
      RECT 11.275 1.799 11.285 2.193 ;
      RECT 11.265 1.793 11.275 2.173 ;
      RECT 11.26 1.789 11.265 2.158 ;
      RECT 11.255 1.787 11.26 2.15 ;
      RECT 11.25 1.785 11.255 2.143 ;
      RECT 11.245 1.783 11.25 2.133 ;
      RECT 11.24 1.781 11.245 2.127 ;
      RECT 11.23 1.78 11.24 2.117 ;
      RECT 11.22 1.78 11.23 2.108 ;
      RECT 11.205 1.78 11.22 2.093 ;
      RECT 11.165 1.78 11.195 2.077 ;
      RECT 11.145 1.782 11.165 2.072 ;
      RECT 11.14 1.787 11.145 2.07 ;
      RECT 11.11 1.795 11.14 2.068 ;
      RECT 11.08 1.81 11.11 2.067 ;
      RECT 11.035 1.832 11.08 2.072 ;
      RECT 11.03 1.847 11.035 2.076 ;
      RECT 11.015 1.852 11.03 2.078 ;
      RECT 11.01 1.856 11.015 2.08 ;
      RECT 10.95 1.879 11.01 2.089 ;
      RECT 10.93 1.905 10.95 2.102 ;
      RECT 10.92 1.912 10.93 2.106 ;
      RECT 10.905 1.919 10.92 2.109 ;
      RECT 10.885 1.929 10.905 2.112 ;
      RECT 10.88 1.937 10.885 2.115 ;
      RECT 10.835 1.942 10.88 2.122 ;
      RECT 10.825 1.945 10.835 2.129 ;
      RECT 10.815 1.945 10.825 2.133 ;
      RECT 10.78 1.947 10.815 2.145 ;
      RECT 10.76 1.95 10.78 2.158 ;
      RECT 10.72 1.953 10.76 2.169 ;
      RECT 10.705 1.955 10.72 2.182 ;
      RECT 10.695 1.955 10.705 2.187 ;
      RECT 10.67 1.956 10.695 2.195 ;
      RECT 10.66 1.958 10.67 2.2 ;
      RECT 10.655 1.959 10.66 2.203 ;
      RECT 10.63 1.957 10.655 2.206 ;
      RECT 10.615 1.955 10.63 2.207 ;
      RECT 10.595 1.952 10.615 2.209 ;
      RECT 10.575 1.947 10.595 2.209 ;
      RECT 10.515 1.942 10.575 2.206 ;
      RECT 10.48 1.917 10.515 2.202 ;
      RECT 10.47 1.894 10.48 2.2 ;
      RECT 10.44 1.871 10.47 2.2 ;
      RECT 10.43 1.85 10.44 2.2 ;
      RECT 10.405 1.832 10.43 2.198 ;
      RECT 10.39 1.81 10.405 2.195 ;
      RECT 10.375 1.792 10.39 2.193 ;
      RECT 10.355 1.782 10.375 2.191 ;
      RECT 10.34 1.777 10.355 2.19 ;
      RECT 10.325 1.775 10.34 2.189 ;
      RECT 10.295 1.776 10.325 2.187 ;
      RECT 10.275 1.779 10.295 2.185 ;
      RECT 10.218 1.783 10.275 2.185 ;
      RECT 10.132 1.792 10.218 2.185 ;
      RECT 10.046 1.803 10.132 2.185 ;
      RECT 9.96 1.814 10.046 2.185 ;
      RECT 9.94 1.821 9.96 2.193 ;
      RECT 9.93 1.824 9.94 2.2 ;
      RECT 9.865 1.829 9.93 2.218 ;
      RECT 9.835 1.836 9.865 2.243 ;
      RECT 9.825 1.839 9.835 2.25 ;
      RECT 9.78 1.843 9.825 2.255 ;
      RECT 9.75 1.848 9.78 2.26 ;
      RECT 9.749 1.85 9.75 2.26 ;
      RECT 9.663 1.856 9.749 2.26 ;
      RECT 9.577 1.867 9.663 2.26 ;
      RECT 9.491 1.879 9.577 2.26 ;
      RECT 9.405 1.89 9.491 2.26 ;
      RECT 9.39 1.897 9.405 2.255 ;
      RECT 9.385 1.899 9.39 2.249 ;
      RECT 9.365 1.91 9.385 2.244 ;
      RECT 9.355 1.928 9.365 2.238 ;
      RECT 9.35 1.94 9.355 2.038 ;
      RECT 11.645 0.693 11.665 0.78 ;
      RECT 11.64 0.628 11.645 0.812 ;
      RECT 11.63 0.595 11.64 0.817 ;
      RECT 11.625 0.575 11.63 0.823 ;
      RECT 11.595 0.575 11.625 0.84 ;
      RECT 11.546 0.575 11.595 0.876 ;
      RECT 11.46 0.575 11.546 0.934 ;
      RECT 11.431 0.585 11.46 0.983 ;
      RECT 11.345 0.627 11.431 1.036 ;
      RECT 11.325 0.665 11.345 1.083 ;
      RECT 11.3 0.682 11.325 1.103 ;
      RECT 11.29 0.696 11.3 1.123 ;
      RECT 11.285 0.702 11.29 1.133 ;
      RECT 11.28 0.706 11.285 1.14 ;
      RECT 11.23 0.726 11.28 1.145 ;
      RECT 11.165 0.77 11.23 1.145 ;
      RECT 11.14 0.82 11.165 1.145 ;
      RECT 11.13 0.85 11.14 1.145 ;
      RECT 11.125 0.877 11.13 1.145 ;
      RECT 11.12 0.895 11.125 1.145 ;
      RECT 11.11 0.937 11.12 1.145 ;
      RECT 11.46 1.495 11.63 1.67 ;
      RECT 11.4 1.323 11.46 1.658 ;
      RECT 11.39 1.316 11.4 1.641 ;
      RECT 11.345 1.495 11.63 1.621 ;
      RECT 11.326 1.495 11.63 1.599 ;
      RECT 11.24 1.495 11.63 1.564 ;
      RECT 11.22 1.315 11.39 1.52 ;
      RECT 11.22 1.462 11.625 1.52 ;
      RECT 11.22 1.41 11.6 1.52 ;
      RECT 11.22 1.365 11.565 1.52 ;
      RECT 11.22 1.347 11.53 1.52 ;
      RECT 11.22 1.337 11.525 1.52 ;
      RECT 10.94 2.295 11.13 2.52 ;
      RECT 10.93 2.296 11.135 2.515 ;
      RECT 10.93 2.298 11.145 2.495 ;
      RECT 10.93 2.302 11.15 2.48 ;
      RECT 10.93 2.289 11.1 2.515 ;
      RECT 10.93 2.292 11.125 2.515 ;
      RECT 10.94 2.288 11.1 2.52 ;
      RECT 11.026 2.286 11.1 2.52 ;
      RECT 10.65 1.537 10.82 1.775 ;
      RECT 10.65 1.537 10.906 1.689 ;
      RECT 10.65 1.537 10.91 1.599 ;
      RECT 10.7 1.31 10.92 1.578 ;
      RECT 10.695 1.327 10.925 1.551 ;
      RECT 10.66 1.485 10.925 1.551 ;
      RECT 10.68 1.335 10.82 1.775 ;
      RECT 10.67 1.417 10.93 1.534 ;
      RECT 10.665 1.465 10.93 1.534 ;
      RECT 10.67 1.375 10.925 1.551 ;
      RECT 10.695 1.312 10.92 1.578 ;
      RECT 10.26 1.287 10.43 1.485 ;
      RECT 10.26 1.287 10.475 1.46 ;
      RECT 10.33 1.23 10.5 1.418 ;
      RECT 10.305 1.245 10.5 1.418 ;
      RECT 9.92 1.291 9.95 1.485 ;
      RECT 9.915 1.263 9.92 1.485 ;
      RECT 9.885 1.237 9.915 1.487 ;
      RECT 9.86 1.195 9.885 1.49 ;
      RECT 9.85 1.167 9.86 1.492 ;
      RECT 9.815 1.147 9.85 1.494 ;
      RECT 9.75 1.132 9.815 1.5 ;
      RECT 9.7 1.13 9.75 1.506 ;
      RECT 9.677 1.132 9.7 1.511 ;
      RECT 9.591 1.143 9.677 1.517 ;
      RECT 9.505 1.161 9.591 1.527 ;
      RECT 9.49 1.172 9.505 1.533 ;
      RECT 9.42 1.195 9.49 1.539 ;
      RECT 9.365 1.227 9.42 1.547 ;
      RECT 9.325 1.25 9.365 1.553 ;
      RECT 9.311 1.263 9.325 1.556 ;
      RECT 9.225 1.285 9.311 1.562 ;
      RECT 9.21 1.31 9.225 1.568 ;
      RECT 9.17 1.325 9.21 1.572 ;
      RECT 9.12 1.34 9.17 1.577 ;
      RECT 9.095 1.347 9.12 1.581 ;
      RECT 9.035 1.342 9.095 1.585 ;
      RECT 9.02 1.333 9.035 1.589 ;
      RECT 8.95 1.323 9.02 1.585 ;
      RECT 8.925 1.315 8.945 1.575 ;
      RECT 8.866 1.315 8.925 1.553 ;
      RECT 8.78 1.315 8.866 1.51 ;
      RECT 8.945 1.315 8.95 1.58 ;
      RECT 9.64 0.546 9.81 0.88 ;
      RECT 9.61 0.546 9.81 0.875 ;
      RECT 9.55 0.513 9.61 0.863 ;
      RECT 9.55 0.569 9.82 0.858 ;
      RECT 9.525 0.569 9.82 0.852 ;
      RECT 9.52 0.51 9.55 0.849 ;
      RECT 9.505 0.516 9.64 0.847 ;
      RECT 9.5 0.524 9.725 0.835 ;
      RECT 9.5 0.576 9.835 0.788 ;
      RECT 9.485 0.532 9.725 0.783 ;
      RECT 9.485 0.602 9.845 0.724 ;
      RECT 9.455 0.552 9.81 0.685 ;
      RECT 9.455 0.642 9.855 0.681 ;
      RECT 9.505 0.521 9.725 0.847 ;
      RECT 8.845 0.851 8.9 1.115 ;
      RECT 8.845 0.851 8.965 1.114 ;
      RECT 8.845 0.851 8.99 1.113 ;
      RECT 8.845 0.851 9.055 1.112 ;
      RECT 8.99 0.817 9.07 1.111 ;
      RECT 8.805 0.861 9.215 1.11 ;
      RECT 8.845 0.858 9.215 1.11 ;
      RECT 8.805 0.866 9.22 1.103 ;
      RECT 8.79 0.868 9.22 1.102 ;
      RECT 8.79 0.875 9.225 1.098 ;
      RECT 8.77 0.874 9.22 1.094 ;
      RECT 8.77 0.882 9.23 1.093 ;
      RECT 8.765 0.879 9.225 1.089 ;
      RECT 8.765 0.892 9.24 1.088 ;
      RECT 8.75 0.882 9.23 1.087 ;
      RECT 8.715 0.895 9.24 1.08 ;
      RECT 8.9 0.85 9.21 1.11 ;
      RECT 8.9 0.835 9.16 1.11 ;
      RECT 8.965 0.822 9.095 1.11 ;
      RECT 8.51 1.911 8.525 2.304 ;
      RECT 8.475 1.916 8.525 2.303 ;
      RECT 8.51 1.915 8.57 2.302 ;
      RECT 8.455 1.926 8.57 2.301 ;
      RECT 8.47 1.922 8.57 2.301 ;
      RECT 8.435 1.932 8.645 2.298 ;
      RECT 8.435 1.951 8.69 2.296 ;
      RECT 8.435 1.958 8.695 2.293 ;
      RECT 8.42 1.935 8.645 2.29 ;
      RECT 8.4 1.94 8.645 2.283 ;
      RECT 8.395 1.944 8.645 2.279 ;
      RECT 8.395 1.961 8.705 2.278 ;
      RECT 8.375 1.955 8.69 2.274 ;
      RECT 8.375 1.964 8.71 2.268 ;
      RECT 8.37 1.97 8.71 2.04 ;
      RECT 8.435 1.93 8.57 2.298 ;
      RECT 8.31 1.293 8.51 1.605 ;
      RECT 8.385 1.271 8.51 1.605 ;
      RECT 8.325 1.29 8.515 1.59 ;
      RECT 8.295 1.301 8.515 1.588 ;
      RECT 8.31 1.296 8.52 1.554 ;
      RECT 8.295 1.4 8.525 1.521 ;
      RECT 8.325 1.272 8.51 1.605 ;
      RECT 8.385 1.25 8.485 1.605 ;
      RECT 8.41 1.247 8.485 1.605 ;
      RECT 8.41 1.242 8.43 1.605 ;
      RECT 7.815 1.31 7.99 1.485 ;
      RECT 7.81 1.31 7.99 1.483 ;
      RECT 7.785 1.31 7.99 1.478 ;
      RECT 7.73 1.29 7.9 1.468 ;
      RECT 7.73 1.297 7.965 1.468 ;
      RECT 7.815 1.977 7.83 2.16 ;
      RECT 7.805 1.955 7.815 2.16 ;
      RECT 7.79 1.935 7.805 2.16 ;
      RECT 7.78 1.91 7.79 2.16 ;
      RECT 7.75 1.875 7.78 2.16 ;
      RECT 7.715 1.815 7.75 2.16 ;
      RECT 7.71 1.777 7.715 2.16 ;
      RECT 7.66 1.728 7.71 2.16 ;
      RECT 7.65 1.678 7.66 2.148 ;
      RECT 7.635 1.657 7.65 2.108 ;
      RECT 7.615 1.625 7.635 2.058 ;
      RECT 7.59 1.581 7.615 1.998 ;
      RECT 7.585 1.553 7.59 1.953 ;
      RECT 7.58 1.544 7.585 1.939 ;
      RECT 7.575 1.537 7.58 1.926 ;
      RECT 7.57 1.532 7.575 1.915 ;
      RECT 7.565 1.517 7.57 1.905 ;
      RECT 7.56 1.495 7.565 1.892 ;
      RECT 7.55 1.455 7.56 1.867 ;
      RECT 7.525 1.385 7.55 1.823 ;
      RECT 7.52 1.325 7.525 1.788 ;
      RECT 7.505 1.305 7.52 1.755 ;
      RECT 7.5 1.305 7.505 1.73 ;
      RECT 7.47 1.305 7.5 1.685 ;
      RECT 7.425 1.305 7.47 1.625 ;
      RECT 7.35 1.305 7.425 1.573 ;
      RECT 7.345 1.305 7.35 1.538 ;
      RECT 7.34 1.305 7.345 1.528 ;
      RECT 7.335 1.305 7.34 1.508 ;
      RECT 7.6 0.525 7.77 0.995 ;
      RECT 7.545 0.518 7.74 0.979 ;
      RECT 7.545 0.532 7.775 0.978 ;
      RECT 7.53 0.533 7.775 0.959 ;
      RECT 7.525 0.551 7.775 0.945 ;
      RECT 7.53 0.534 7.78 0.943 ;
      RECT 7.515 0.565 7.78 0.928 ;
      RECT 7.53 0.54 7.785 0.913 ;
      RECT 7.51 0.58 7.785 0.91 ;
      RECT 7.525 0.552 7.79 0.895 ;
      RECT 7.525 0.564 7.795 0.875 ;
      RECT 7.51 0.58 7.8 0.858 ;
      RECT 7.51 0.59 7.805 0.713 ;
      RECT 7.505 0.59 7.805 0.67 ;
      RECT 7.505 0.605 7.81 0.648 ;
      RECT 7.6 0.515 7.74 0.995 ;
      RECT 7.6 0.513 7.71 0.995 ;
      RECT 7.686 0.51 7.71 0.995 ;
      RECT 7.345 2.177 7.35 2.223 ;
      RECT 7.335 2.025 7.345 2.247 ;
      RECT 7.33 1.87 7.335 2.272 ;
      RECT 7.315 1.832 7.33 2.283 ;
      RECT 7.31 1.815 7.315 2.29 ;
      RECT 7.3 1.803 7.31 2.297 ;
      RECT 7.295 1.794 7.3 2.299 ;
      RECT 7.29 1.792 7.295 2.303 ;
      RECT 7.245 1.783 7.29 2.318 ;
      RECT 7.24 1.775 7.245 2.332 ;
      RECT 7.235 1.772 7.24 2.336 ;
      RECT 7.22 1.767 7.235 2.344 ;
      RECT 7.165 1.757 7.22 2.355 ;
      RECT 7.13 1.745 7.165 2.356 ;
      RECT 7.121 1.74 7.13 2.35 ;
      RECT 7.035 1.74 7.121 2.34 ;
      RECT 7.005 1.74 7.035 2.318 ;
      RECT 6.995 1.74 7 2.298 ;
      RECT 6.99 1.74 6.995 2.26 ;
      RECT 6.985 1.74 6.99 2.218 ;
      RECT 6.98 1.74 6.985 2.178 ;
      RECT 6.975 1.74 6.98 2.108 ;
      RECT 6.965 1.74 6.975 2.03 ;
      RECT 6.96 1.74 6.965 1.93 ;
      RECT 7 1.74 7.005 2.3 ;
      RECT 6.495 1.822 6.585 2.3 ;
      RECT 6.48 1.825 6.6 2.298 ;
      RECT 6.495 1.824 6.6 2.298 ;
      RECT 6.46 1.831 6.625 2.288 ;
      RECT 6.48 1.825 6.625 2.288 ;
      RECT 6.445 1.837 6.625 2.276 ;
      RECT 6.48 1.828 6.675 2.269 ;
      RECT 6.431 1.845 6.675 2.267 ;
      RECT 6.46 1.835 6.685 2.255 ;
      RECT 6.431 1.856 6.715 2.246 ;
      RECT 6.345 1.88 6.715 2.24 ;
      RECT 6.345 1.893 6.755 2.223 ;
      RECT 6.34 1.915 6.755 2.216 ;
      RECT 6.31 1.93 6.755 2.206 ;
      RECT 6.305 1.941 6.755 2.196 ;
      RECT 6.275 1.954 6.755 2.187 ;
      RECT 6.26 1.972 6.755 2.176 ;
      RECT 6.235 1.985 6.755 2.166 ;
      RECT 6.495 1.821 6.505 2.3 ;
      RECT 6.541 1.245 6.58 1.49 ;
      RECT 6.455 1.245 6.59 1.488 ;
      RECT 6.34 1.27 6.59 1.485 ;
      RECT 6.34 1.27 6.595 1.483 ;
      RECT 6.34 1.27 6.61 1.478 ;
      RECT 6.446 1.245 6.625 1.458 ;
      RECT 6.36 1.253 6.625 1.458 ;
      RECT 6.03 0.605 6.2 1.04 ;
      RECT 6.02 0.639 6.2 1.023 ;
      RECT 6.1 0.575 6.27 1.01 ;
      RECT 6.005 0.65 6.27 0.988 ;
      RECT 6.1 0.585 6.275 0.978 ;
      RECT 6.03 0.637 6.305 0.963 ;
      RECT 5.99 0.663 6.305 0.948 ;
      RECT 5.99 0.705 6.315 0.928 ;
      RECT 5.985 0.73 6.32 0.91 ;
      RECT 5.985 0.74 6.325 0.895 ;
      RECT 5.98 0.677 6.305 0.893 ;
      RECT 5.98 0.75 6.33 0.878 ;
      RECT 5.975 0.687 6.305 0.875 ;
      RECT 5.97 0.771 6.335 0.858 ;
      RECT 5.97 0.803 6.34 0.838 ;
      RECT 5.965 0.717 6.315 0.83 ;
      RECT 5.97 0.702 6.305 0.858 ;
      RECT 5.985 0.672 6.305 0.91 ;
      RECT 5.83 1.259 6.055 1.515 ;
      RECT 5.83 1.292 6.075 1.505 ;
      RECT 5.795 1.292 6.075 1.503 ;
      RECT 5.795 1.305 6.08 1.493 ;
      RECT 5.795 1.325 6.09 1.485 ;
      RECT 5.795 1.422 6.095 1.478 ;
      RECT 5.775 1.17 5.905 1.468 ;
      RECT 5.73 1.325 6.09 1.41 ;
      RECT 5.72 1.17 5.905 1.355 ;
      RECT 5.72 1.202 5.991 1.355 ;
      RECT 5.685 1.732 5.705 1.91 ;
      RECT 5.65 1.685 5.685 1.91 ;
      RECT 5.635 1.625 5.65 1.91 ;
      RECT 5.61 1.572 5.635 1.91 ;
      RECT 5.595 1.525 5.61 1.91 ;
      RECT 5.575 1.502 5.595 1.91 ;
      RECT 5.55 1.467 5.575 1.91 ;
      RECT 5.54 1.313 5.55 1.91 ;
      RECT 5.51 1.308 5.54 1.901 ;
      RECT 5.505 1.305 5.51 1.891 ;
      RECT 5.49 1.305 5.505 1.865 ;
      RECT 5.485 1.305 5.49 1.828 ;
      RECT 5.46 1.305 5.485 1.78 ;
      RECT 5.44 1.305 5.46 1.705 ;
      RECT 5.43 1.305 5.44 1.665 ;
      RECT 5.425 1.305 5.43 1.64 ;
      RECT 5.42 1.305 5.425 1.623 ;
      RECT 5.415 1.305 5.42 1.605 ;
      RECT 5.41 1.306 5.415 1.595 ;
      RECT 5.4 1.308 5.41 1.563 ;
      RECT 5.39 1.31 5.4 1.53 ;
      RECT 5.38 1.313 5.39 1.503 ;
      RECT 5.705 1.74 5.93 1.91 ;
      RECT 5.035 0.552 5.205 1.005 ;
      RECT 5.035 0.552 5.295 0.971 ;
      RECT 5.035 0.552 5.325 0.955 ;
      RECT 5.035 0.552 5.355 0.928 ;
      RECT 5.291 0.53 5.37 0.91 ;
      RECT 5.07 0.537 5.375 0.895 ;
      RECT 5.07 0.545 5.385 0.858 ;
      RECT 5.03 0.572 5.385 0.83 ;
      RECT 5.015 0.585 5.385 0.795 ;
      RECT 5.035 0.56 5.405 0.785 ;
      RECT 5.01 0.625 5.405 0.755 ;
      RECT 5.01 0.655 5.41 0.738 ;
      RECT 5.005 0.685 5.41 0.725 ;
      RECT 5.07 0.534 5.37 0.91 ;
      RECT 5.205 0.531 5.291 0.989 ;
      RECT 5.156 0.532 5.37 0.91 ;
      RECT 5.3 2.192 5.345 2.385 ;
      RECT 5.29 2.162 5.3 2.385 ;
      RECT 5.285 2.147 5.29 2.385 ;
      RECT 5.245 2.057 5.285 2.385 ;
      RECT 5.24 1.97 5.245 2.385 ;
      RECT 5.23 1.94 5.24 2.385 ;
      RECT 5.225 1.9 5.23 2.385 ;
      RECT 5.215 1.862 5.225 2.385 ;
      RECT 5.21 1.827 5.215 2.385 ;
      RECT 5.19 1.78 5.21 2.385 ;
      RECT 5.175 1.705 5.19 2.385 ;
      RECT 5.17 1.66 5.175 2.38 ;
      RECT 5.165 1.64 5.17 2.353 ;
      RECT 5.16 1.62 5.165 2.338 ;
      RECT 5.155 1.595 5.16 2.318 ;
      RECT 5.15 1.573 5.155 2.303 ;
      RECT 5.145 1.551 5.15 2.285 ;
      RECT 5.14 1.53 5.145 2.275 ;
      RECT 5.13 1.502 5.14 2.245 ;
      RECT 5.12 1.465 5.13 2.213 ;
      RECT 5.11 1.425 5.12 2.18 ;
      RECT 5.1 1.403 5.11 2.15 ;
      RECT 5.07 1.355 5.1 2.082 ;
      RECT 5.055 1.315 5.07 2.009 ;
      RECT 5.045 1.315 5.055 1.975 ;
      RECT 5.04 1.315 5.045 1.95 ;
      RECT 5.035 1.315 5.04 1.935 ;
      RECT 5.03 1.315 5.035 1.913 ;
      RECT 5.025 1.315 5.03 1.9 ;
      RECT 5.01 1.315 5.025 1.865 ;
      RECT 4.99 1.315 5.01 1.805 ;
      RECT 4.98 1.315 4.99 1.755 ;
      RECT 4.96 1.315 4.98 1.703 ;
      RECT 4.94 1.315 4.96 1.66 ;
      RECT 4.93 1.315 4.94 1.648 ;
      RECT 4.9 1.315 4.93 1.635 ;
      RECT 4.87 1.336 4.9 1.615 ;
      RECT 4.86 1.364 4.87 1.595 ;
      RECT 4.845 1.381 4.86 1.563 ;
      RECT 4.84 1.395 4.845 1.53 ;
      RECT 4.835 1.403 4.84 1.503 ;
      RECT 4.83 1.411 4.835 1.465 ;
      RECT 4.835 1.935 4.84 2.27 ;
      RECT 4.8 1.922 4.835 2.269 ;
      RECT 4.73 1.862 4.8 2.268 ;
      RECT 4.65 1.805 4.73 2.267 ;
      RECT 4.515 1.765 4.65 2.266 ;
      RECT 4.515 1.952 4.85 2.255 ;
      RECT 4.475 1.952 4.85 2.245 ;
      RECT 4.475 1.97 4.855 2.24 ;
      RECT 4.475 2.06 4.86 2.23 ;
      RECT 4.47 1.755 4.635 2.21 ;
      RECT 4.465 1.755 4.635 1.953 ;
      RECT 4.465 1.912 4.83 1.953 ;
      RECT 4.465 1.9 4.825 1.953 ;
      RECT 3.73 2.115 4.245 2.525 ;
      RECT 3.905 1.135 4.245 2.525 ;
      RECT 3.015 1.135 4.245 1.305 ;
      RECT 3.725 0.53 3.97 1.305 ;
      RECT 1.125 2.535 3.155 2.705 ;
      RECT 2.985 1.68 3.155 2.705 ;
      RECT 1.125 1.235 1.295 2.705 ;
      RECT 2.985 1.68 3.735 1.87 ;
      RECT 1.1 1.235 1.295 1.565 ;
      RECT 1.805 1.855 2.815 2.025 ;
      RECT 2.625 0.495 2.815 2.025 ;
      RECT 1.805 1.055 1.975 2.025 ;
      RECT 1.465 2.195 2.59 2.365 ;
      RECT 1.465 0.495 1.635 2.365 ;
      RECT 0.62 1.235 0.875 1.565 ;
      RECT 0.705 0.895 0.875 1.565 ;
      RECT 0.705 0.895 1.635 1.065 ;
      RECT 1.46 0.495 1.635 1.065 ;
      RECT 1.46 0.495 1.99 0.86 ;
      RECT 0.28 1.735 0.615 2.705 ;
      RECT 0.28 0.495 0.45 2.705 ;
      RECT 0.28 0.495 0.535 1.065 ;
      RECT -0.41 2.115 0.105 2.525 ;
      RECT -0.235 1.135 0.105 2.525 ;
      RECT -1.125 1.135 0.105 1.305 ;
      RECT -0.415 0.53 -0.17 1.305 ;
      RECT -3.015 2.535 -0.985 2.705 ;
      RECT -1.155 1.68 -0.985 2.705 ;
      RECT -3.015 1.235 -2.845 2.705 ;
      RECT -1.155 1.68 -0.405 1.87 ;
      RECT -3.04 1.235 -2.845 1.565 ;
      RECT -2.335 1.855 -1.325 2.025 ;
      RECT -1.515 0.495 -1.325 2.025 ;
      RECT -2.335 1.055 -2.165 2.025 ;
      RECT -2.675 2.195 -1.55 2.365 ;
      RECT -2.675 0.495 -2.505 2.365 ;
      RECT -3.52 1.235 -3.265 1.565 ;
      RECT -3.435 0.895 -3.265 1.565 ;
      RECT -3.435 0.895 -2.505 1.065 ;
      RECT -2.68 0.495 -2.505 1.065 ;
      RECT -2.68 0.495 -2.15 0.86 ;
      RECT -3.86 1.735 -3.525 2.705 ;
      RECT -3.86 0.495 -3.69 2.705 ;
      RECT -3.86 0.495 -3.605 1.065 ;
      RECT 135.725 1.315 136.055 1.555 ;
      RECT 132.965 1.315 133.295 1.555 ;
      RECT 130.495 0.495 130.77 1.655 ;
      RECT 126.36 0.495 126.635 1.655 ;
      RECT 108.13 1.315 108.46 1.555 ;
      RECT 105.37 1.315 105.7 1.555 ;
      RECT 102.9 0.495 103.175 1.655 ;
      RECT 98.765 0.495 99.04 1.655 ;
      RECT 80.535 1.315 80.865 1.555 ;
      RECT 77.775 1.315 78.105 1.555 ;
      RECT 75.305 0.495 75.58 1.655 ;
      RECT 71.17 0.495 71.445 1.655 ;
      RECT 52.94 1.315 53.27 1.555 ;
      RECT 50.18 1.315 50.51 1.555 ;
      RECT 47.71 0.495 47.985 1.655 ;
      RECT 43.575 0.495 43.85 1.655 ;
      RECT 25.345 1.315 25.675 1.555 ;
      RECT 22.585 1.315 22.915 1.555 ;
      RECT 20.115 0.495 20.39 1.655 ;
      RECT 15.98 0.495 16.255 1.655 ;
      RECT -1.96 0.495 -1.685 1.655 ;
  END
END sky130_osu_ring_oscillator_mpr2aa_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ca_8_b0r1
  CLASS CORE ;
  ORIGIN 4.14 -0.06 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ca_8_b0r1 -4.14 0.06 ;
  SIZE 94.215 BY 5.92 ;
  SYMMETRY X Y ;
  SITE b0r1_b0r2_HFix ;
  OBS
    LAYER met4 ;
      RECT 89.245 4.855 89.67 5.28 ;
      RECT -0.01 4.85 0.415 5.275 ;
      RECT -0.01 4.91 89.67 5.23 ;
      RECT -0.015 4.905 0.415 5.225 ;
      RECT 74.18 1.1 74.56 1.48 ;
      RECT 84.935 1.09 85.315 1.47 ;
      RECT 74.18 1.135 85.315 1.44 ;
      RECT 56.24 1.1 56.62 1.48 ;
      RECT 66.995 1.09 67.375 1.47 ;
      RECT 56.24 1.135 67.375 1.44 ;
      RECT 38.305 1.1 38.685 1.48 ;
      RECT 49.06 1.09 49.44 1.47 ;
      RECT 38.305 1.135 49.44 1.44 ;
      RECT 20.365 1.1 20.745 1.48 ;
      RECT 31.12 1.09 31.5 1.47 ;
      RECT 20.365 1.135 31.5 1.44 ;
      RECT 2.425 1.1 2.805 1.48 ;
      RECT 13.18 1.09 13.56 1.47 ;
      RECT 2.425 1.135 13.56 1.44 ;
    LAYER via3 ;
      RECT 89.36 4.97 89.56 5.17 ;
      RECT 85.025 1.18 85.225 1.38 ;
      RECT 74.27 1.19 74.47 1.39 ;
      RECT 67.085 1.18 67.285 1.38 ;
      RECT 56.33 1.19 56.53 1.39 ;
      RECT 49.15 1.18 49.35 1.38 ;
      RECT 38.395 1.19 38.595 1.39 ;
      RECT 31.21 1.18 31.41 1.38 ;
      RECT 20.455 1.19 20.655 1.39 ;
      RECT 13.27 1.18 13.47 1.38 ;
      RECT 2.515 1.19 2.715 1.39 ;
      RECT 0.105 4.965 0.305 5.165 ;
    LAYER met3 ;
      RECT 89.245 4.855 89.665 5.28 ;
      RECT 88.93 4.9 89.96 5.245 ;
      RECT 84.935 1.09 85.315 1.47 ;
      RECT 84.675 1.125 85.58 1.435 ;
      RECT 72.525 4.02 72.895 4.39 ;
      RECT 72.525 4.055 73.2 4.355 ;
      RECT 72.855 0.24 73.155 4.355 ;
      RECT 83.81 1.28 84.18 1.65 ;
      RECT 83.875 0.275 84.175 1.65 ;
      RECT 72.855 0.275 84.185 0.575 ;
      RECT 80.86 1.325 81.19 1.655 ;
      RECT 80.86 1.34 81.66 1.64 ;
      RECT 75.76 4.38 76.13 4.75 ;
      RECT 80.18 4.385 80.51 4.715 ;
      RECT 79.135 4.385 79.465 4.715 ;
      RECT 79.135 4.41 80.51 4.71 ;
      RECT 75.76 4.41 80.98 4.7 ;
      RECT 80.86 2.345 81.185 4.695 ;
      RECT 80.18 4.4 81.185 4.695 ;
      RECT 80.855 2.63 80.98 4.7 ;
      RECT 75.76 4.4 79.465 4.7 ;
      RECT 80.185 4.38 80.485 4.715 ;
      RECT 80.86 2.345 81.19 2.675 ;
      RECT 80.86 2.36 81.66 2.66 ;
      RECT 80.865 2.295 81.165 4.695 ;
      RECT 80.16 1.665 80.49 1.995 ;
      RECT 79.69 1.68 80.49 1.98 ;
      RECT 80.185 1.65 80.485 1.995 ;
      RECT 79.5 3.365 79.83 3.695 ;
      RECT 79.5 3.38 80.3 3.68 ;
      RECT 78.82 0.98 79.15 1.31 ;
      RECT 78.35 1 78.71 1.3 ;
      RECT 78.71 0.995 79.15 1.295 ;
      RECT 78.43 5.08 78.73 5.495 ;
      RECT 78.46 5.065 78.79 5.395 ;
      RECT 77.99 5.08 78.79 5.38 ;
      RECT 74.23 3.875 74.6 4.245 ;
      RECT 74.21 1.1 74.51 4.055 ;
      RECT 74.18 1.1 74.56 1.48 ;
      RECT 66.995 1.09 67.375 1.47 ;
      RECT 66.735 1.125 67.64 1.435 ;
      RECT 54.585 4.02 54.955 4.39 ;
      RECT 54.585 4.055 55.26 4.355 ;
      RECT 54.915 0.24 55.215 4.355 ;
      RECT 65.87 1.28 66.24 1.65 ;
      RECT 65.935 0.275 66.235 1.65 ;
      RECT 54.915 0.275 66.245 0.575 ;
      RECT 62.92 1.325 63.25 1.655 ;
      RECT 62.92 1.34 63.72 1.64 ;
      RECT 57.82 4.38 58.19 4.75 ;
      RECT 62.24 4.385 62.57 4.715 ;
      RECT 61.195 4.385 61.525 4.715 ;
      RECT 61.195 4.41 62.57 4.71 ;
      RECT 57.82 4.41 63.04 4.7 ;
      RECT 62.92 2.345 63.245 4.695 ;
      RECT 62.24 4.4 63.245 4.695 ;
      RECT 62.915 2.63 63.04 4.7 ;
      RECT 57.82 4.4 61.525 4.7 ;
      RECT 62.245 4.38 62.545 4.715 ;
      RECT 62.92 2.345 63.25 2.675 ;
      RECT 62.92 2.36 63.72 2.66 ;
      RECT 62.925 2.295 63.225 4.695 ;
      RECT 62.22 1.665 62.55 1.995 ;
      RECT 61.75 1.68 62.55 1.98 ;
      RECT 62.245 1.65 62.545 1.995 ;
      RECT 61.56 3.365 61.89 3.695 ;
      RECT 61.56 3.38 62.36 3.68 ;
      RECT 60.88 0.98 61.21 1.31 ;
      RECT 60.41 1 60.77 1.3 ;
      RECT 60.77 0.995 61.21 1.295 ;
      RECT 60.49 5.08 60.79 5.495 ;
      RECT 60.52 5.065 60.85 5.395 ;
      RECT 60.05 5.08 60.85 5.38 ;
      RECT 56.29 3.875 56.66 4.245 ;
      RECT 56.27 1.1 56.57 4.055 ;
      RECT 56.24 1.1 56.62 1.48 ;
      RECT 49.06 1.09 49.44 1.47 ;
      RECT 48.8 1.125 49.705 1.435 ;
      RECT 36.65 4.02 37.02 4.39 ;
      RECT 36.65 4.055 37.325 4.355 ;
      RECT 36.98 0.24 37.28 4.355 ;
      RECT 47.935 1.28 48.305 1.65 ;
      RECT 48 0.275 48.3 1.65 ;
      RECT 36.98 0.275 48.31 0.575 ;
      RECT 44.985 1.325 45.315 1.655 ;
      RECT 44.985 1.34 45.785 1.64 ;
      RECT 39.885 4.38 40.255 4.75 ;
      RECT 44.305 4.385 44.635 4.715 ;
      RECT 43.26 4.385 43.59 4.715 ;
      RECT 43.26 4.41 44.635 4.71 ;
      RECT 39.885 4.41 45.105 4.7 ;
      RECT 44.985 2.345 45.31 4.695 ;
      RECT 44.305 4.4 45.31 4.695 ;
      RECT 44.98 2.63 45.105 4.7 ;
      RECT 39.885 4.4 43.59 4.7 ;
      RECT 44.31 4.38 44.61 4.715 ;
      RECT 44.985 2.345 45.315 2.675 ;
      RECT 44.985 2.36 45.785 2.66 ;
      RECT 44.99 2.295 45.29 4.695 ;
      RECT 44.285 1.665 44.615 1.995 ;
      RECT 43.815 1.68 44.615 1.98 ;
      RECT 44.31 1.65 44.61 1.995 ;
      RECT 43.625 3.365 43.955 3.695 ;
      RECT 43.625 3.38 44.425 3.68 ;
      RECT 42.945 0.98 43.275 1.31 ;
      RECT 42.475 1 42.835 1.3 ;
      RECT 42.835 0.995 43.275 1.295 ;
      RECT 42.555 5.08 42.855 5.495 ;
      RECT 42.585 5.065 42.915 5.395 ;
      RECT 42.115 5.08 42.915 5.38 ;
      RECT 38.355 3.875 38.725 4.245 ;
      RECT 38.335 1.1 38.635 4.055 ;
      RECT 38.305 1.1 38.685 1.48 ;
      RECT 31.12 1.09 31.5 1.47 ;
      RECT 30.86 1.125 31.765 1.435 ;
      RECT 18.71 4.02 19.08 4.39 ;
      RECT 18.71 4.055 19.385 4.355 ;
      RECT 19.04 0.24 19.34 4.355 ;
      RECT 29.995 1.28 30.365 1.65 ;
      RECT 30.06 0.275 30.36 1.65 ;
      RECT 19.04 0.275 30.37 0.575 ;
      RECT 27.045 1.325 27.375 1.655 ;
      RECT 27.045 1.34 27.845 1.64 ;
      RECT 21.945 4.38 22.315 4.75 ;
      RECT 26.365 4.385 26.695 4.715 ;
      RECT 25.32 4.385 25.65 4.715 ;
      RECT 25.32 4.41 26.695 4.71 ;
      RECT 21.945 4.41 27.165 4.7 ;
      RECT 27.045 2.345 27.37 4.695 ;
      RECT 26.365 4.4 27.37 4.695 ;
      RECT 27.04 2.63 27.165 4.7 ;
      RECT 21.945 4.4 25.65 4.7 ;
      RECT 26.37 4.38 26.67 4.715 ;
      RECT 27.045 2.345 27.375 2.675 ;
      RECT 27.045 2.36 27.845 2.66 ;
      RECT 27.05 2.295 27.35 4.695 ;
      RECT 26.345 1.665 26.675 1.995 ;
      RECT 25.875 1.68 26.675 1.98 ;
      RECT 26.37 1.65 26.67 1.995 ;
      RECT 25.685 3.365 26.015 3.695 ;
      RECT 25.685 3.38 26.485 3.68 ;
      RECT 25.005 0.98 25.335 1.31 ;
      RECT 24.535 1 24.895 1.3 ;
      RECT 24.895 0.995 25.335 1.295 ;
      RECT 24.615 5.08 24.915 5.495 ;
      RECT 24.645 5.065 24.975 5.395 ;
      RECT 24.175 5.08 24.975 5.38 ;
      RECT 20.415 3.875 20.785 4.245 ;
      RECT 20.395 1.1 20.695 4.055 ;
      RECT 20.365 1.1 20.745 1.48 ;
      RECT 13.18 1.09 13.56 1.47 ;
      RECT 12.92 1.125 13.825 1.435 ;
      RECT 0.77 4.02 1.14 4.39 ;
      RECT 0.77 4.055 1.445 4.355 ;
      RECT 1.1 0.24 1.4 4.355 ;
      RECT 12.055 1.28 12.425 1.65 ;
      RECT 12.12 0.275 12.42 1.65 ;
      RECT 1.1 0.275 12.43 0.575 ;
      RECT 9.105 1.325 9.435 1.655 ;
      RECT 9.105 1.34 9.905 1.64 ;
      RECT 4.005 4.38 4.375 4.75 ;
      RECT 8.425 4.385 8.755 4.715 ;
      RECT 7.38 4.385 7.71 4.715 ;
      RECT 7.38 4.41 8.755 4.71 ;
      RECT 4.005 4.41 9.225 4.7 ;
      RECT 9.105 2.345 9.43 4.695 ;
      RECT 8.425 4.4 9.43 4.695 ;
      RECT 9.1 2.63 9.225 4.7 ;
      RECT 4.005 4.4 7.71 4.7 ;
      RECT 8.43 4.38 8.73 4.715 ;
      RECT 9.105 2.345 9.435 2.675 ;
      RECT 9.105 2.36 9.905 2.66 ;
      RECT 9.11 2.295 9.41 4.695 ;
      RECT 8.405 1.665 8.735 1.995 ;
      RECT 7.935 1.68 8.735 1.98 ;
      RECT 8.43 1.65 8.73 1.995 ;
      RECT 7.745 3.365 8.075 3.695 ;
      RECT 7.745 3.38 8.545 3.68 ;
      RECT 7.065 0.98 7.395 1.31 ;
      RECT 6.595 1 6.955 1.3 ;
      RECT 6.955 0.995 7.395 1.295 ;
      RECT 6.675 5.08 6.975 5.495 ;
      RECT 6.705 5.065 7.035 5.395 ;
      RECT 6.235 5.08 7.035 5.38 ;
      RECT 2.475 3.875 2.845 4.245 ;
      RECT 2.455 1.1 2.755 4.055 ;
      RECT 2.425 1.1 2.805 1.48 ;
      RECT -0.01 4.85 0.41 5.275 ;
      RECT -0.325 4.895 0.705 5.24 ;
    LAYER via2 ;
      RECT 89.36 4.97 89.56 5.17 ;
      RECT 85.03 1.18 85.23 1.38 ;
      RECT 83.895 1.365 84.095 1.565 ;
      RECT 80.925 1.39 81.125 1.59 ;
      RECT 80.925 2.41 81.125 2.61 ;
      RECT 80.245 4.45 80.445 4.65 ;
      RECT 80.225 1.73 80.425 1.93 ;
      RECT 79.565 3.43 79.765 3.63 ;
      RECT 79.2 4.45 79.4 4.65 ;
      RECT 78.885 1.045 79.085 1.245 ;
      RECT 78.525 5.13 78.725 5.33 ;
      RECT 75.845 4.465 76.045 4.665 ;
      RECT 74.315 3.96 74.515 4.16 ;
      RECT 72.61 4.105 72.81 4.305 ;
      RECT 67.09 1.18 67.29 1.38 ;
      RECT 65.955 1.365 66.155 1.565 ;
      RECT 62.985 1.39 63.185 1.59 ;
      RECT 62.985 2.41 63.185 2.61 ;
      RECT 62.305 4.45 62.505 4.65 ;
      RECT 62.285 1.73 62.485 1.93 ;
      RECT 61.625 3.43 61.825 3.63 ;
      RECT 61.26 4.45 61.46 4.65 ;
      RECT 60.945 1.045 61.145 1.245 ;
      RECT 60.585 5.13 60.785 5.33 ;
      RECT 57.905 4.465 58.105 4.665 ;
      RECT 56.375 3.96 56.575 4.16 ;
      RECT 54.67 4.105 54.87 4.305 ;
      RECT 49.155 1.18 49.355 1.38 ;
      RECT 48.02 1.365 48.22 1.565 ;
      RECT 45.05 1.39 45.25 1.59 ;
      RECT 45.05 2.41 45.25 2.61 ;
      RECT 44.37 4.45 44.57 4.65 ;
      RECT 44.35 1.73 44.55 1.93 ;
      RECT 43.69 3.43 43.89 3.63 ;
      RECT 43.325 4.45 43.525 4.65 ;
      RECT 43.01 1.045 43.21 1.245 ;
      RECT 42.65 5.13 42.85 5.33 ;
      RECT 39.97 4.465 40.17 4.665 ;
      RECT 38.44 3.96 38.64 4.16 ;
      RECT 36.735 4.105 36.935 4.305 ;
      RECT 31.215 1.18 31.415 1.38 ;
      RECT 30.08 1.365 30.28 1.565 ;
      RECT 27.11 1.39 27.31 1.59 ;
      RECT 27.11 2.41 27.31 2.61 ;
      RECT 26.43 4.45 26.63 4.65 ;
      RECT 26.41 1.73 26.61 1.93 ;
      RECT 25.75 3.43 25.95 3.63 ;
      RECT 25.385 4.45 25.585 4.65 ;
      RECT 25.07 1.045 25.27 1.245 ;
      RECT 24.71 5.13 24.91 5.33 ;
      RECT 22.03 4.465 22.23 4.665 ;
      RECT 20.5 3.96 20.7 4.16 ;
      RECT 18.795 4.105 18.995 4.305 ;
      RECT 13.275 1.18 13.475 1.38 ;
      RECT 12.14 1.365 12.34 1.565 ;
      RECT 9.17 1.39 9.37 1.59 ;
      RECT 9.17 2.41 9.37 2.61 ;
      RECT 8.49 4.45 8.69 4.65 ;
      RECT 8.47 1.73 8.67 1.93 ;
      RECT 7.81 3.43 8.01 3.63 ;
      RECT 7.445 4.45 7.645 4.65 ;
      RECT 7.13 1.045 7.33 1.245 ;
      RECT 6.77 5.13 6.97 5.33 ;
      RECT 4.09 4.465 4.29 4.665 ;
      RECT 2.56 3.96 2.76 4.16 ;
      RECT 0.855 4.105 1.055 4.305 ;
      RECT 0.105 4.965 0.305 5.165 ;
    LAYER met2 ;
      RECT 84.945 4.575 85.285 4.915 ;
      RECT 84.945 4.705 86.22 4.895 ;
      RECT 86.03 3.47 86.22 4.895 ;
      RECT 85.56 3.47 86.22 3.66 ;
      RECT 85.56 1.7 85.75 3.66 ;
      RECT 85.41 1.7 85.75 2.04 ;
      RECT 81.95 1.7 82.29 2.04 ;
      RECT 82.24 0.67 82.38 1.995 ;
      RECT 85.605 0.67 85.745 3.66 ;
      RECT 82.24 0.67 85.745 0.81 ;
      RECT 85.365 3.97 85.705 4.31 ;
      RECT 84.59 3.97 85.705 4.14 ;
      RECT 84.59 1.2 84.76 4.14 ;
      RECT 84.945 1.095 85.315 1.465 ;
      RECT 84.59 1.2 85.315 1.37 ;
      RECT 83.81 4.415 84.15 4.755 ;
      RECT 83.92 1.28 84.09 4.755 ;
      RECT 83.81 1.28 84.18 1.65 ;
      RECT 82.585 3.37 82.845 3.69 ;
      RECT 82.645 1.33 82.785 3.69 ;
      RECT 82.585 1.33 82.845 1.65 ;
      RECT 81.565 4.39 81.825 4.71 ;
      RECT 80.945 4.48 81.825 4.62 ;
      RECT 80.945 2.325 81.085 4.62 ;
      RECT 80.885 2.325 81.165 2.695 ;
      RECT 80.205 4.365 80.485 4.735 ;
      RECT 80.265 2.44 80.405 4.735 ;
      RECT 80.265 2.44 80.745 2.58 ;
      RECT 80.605 0.65 80.745 2.58 ;
      RECT 80.545 0.65 80.805 0.97 ;
      RECT 79.525 3.345 79.805 3.715 ;
      RECT 79.585 0.99 79.725 3.715 ;
      RECT 79.525 0.99 79.785 1.31 ;
      RECT 79.16 4.365 79.44 4.735 ;
      RECT 79.16 4.39 79.445 4.71 ;
      RECT 67.005 4.575 67.345 4.915 ;
      RECT 67.005 4.705 68.28 4.895 ;
      RECT 68.09 3.47 68.28 4.895 ;
      RECT 67.62 3.47 68.28 3.66 ;
      RECT 67.62 1.7 67.81 3.66 ;
      RECT 67.47 1.7 67.81 2.04 ;
      RECT 64.01 1.7 64.35 2.04 ;
      RECT 64.3 0.67 64.44 1.995 ;
      RECT 67.665 0.67 67.805 3.66 ;
      RECT 64.3 0.67 67.805 0.81 ;
      RECT 67.425 3.97 67.765 4.31 ;
      RECT 66.65 3.97 67.765 4.14 ;
      RECT 66.65 1.2 66.82 4.14 ;
      RECT 67.005 1.095 67.375 1.465 ;
      RECT 66.65 1.2 67.375 1.37 ;
      RECT 65.87 4.415 66.21 4.755 ;
      RECT 65.98 1.28 66.15 4.755 ;
      RECT 65.87 1.28 66.24 1.65 ;
      RECT 64.645 3.37 64.905 3.69 ;
      RECT 64.705 1.33 64.845 3.69 ;
      RECT 64.645 1.33 64.905 1.65 ;
      RECT 63.625 4.39 63.885 4.71 ;
      RECT 63.005 4.48 63.885 4.62 ;
      RECT 63.005 2.325 63.145 4.62 ;
      RECT 62.945 2.325 63.225 2.695 ;
      RECT 62.265 4.365 62.545 4.735 ;
      RECT 62.325 2.44 62.465 4.735 ;
      RECT 62.325 2.44 62.805 2.58 ;
      RECT 62.665 0.65 62.805 2.58 ;
      RECT 62.605 0.65 62.865 0.97 ;
      RECT 61.585 3.345 61.865 3.715 ;
      RECT 61.645 0.99 61.785 3.715 ;
      RECT 61.585 0.99 61.845 1.31 ;
      RECT 61.22 4.365 61.5 4.735 ;
      RECT 61.22 4.39 61.505 4.71 ;
      RECT 49.07 4.575 49.41 4.915 ;
      RECT 49.07 4.705 50.345 4.895 ;
      RECT 50.155 3.47 50.345 4.895 ;
      RECT 49.685 3.47 50.345 3.66 ;
      RECT 49.685 1.7 49.875 3.66 ;
      RECT 49.535 1.7 49.875 2.04 ;
      RECT 46.075 1.7 46.415 2.04 ;
      RECT 46.365 0.67 46.505 1.995 ;
      RECT 49.73 0.67 49.87 3.66 ;
      RECT 46.365 0.67 49.87 0.81 ;
      RECT 49.49 3.97 49.83 4.31 ;
      RECT 48.715 3.97 49.83 4.14 ;
      RECT 48.715 1.2 48.885 4.14 ;
      RECT 49.07 1.095 49.44 1.465 ;
      RECT 48.715 1.2 49.44 1.37 ;
      RECT 47.935 4.415 48.275 4.755 ;
      RECT 48.045 1.28 48.215 4.755 ;
      RECT 47.935 1.28 48.305 1.65 ;
      RECT 46.71 3.37 46.97 3.69 ;
      RECT 46.77 1.33 46.91 3.69 ;
      RECT 46.71 1.33 46.97 1.65 ;
      RECT 45.69 4.39 45.95 4.71 ;
      RECT 45.07 4.48 45.95 4.62 ;
      RECT 45.07 2.325 45.21 4.62 ;
      RECT 45.01 2.325 45.29 2.695 ;
      RECT 44.33 4.365 44.61 4.735 ;
      RECT 44.39 2.44 44.53 4.735 ;
      RECT 44.39 2.44 44.87 2.58 ;
      RECT 44.73 0.65 44.87 2.58 ;
      RECT 44.67 0.65 44.93 0.97 ;
      RECT 43.65 3.345 43.93 3.715 ;
      RECT 43.71 0.99 43.85 3.715 ;
      RECT 43.65 0.99 43.91 1.31 ;
      RECT 43.285 4.365 43.565 4.735 ;
      RECT 43.285 4.39 43.57 4.71 ;
      RECT 31.13 4.575 31.47 4.915 ;
      RECT 31.13 4.705 32.405 4.895 ;
      RECT 32.215 3.47 32.405 4.895 ;
      RECT 31.745 3.47 32.405 3.66 ;
      RECT 31.745 1.7 31.935 3.66 ;
      RECT 31.595 1.7 31.935 2.04 ;
      RECT 28.135 1.7 28.475 2.04 ;
      RECT 28.425 0.67 28.565 1.995 ;
      RECT 31.79 0.67 31.93 3.66 ;
      RECT 28.425 0.67 31.93 0.81 ;
      RECT 31.55 3.97 31.89 4.31 ;
      RECT 30.775 3.97 31.89 4.14 ;
      RECT 30.775 1.2 30.945 4.14 ;
      RECT 31.13 1.095 31.5 1.465 ;
      RECT 30.775 1.2 31.5 1.37 ;
      RECT 29.995 4.415 30.335 4.755 ;
      RECT 30.105 1.28 30.275 4.755 ;
      RECT 29.995 1.28 30.365 1.65 ;
      RECT 28.77 3.37 29.03 3.69 ;
      RECT 28.83 1.33 28.97 3.69 ;
      RECT 28.77 1.33 29.03 1.65 ;
      RECT 27.75 4.39 28.01 4.71 ;
      RECT 27.13 4.48 28.01 4.62 ;
      RECT 27.13 2.325 27.27 4.62 ;
      RECT 27.07 2.325 27.35 2.695 ;
      RECT 26.39 4.365 26.67 4.735 ;
      RECT 26.45 2.44 26.59 4.735 ;
      RECT 26.45 2.44 26.93 2.58 ;
      RECT 26.79 0.65 26.93 2.58 ;
      RECT 26.73 0.65 26.99 0.97 ;
      RECT 25.71 3.345 25.99 3.715 ;
      RECT 25.77 0.99 25.91 3.715 ;
      RECT 25.71 0.99 25.97 1.31 ;
      RECT 25.345 4.365 25.625 4.735 ;
      RECT 25.345 4.39 25.63 4.71 ;
      RECT 13.19 4.575 13.53 4.915 ;
      RECT 13.19 4.705 14.465 4.895 ;
      RECT 14.275 3.47 14.465 4.895 ;
      RECT 13.805 3.47 14.465 3.66 ;
      RECT 13.805 1.7 13.995 3.66 ;
      RECT 13.655 1.7 13.995 2.04 ;
      RECT 10.195 1.7 10.535 2.04 ;
      RECT 10.485 0.67 10.625 1.995 ;
      RECT 13.85 0.67 13.99 3.66 ;
      RECT 10.485 0.67 13.99 0.81 ;
      RECT 13.61 3.97 13.95 4.31 ;
      RECT 12.835 3.97 13.95 4.14 ;
      RECT 12.835 1.2 13.005 4.14 ;
      RECT 13.19 1.095 13.56 1.465 ;
      RECT 12.835 1.2 13.56 1.37 ;
      RECT 12.055 4.415 12.395 4.755 ;
      RECT 12.165 1.28 12.335 4.755 ;
      RECT 12.055 1.28 12.425 1.65 ;
      RECT 10.83 3.37 11.09 3.69 ;
      RECT 10.89 1.33 11.03 3.69 ;
      RECT 10.83 1.33 11.09 1.65 ;
      RECT 9.81 4.39 10.07 4.71 ;
      RECT 9.19 4.48 10.07 4.62 ;
      RECT 9.19 2.325 9.33 4.62 ;
      RECT 9.13 2.325 9.41 2.695 ;
      RECT 8.45 4.365 8.73 4.735 ;
      RECT 8.51 2.44 8.65 4.735 ;
      RECT 8.51 2.44 8.99 2.58 ;
      RECT 8.85 0.65 8.99 2.58 ;
      RECT 8.79 0.65 9.05 0.97 ;
      RECT 7.77 3.345 8.05 3.715 ;
      RECT 7.83 0.99 7.97 3.715 ;
      RECT 7.77 0.99 8.03 1.31 ;
      RECT 7.405 4.365 7.685 4.735 ;
      RECT 7.405 4.39 7.69 4.71 ;
      RECT 2.475 3.875 2.845 4.245 ;
      RECT -3.885 3.55 -3.505 3.93 ;
      RECT 2.52 3.55 2.66 4.245 ;
      RECT -3.885 3.55 2.66 3.69 ;
      RECT 89.24 4.86 89.67 5.28 ;
      RECT 80.885 1.305 81.165 1.675 ;
      RECT 80.185 1.645 80.465 2.015 ;
      RECT 78.845 0.96 79.125 1.33 ;
      RECT 78.485 5.045 78.765 5.415 ;
      RECT 75.76 4.38 76.13 4.75 ;
      RECT 74.23 3.875 74.6 4.245 ;
      RECT 72.525 4.02 72.895 4.39 ;
      RECT 62.945 1.305 63.225 1.675 ;
      RECT 62.245 1.645 62.525 2.015 ;
      RECT 60.905 0.96 61.185 1.33 ;
      RECT 60.545 5.045 60.825 5.415 ;
      RECT 57.82 4.38 58.19 4.75 ;
      RECT 56.29 3.875 56.66 4.245 ;
      RECT 54.585 4.02 54.955 4.39 ;
      RECT 45.01 1.305 45.29 1.675 ;
      RECT 44.31 1.645 44.59 2.015 ;
      RECT 42.97 0.96 43.25 1.33 ;
      RECT 42.61 5.045 42.89 5.415 ;
      RECT 39.885 4.38 40.255 4.75 ;
      RECT 38.355 3.875 38.725 4.245 ;
      RECT 36.65 4.02 37.02 4.39 ;
      RECT 27.07 1.305 27.35 1.675 ;
      RECT 26.37 1.645 26.65 2.015 ;
      RECT 25.03 0.96 25.31 1.33 ;
      RECT 24.67 5.045 24.95 5.415 ;
      RECT 21.945 4.38 22.315 4.75 ;
      RECT 20.415 3.875 20.785 4.245 ;
      RECT 18.71 4.02 19.08 4.39 ;
      RECT 9.13 1.305 9.41 1.675 ;
      RECT 8.43 1.645 8.71 2.015 ;
      RECT 7.09 0.96 7.37 1.33 ;
      RECT 6.73 5.045 7.01 5.415 ;
      RECT 4.005 4.38 4.375 4.75 ;
      RECT 0.77 4.02 1.14 4.39 ;
      RECT -0.015 4.855 0.415 5.275 ;
    LAYER via1 ;
      RECT 89.385 4.995 89.535 5.145 ;
      RECT 85.505 1.795 85.655 1.945 ;
      RECT 85.46 4.065 85.61 4.215 ;
      RECT 85.055 1.205 85.205 1.355 ;
      RECT 85.04 4.67 85.19 4.82 ;
      RECT 83.91 1.38 84.06 1.53 ;
      RECT 83.905 4.51 84.055 4.66 ;
      RECT 82.64 1.415 82.79 1.565 ;
      RECT 82.64 3.455 82.79 3.605 ;
      RECT 82.045 1.795 82.195 1.945 ;
      RECT 81.62 4.475 81.77 4.625 ;
      RECT 80.94 1.415 81.09 1.565 ;
      RECT 80.94 2.435 81.09 2.585 ;
      RECT 80.6 0.735 80.75 0.885 ;
      RECT 80.26 1.755 80.41 1.905 ;
      RECT 80.26 4.475 80.41 4.625 ;
      RECT 79.58 1.075 79.73 1.225 ;
      RECT 79.58 3.455 79.73 3.605 ;
      RECT 79.24 4.475 79.39 4.625 ;
      RECT 78.9 1.07 79.05 1.22 ;
      RECT 78.56 5.155 78.71 5.305 ;
      RECT 75.87 4.49 76.02 4.64 ;
      RECT 74.34 3.985 74.49 4.135 ;
      RECT 72.635 4.13 72.785 4.28 ;
      RECT 67.565 1.795 67.715 1.945 ;
      RECT 67.52 4.065 67.67 4.215 ;
      RECT 67.115 1.205 67.265 1.355 ;
      RECT 67.1 4.67 67.25 4.82 ;
      RECT 65.97 1.38 66.12 1.53 ;
      RECT 65.965 4.51 66.115 4.66 ;
      RECT 64.7 1.415 64.85 1.565 ;
      RECT 64.7 3.455 64.85 3.605 ;
      RECT 64.105 1.795 64.255 1.945 ;
      RECT 63.68 4.475 63.83 4.625 ;
      RECT 63 1.415 63.15 1.565 ;
      RECT 63 2.435 63.15 2.585 ;
      RECT 62.66 0.735 62.81 0.885 ;
      RECT 62.32 1.755 62.47 1.905 ;
      RECT 62.32 4.475 62.47 4.625 ;
      RECT 61.64 1.075 61.79 1.225 ;
      RECT 61.64 3.455 61.79 3.605 ;
      RECT 61.3 4.475 61.45 4.625 ;
      RECT 60.96 1.07 61.11 1.22 ;
      RECT 60.62 5.155 60.77 5.305 ;
      RECT 57.93 4.49 58.08 4.64 ;
      RECT 56.4 3.985 56.55 4.135 ;
      RECT 54.695 4.13 54.845 4.28 ;
      RECT 49.63 1.795 49.78 1.945 ;
      RECT 49.585 4.065 49.735 4.215 ;
      RECT 49.18 1.205 49.33 1.355 ;
      RECT 49.165 4.67 49.315 4.82 ;
      RECT 48.035 1.38 48.185 1.53 ;
      RECT 48.03 4.51 48.18 4.66 ;
      RECT 46.765 1.415 46.915 1.565 ;
      RECT 46.765 3.455 46.915 3.605 ;
      RECT 46.17 1.795 46.32 1.945 ;
      RECT 45.745 4.475 45.895 4.625 ;
      RECT 45.065 1.415 45.215 1.565 ;
      RECT 45.065 2.435 45.215 2.585 ;
      RECT 44.725 0.735 44.875 0.885 ;
      RECT 44.385 1.755 44.535 1.905 ;
      RECT 44.385 4.475 44.535 4.625 ;
      RECT 43.705 1.075 43.855 1.225 ;
      RECT 43.705 3.455 43.855 3.605 ;
      RECT 43.365 4.475 43.515 4.625 ;
      RECT 43.025 1.07 43.175 1.22 ;
      RECT 42.685 5.155 42.835 5.305 ;
      RECT 39.995 4.49 40.145 4.64 ;
      RECT 38.465 3.985 38.615 4.135 ;
      RECT 36.76 4.13 36.91 4.28 ;
      RECT 31.69 1.795 31.84 1.945 ;
      RECT 31.645 4.065 31.795 4.215 ;
      RECT 31.24 1.205 31.39 1.355 ;
      RECT 31.225 4.67 31.375 4.82 ;
      RECT 30.095 1.38 30.245 1.53 ;
      RECT 30.09 4.51 30.24 4.66 ;
      RECT 28.825 1.415 28.975 1.565 ;
      RECT 28.825 3.455 28.975 3.605 ;
      RECT 28.23 1.795 28.38 1.945 ;
      RECT 27.805 4.475 27.955 4.625 ;
      RECT 27.125 1.415 27.275 1.565 ;
      RECT 27.125 2.435 27.275 2.585 ;
      RECT 26.785 0.735 26.935 0.885 ;
      RECT 26.445 1.755 26.595 1.905 ;
      RECT 26.445 4.475 26.595 4.625 ;
      RECT 25.765 1.075 25.915 1.225 ;
      RECT 25.765 3.455 25.915 3.605 ;
      RECT 25.425 4.475 25.575 4.625 ;
      RECT 25.085 1.07 25.235 1.22 ;
      RECT 24.745 5.155 24.895 5.305 ;
      RECT 22.055 4.49 22.205 4.64 ;
      RECT 20.525 3.985 20.675 4.135 ;
      RECT 18.82 4.13 18.97 4.28 ;
      RECT 13.75 1.795 13.9 1.945 ;
      RECT 13.705 4.065 13.855 4.215 ;
      RECT 13.3 1.205 13.45 1.355 ;
      RECT 13.285 4.67 13.435 4.82 ;
      RECT 12.155 1.38 12.305 1.53 ;
      RECT 12.15 4.51 12.3 4.66 ;
      RECT 10.885 1.415 11.035 1.565 ;
      RECT 10.885 3.455 11.035 3.605 ;
      RECT 10.29 1.795 10.44 1.945 ;
      RECT 9.865 4.475 10.015 4.625 ;
      RECT 9.185 1.415 9.335 1.565 ;
      RECT 9.185 2.435 9.335 2.585 ;
      RECT 8.845 0.735 8.995 0.885 ;
      RECT 8.505 1.755 8.655 1.905 ;
      RECT 8.505 4.475 8.655 4.625 ;
      RECT 7.825 1.075 7.975 1.225 ;
      RECT 7.825 3.455 7.975 3.605 ;
      RECT 7.485 4.475 7.635 4.625 ;
      RECT 7.145 1.07 7.295 1.22 ;
      RECT 6.805 5.155 6.955 5.305 ;
      RECT 4.115 4.49 4.265 4.64 ;
      RECT 2.585 3.985 2.735 4.135 ;
      RECT 0.88 4.13 1.03 4.28 ;
      RECT 0.13 4.99 0.28 5.14 ;
      RECT -3.77 3.665 -3.62 3.815 ;
    LAYER met1 ;
      RECT -1.51 2.78 -1.32 4.365 ;
      RECT -1.53 4.07 -1.29 4.325 ;
      RECT -3.95 2.78 89.885 3.26 ;
      RECT -3.95 5.5 89.885 5.98 ;
      RECT 78.515 5.1 78.76 5.98 ;
      RECT 60.575 5.1 60.82 5.98 ;
      RECT 42.64 5.1 42.885 5.98 ;
      RECT 24.7 5.1 24.945 5.98 ;
      RECT 6.76 5.1 7.005 5.98 ;
      RECT 78.475 5.1 78.795 5.36 ;
      RECT 60.535 5.1 60.855 5.36 ;
      RECT 42.6 5.1 42.92 5.36 ;
      RECT 24.66 5.1 24.98 5.36 ;
      RECT 6.72 5.1 7.04 5.36 ;
      RECT 77.545 5.16 79.895 5.3 ;
      RECT 79.755 4.435 79.895 5.3 ;
      RECT 59.605 5.16 61.955 5.3 ;
      RECT 61.815 4.435 61.955 5.3 ;
      RECT 41.67 5.16 44.02 5.3 ;
      RECT 43.88 4.435 44.02 5.3 ;
      RECT 23.73 5.16 26.08 5.3 ;
      RECT 25.94 4.435 26.08 5.3 ;
      RECT 5.79 5.16 8.14 5.3 ;
      RECT 8 4.435 8.14 5.3 ;
      RECT 77.545 4.435 77.685 5.3 ;
      RECT 59.605 4.435 59.745 5.3 ;
      RECT 41.67 4.435 41.81 5.3 ;
      RECT 23.73 4.435 23.87 5.3 ;
      RECT 5.79 4.435 5.93 5.3 ;
      RECT 79.68 4.435 79.97 4.665 ;
      RECT 77.47 4.435 77.76 4.665 ;
      RECT 61.74 4.435 62.03 4.665 ;
      RECT 59.53 4.435 59.82 4.665 ;
      RECT 43.805 4.435 44.095 4.665 ;
      RECT 41.595 4.435 41.885 4.665 ;
      RECT 25.865 4.435 26.155 4.665 ;
      RECT 23.655 4.435 23.945 4.665 ;
      RECT 7.925 4.435 8.215 4.665 ;
      RECT 5.715 4.435 6.005 4.665 ;
      RECT 83.24 5.185 87.69 5.35 ;
      RECT 87.525 4.435 87.69 5.35 ;
      RECT 83.16 4.97 83.33 5.235 ;
      RECT 83.1 4.99 83.38 5.235 ;
      RECT 87.525 4.435 87.695 4.725 ;
      RECT 87.49 4.465 87.74 4.7 ;
      RECT 87.505 0.7 87.675 1.605 ;
      RECT 87.475 1.345 87.705 1.58 ;
      RECT 83.065 0.82 83.325 1.05 ;
      RECT 83.065 0.85 84.4 1.02 ;
      RECT 84.23 0.7 87.675 0.87 ;
      RECT 82.555 1.36 82.875 1.62 ;
      RECT 82.28 1.42 82.875 1.56 ;
      RECT 81.95 1.7 82.29 2.04 ;
      RECT 80.175 1.7 80.495 1.96 ;
      RECT 81.95 1.715 82.44 1.945 ;
      RECT 80.175 1.76 82.44 1.9 ;
      RECT 81.535 4.42 81.855 4.68 ;
      RECT 81.535 4.48 82.13 4.62 ;
      RECT 80.855 1.36 81.175 1.62 ;
      RECT 76.115 1.375 76.405 1.605 ;
      RECT 76.115 1.42 81.175 1.56 ;
      RECT 80.945 1.08 81.085 1.62 ;
      RECT 80.945 1.08 81.425 1.22 ;
      RECT 81.285 0.695 81.425 1.22 ;
      RECT 81.21 0.695 81.5 0.925 ;
      RECT 80.855 2.38 81.175 2.64 ;
      RECT 80.19 2.395 80.48 2.625 ;
      RECT 77.98 2.395 78.27 2.625 ;
      RECT 77.98 2.44 81.175 2.58 ;
      RECT 79.155 4.42 79.475 4.68 ;
      RECT 80.87 4.435 81.16 4.665 ;
      RECT 78.49 4.435 78.78 4.665 ;
      RECT 78.49 4.48 79.475 4.62 ;
      RECT 80.945 4.14 81.085 4.665 ;
      RECT 79.245 4.14 79.385 4.68 ;
      RECT 79.245 4.14 81.085 4.28 ;
      RECT 78.15 1.035 78.44 1.265 ;
      RECT 78.225 0.74 78.365 1.265 ;
      RECT 80.515 0.68 80.835 0.94 ;
      RECT 80.415 0.695 80.835 0.925 ;
      RECT 78.225 0.74 80.835 0.88 ;
      RECT 79.495 1.02 79.815 1.28 ;
      RECT 79.495 1.08 80.09 1.22 ;
      RECT 79.495 3.4 79.815 3.66 ;
      RECT 76.79 3.415 77.08 3.645 ;
      RECT 76.79 3.46 79.815 3.6 ;
      RECT 78.82 0.98 79.15 1.31 ;
      RECT 78.815 1.015 79.15 1.275 ;
      RECT 79.165 1.035 79.28 1.265 ;
      RECT 78.815 1.03 79.165 1.26 ;
      RECT 78.815 1.08 79.295 1.22 ;
      RECT 78.7 1.08 78.71 1.22 ;
      RECT 78.71 1.075 79.28 1.215 ;
      RECT 74.23 3.875 74.6 4.245 ;
      RECT 74.23 3.655 74.4 4.245 ;
      RECT 71.335 3.625 71.565 3.855 ;
      RECT 71.305 3.655 74.4 3.825 ;
      RECT 65.3 5.185 69.75 5.35 ;
      RECT 69.585 4.435 69.75 5.35 ;
      RECT 65.22 4.97 65.39 5.235 ;
      RECT 65.16 4.99 65.44 5.235 ;
      RECT 69.585 4.435 69.755 4.725 ;
      RECT 69.55 4.465 69.8 4.7 ;
      RECT 69.565 0.7 69.735 1.605 ;
      RECT 69.535 1.345 69.765 1.58 ;
      RECT 65.125 0.82 65.385 1.05 ;
      RECT 65.125 0.85 66.46 1.02 ;
      RECT 66.29 0.7 69.735 0.87 ;
      RECT 64.615 1.36 64.935 1.62 ;
      RECT 64.34 1.42 64.935 1.56 ;
      RECT 64.01 1.7 64.35 2.04 ;
      RECT 62.235 1.7 62.555 1.96 ;
      RECT 64.01 1.715 64.5 1.945 ;
      RECT 62.235 1.76 64.5 1.9 ;
      RECT 63.595 4.42 63.915 4.68 ;
      RECT 63.595 4.48 64.19 4.62 ;
      RECT 62.915 1.36 63.235 1.62 ;
      RECT 58.175 1.375 58.465 1.605 ;
      RECT 58.175 1.42 63.235 1.56 ;
      RECT 63.005 1.08 63.145 1.62 ;
      RECT 63.005 1.08 63.485 1.22 ;
      RECT 63.345 0.695 63.485 1.22 ;
      RECT 63.27 0.695 63.56 0.925 ;
      RECT 62.915 2.38 63.235 2.64 ;
      RECT 62.25 2.395 62.54 2.625 ;
      RECT 60.04 2.395 60.33 2.625 ;
      RECT 60.04 2.44 63.235 2.58 ;
      RECT 61.215 4.42 61.535 4.68 ;
      RECT 62.93 4.435 63.22 4.665 ;
      RECT 60.55 4.435 60.84 4.665 ;
      RECT 60.55 4.48 61.535 4.62 ;
      RECT 63.005 4.14 63.145 4.665 ;
      RECT 61.305 4.14 61.445 4.68 ;
      RECT 61.305 4.14 63.145 4.28 ;
      RECT 60.21 1.035 60.5 1.265 ;
      RECT 60.285 0.74 60.425 1.265 ;
      RECT 62.575 0.68 62.895 0.94 ;
      RECT 62.475 0.695 62.895 0.925 ;
      RECT 60.285 0.74 62.895 0.88 ;
      RECT 61.555 1.02 61.875 1.28 ;
      RECT 61.555 1.08 62.15 1.22 ;
      RECT 61.555 3.4 61.875 3.66 ;
      RECT 58.85 3.415 59.14 3.645 ;
      RECT 58.85 3.46 61.875 3.6 ;
      RECT 60.88 0.98 61.21 1.31 ;
      RECT 60.875 1.015 61.21 1.275 ;
      RECT 61.225 1.035 61.34 1.265 ;
      RECT 60.875 1.03 61.225 1.26 ;
      RECT 60.875 1.08 61.355 1.22 ;
      RECT 60.76 1.08 60.77 1.22 ;
      RECT 60.77 1.075 61.34 1.215 ;
      RECT 56.29 3.875 56.66 4.245 ;
      RECT 56.29 3.655 56.5 4.245 ;
      RECT 53.4 3.625 53.63 3.855 ;
      RECT 53.37 3.655 56.5 3.825 ;
      RECT 47.365 5.185 51.815 5.35 ;
      RECT 51.65 4.435 51.815 5.35 ;
      RECT 47.285 4.97 47.455 5.235 ;
      RECT 47.225 4.99 47.505 5.235 ;
      RECT 51.65 4.435 51.82 4.725 ;
      RECT 51.615 4.465 51.865 4.7 ;
      RECT 51.63 0.7 51.8 1.605 ;
      RECT 51.6 1.345 51.83 1.58 ;
      RECT 47.19 0.82 47.45 1.05 ;
      RECT 47.19 0.85 48.525 1.02 ;
      RECT 48.355 0.7 51.8 0.87 ;
      RECT 46.68 1.36 47 1.62 ;
      RECT 46.405 1.42 47 1.56 ;
      RECT 46.075 1.7 46.415 2.04 ;
      RECT 44.3 1.7 44.62 1.96 ;
      RECT 46.075 1.715 46.565 1.945 ;
      RECT 44.3 1.76 46.565 1.9 ;
      RECT 45.66 4.42 45.98 4.68 ;
      RECT 45.66 4.48 46.255 4.62 ;
      RECT 44.98 1.36 45.3 1.62 ;
      RECT 40.24 1.375 40.53 1.605 ;
      RECT 40.24 1.42 45.3 1.56 ;
      RECT 45.07 1.08 45.21 1.62 ;
      RECT 45.07 1.08 45.55 1.22 ;
      RECT 45.41 0.695 45.55 1.22 ;
      RECT 45.335 0.695 45.625 0.925 ;
      RECT 44.98 2.38 45.3 2.64 ;
      RECT 44.315 2.395 44.605 2.625 ;
      RECT 42.105 2.395 42.395 2.625 ;
      RECT 42.105 2.44 45.3 2.58 ;
      RECT 43.28 4.42 43.6 4.68 ;
      RECT 44.995 4.435 45.285 4.665 ;
      RECT 42.615 4.435 42.905 4.665 ;
      RECT 42.615 4.48 43.6 4.62 ;
      RECT 45.07 4.14 45.21 4.665 ;
      RECT 43.37 4.14 43.51 4.68 ;
      RECT 43.37 4.14 45.21 4.28 ;
      RECT 42.275 1.035 42.565 1.265 ;
      RECT 42.35 0.74 42.49 1.265 ;
      RECT 44.64 0.68 44.96 0.94 ;
      RECT 44.54 0.695 44.96 0.925 ;
      RECT 42.35 0.74 44.96 0.88 ;
      RECT 43.62 1.02 43.94 1.28 ;
      RECT 43.62 1.08 44.215 1.22 ;
      RECT 43.62 3.4 43.94 3.66 ;
      RECT 40.915 3.415 41.205 3.645 ;
      RECT 40.915 3.46 43.94 3.6 ;
      RECT 42.945 0.98 43.275 1.31 ;
      RECT 42.94 1.015 43.275 1.275 ;
      RECT 43.29 1.035 43.405 1.265 ;
      RECT 42.94 1.03 43.29 1.26 ;
      RECT 42.94 1.08 43.42 1.22 ;
      RECT 42.825 1.08 42.835 1.22 ;
      RECT 42.835 1.075 43.405 1.215 ;
      RECT 38.355 3.875 38.725 4.245 ;
      RECT 38.35 3.655 38.52 3.93 ;
      RECT 35.46 3.625 35.69 3.855 ;
      RECT 35.43 3.655 38.52 3.825 ;
      RECT 29.425 5.185 33.875 5.35 ;
      RECT 33.71 4.435 33.875 5.35 ;
      RECT 29.345 4.97 29.515 5.235 ;
      RECT 29.285 4.99 29.565 5.235 ;
      RECT 33.71 4.435 33.88 4.725 ;
      RECT 33.675 4.465 33.925 4.7 ;
      RECT 33.69 0.7 33.86 1.605 ;
      RECT 33.66 1.345 33.89 1.58 ;
      RECT 29.25 0.82 29.51 1.05 ;
      RECT 29.25 0.85 30.585 1.02 ;
      RECT 30.415 0.7 33.86 0.87 ;
      RECT 28.74 1.36 29.06 1.62 ;
      RECT 28.465 1.42 29.06 1.56 ;
      RECT 28.135 1.7 28.475 2.04 ;
      RECT 26.36 1.7 26.68 1.96 ;
      RECT 28.135 1.715 28.625 1.945 ;
      RECT 26.36 1.76 28.625 1.9 ;
      RECT 27.72 4.42 28.04 4.68 ;
      RECT 27.72 4.48 28.315 4.62 ;
      RECT 27.04 1.36 27.36 1.62 ;
      RECT 22.3 1.375 22.59 1.605 ;
      RECT 22.3 1.42 27.36 1.56 ;
      RECT 27.13 1.08 27.27 1.62 ;
      RECT 27.13 1.08 27.61 1.22 ;
      RECT 27.47 0.695 27.61 1.22 ;
      RECT 27.395 0.695 27.685 0.925 ;
      RECT 27.04 2.38 27.36 2.64 ;
      RECT 26.375 2.395 26.665 2.625 ;
      RECT 24.165 2.395 24.455 2.625 ;
      RECT 24.165 2.44 27.36 2.58 ;
      RECT 25.34 4.42 25.66 4.68 ;
      RECT 27.055 4.435 27.345 4.665 ;
      RECT 24.675 4.435 24.965 4.665 ;
      RECT 24.675 4.48 25.66 4.62 ;
      RECT 27.13 4.14 27.27 4.665 ;
      RECT 25.43 4.14 25.57 4.68 ;
      RECT 25.43 4.14 27.27 4.28 ;
      RECT 24.335 1.035 24.625 1.265 ;
      RECT 24.41 0.74 24.55 1.265 ;
      RECT 26.7 0.68 27.02 0.94 ;
      RECT 26.6 0.695 27.02 0.925 ;
      RECT 24.41 0.74 27.02 0.88 ;
      RECT 25.68 1.02 26 1.28 ;
      RECT 25.68 1.08 26.275 1.22 ;
      RECT 25.68 3.4 26 3.66 ;
      RECT 22.975 3.415 23.265 3.645 ;
      RECT 22.975 3.46 26 3.6 ;
      RECT 25.005 0.98 25.335 1.31 ;
      RECT 25 1.015 25.335 1.275 ;
      RECT 25.35 1.035 25.465 1.265 ;
      RECT 25 1.03 25.35 1.26 ;
      RECT 25 1.08 25.48 1.22 ;
      RECT 24.885 1.08 24.895 1.22 ;
      RECT 24.895 1.075 25.465 1.215 ;
      RECT 20.415 3.875 20.785 4.245 ;
      RECT 20.415 3.655 20.685 4.245 ;
      RECT 17.505 3.61 17.765 3.86 ;
      RECT 17.49 3.655 20.685 3.825 ;
      RECT 11.485 5.185 15.935 5.35 ;
      RECT 15.77 4.435 15.935 5.35 ;
      RECT 11.405 4.97 11.575 5.235 ;
      RECT 11.345 4.99 11.625 5.235 ;
      RECT 15.77 4.435 15.94 4.725 ;
      RECT 15.735 4.465 15.985 4.7 ;
      RECT 15.75 0.7 15.92 1.605 ;
      RECT 15.72 1.345 15.95 1.58 ;
      RECT 11.31 0.82 11.57 1.05 ;
      RECT 11.31 0.85 12.645 1.02 ;
      RECT 12.475 0.7 15.92 0.87 ;
      RECT 10.8 1.36 11.12 1.62 ;
      RECT 10.525 1.42 11.12 1.56 ;
      RECT 10.195 1.7 10.535 2.04 ;
      RECT 8.42 1.7 8.74 1.96 ;
      RECT 10.195 1.715 10.685 1.945 ;
      RECT 8.42 1.76 10.685 1.9 ;
      RECT 9.78 4.42 10.1 4.68 ;
      RECT 9.78 4.48 10.375 4.62 ;
      RECT 9.1 1.36 9.42 1.62 ;
      RECT 4.36 1.375 4.65 1.605 ;
      RECT 4.36 1.42 9.42 1.56 ;
      RECT 9.19 1.08 9.33 1.62 ;
      RECT 9.19 1.08 9.67 1.22 ;
      RECT 9.53 0.695 9.67 1.22 ;
      RECT 9.455 0.695 9.745 0.925 ;
      RECT 9.1 2.38 9.42 2.64 ;
      RECT 8.435 2.395 8.725 2.625 ;
      RECT 6.225 2.395 6.515 2.625 ;
      RECT 6.225 2.44 9.42 2.58 ;
      RECT 7.4 4.42 7.72 4.68 ;
      RECT 9.115 4.435 9.405 4.665 ;
      RECT 6.735 4.435 7.025 4.665 ;
      RECT 6.735 4.48 7.72 4.62 ;
      RECT 9.19 4.14 9.33 4.665 ;
      RECT 7.49 4.14 7.63 4.68 ;
      RECT 7.49 4.14 9.33 4.28 ;
      RECT 6.395 1.035 6.685 1.265 ;
      RECT 6.47 0.74 6.61 1.265 ;
      RECT 8.76 0.68 9.08 0.94 ;
      RECT 8.66 0.695 9.08 0.925 ;
      RECT 6.47 0.74 9.08 0.88 ;
      RECT 7.74 1.02 8.06 1.28 ;
      RECT 7.74 1.08 8.335 1.22 ;
      RECT 7.74 3.4 8.06 3.66 ;
      RECT 5.035 3.415 5.325 3.645 ;
      RECT 5.035 3.46 8.06 3.6 ;
      RECT 7.065 0.98 7.395 1.31 ;
      RECT 7.06 1.015 7.395 1.275 ;
      RECT 7.41 1.035 7.525 1.265 ;
      RECT 7.06 1.03 7.41 1.26 ;
      RECT 7.06 1.08 7.54 1.22 ;
      RECT 6.945 1.08 6.955 1.22 ;
      RECT 6.955 1.075 7.525 1.215 ;
      RECT -0.015 4.855 0.415 5.275 ;
      RECT -1.855 4.925 0.415 5.115 ;
      RECT -1.855 4.645 -1.65 5.115 ;
      RECT -1.885 4.645 -1.65 4.875 ;
      RECT -1.855 4.615 -1.685 5.115 ;
      RECT -3.95 0.06 89.885 0.54 ;
      RECT 89.24 4.86 89.67 5.28 ;
      RECT 85.41 1.7 85.75 2.04 ;
      RECT 85.365 3.97 85.705 4.31 ;
      RECT 84.96 1.11 85.3 1.45 ;
      RECT 84.945 4.575 85.285 4.915 ;
      RECT 83.81 4.415 84.15 4.755 ;
      RECT 83.825 1.295 84.145 1.615 ;
      RECT 82.23 3.4 82.875 3.66 ;
      RECT 80.175 4.42 80.495 4.68 ;
      RECT 75.76 4.38 76.13 4.75 ;
      RECT 72.525 4.02 72.895 4.39 ;
      RECT 67.47 1.7 67.81 2.04 ;
      RECT 67.425 3.97 67.765 4.31 ;
      RECT 67.02 1.11 67.36 1.45 ;
      RECT 67.005 4.575 67.345 4.915 ;
      RECT 65.87 4.415 66.21 4.755 ;
      RECT 65.885 1.295 66.205 1.615 ;
      RECT 64.29 3.4 64.935 3.66 ;
      RECT 62.235 4.42 62.555 4.68 ;
      RECT 57.82 4.38 58.19 4.75 ;
      RECT 54.585 4.02 54.955 4.39 ;
      RECT 49.535 1.7 49.875 2.04 ;
      RECT 49.49 3.97 49.83 4.31 ;
      RECT 49.085 1.11 49.425 1.45 ;
      RECT 49.07 4.575 49.41 4.915 ;
      RECT 47.935 4.415 48.275 4.755 ;
      RECT 47.95 1.295 48.27 1.615 ;
      RECT 46.355 3.4 47 3.66 ;
      RECT 44.3 4.42 44.62 4.68 ;
      RECT 39.885 4.38 40.255 4.75 ;
      RECT 36.65 4.02 37.02 4.39 ;
      RECT 31.595 1.7 31.935 2.04 ;
      RECT 31.55 3.97 31.89 4.31 ;
      RECT 31.145 1.11 31.485 1.45 ;
      RECT 31.13 4.575 31.47 4.915 ;
      RECT 29.995 4.415 30.335 4.755 ;
      RECT 30.01 1.295 30.33 1.615 ;
      RECT 28.415 3.4 29.06 3.66 ;
      RECT 26.36 4.42 26.68 4.68 ;
      RECT 21.945 4.38 22.315 4.75 ;
      RECT 18.71 4.02 19.08 4.39 ;
      RECT 13.655 1.7 13.995 2.04 ;
      RECT 13.61 3.97 13.95 4.31 ;
      RECT 13.205 1.11 13.545 1.45 ;
      RECT 13.19 4.575 13.53 4.915 ;
      RECT 12.055 4.415 12.395 4.755 ;
      RECT 12.07 1.295 12.39 1.615 ;
      RECT 10.475 3.4 11.12 3.66 ;
      RECT 8.42 4.42 8.74 4.68 ;
      RECT 4.005 4.38 4.375 4.75 ;
      RECT 2.475 3.875 2.845 4.245 ;
      RECT 0.77 4.02 1.14 4.39 ;
      RECT -3.885 3.55 -3.505 3.93 ;
    LAYER mcon ;
      RECT 89.57 0.215 89.74 0.385 ;
      RECT 89.57 2.935 89.74 3.105 ;
      RECT 89.57 5.655 89.74 5.825 ;
      RECT 89.305 4.915 89.475 5.085 ;
      RECT 89.11 0.215 89.28 0.385 ;
      RECT 89.11 2.935 89.28 3.105 ;
      RECT 89.11 5.655 89.28 5.825 ;
      RECT 88.65 0.215 88.82 0.385 ;
      RECT 88.65 2.935 88.82 3.105 ;
      RECT 88.65 5.655 88.82 5.825 ;
      RECT 88.19 0.215 88.36 0.385 ;
      RECT 88.19 2.935 88.36 3.105 ;
      RECT 88.19 5.655 88.36 5.825 ;
      RECT 87.73 0.215 87.9 0.385 ;
      RECT 87.73 2.935 87.9 3.105 ;
      RECT 87.73 5.655 87.9 5.825 ;
      RECT 87.525 4.495 87.695 4.665 ;
      RECT 87.505 1.375 87.675 1.545 ;
      RECT 87.27 0.215 87.44 0.385 ;
      RECT 87.27 2.935 87.44 3.105 ;
      RECT 87.27 5.655 87.44 5.825 ;
      RECT 86.81 0.215 86.98 0.385 ;
      RECT 86.81 2.935 86.98 3.105 ;
      RECT 86.81 5.655 86.98 5.825 ;
      RECT 86.35 0.215 86.52 0.385 ;
      RECT 86.35 2.935 86.52 3.105 ;
      RECT 86.35 5.655 86.52 5.825 ;
      RECT 85.89 0.215 86.06 0.385 ;
      RECT 85.89 2.935 86.06 3.105 ;
      RECT 85.89 5.655 86.06 5.825 ;
      RECT 85.44 1.76 85.61 1.93 ;
      RECT 85.44 4.11 85.61 4.28 ;
      RECT 85.43 0.215 85.6 0.385 ;
      RECT 85.43 2.935 85.6 3.105 ;
      RECT 85.43 5.655 85.6 5.825 ;
      RECT 85.08 1.195 85.25 1.365 ;
      RECT 85.08 4.675 85.25 4.845 ;
      RECT 84.97 0.215 85.14 0.385 ;
      RECT 84.97 2.935 85.14 3.105 ;
      RECT 84.97 5.655 85.14 5.825 ;
      RECT 84.51 0.215 84.68 0.385 ;
      RECT 84.51 2.935 84.68 3.105 ;
      RECT 84.51 5.655 84.68 5.825 ;
      RECT 84.05 0.215 84.22 0.385 ;
      RECT 84.05 2.935 84.22 3.105 ;
      RECT 84.05 5.655 84.22 5.825 ;
      RECT 83.895 1.375 84.065 1.545 ;
      RECT 83.895 4.495 84.065 4.665 ;
      RECT 83.59 0.215 83.76 0.385 ;
      RECT 83.59 2.935 83.76 3.105 ;
      RECT 83.59 5.655 83.76 5.825 ;
      RECT 83.16 5.03 83.33 5.2 ;
      RECT 83.13 0.215 83.3 0.385 ;
      RECT 83.13 2.935 83.3 3.105 ;
      RECT 83.13 5.655 83.3 5.825 ;
      RECT 83.125 0.85 83.295 1.02 ;
      RECT 82.67 0.215 82.84 0.385 ;
      RECT 82.67 2.935 82.84 3.105 ;
      RECT 82.67 5.655 82.84 5.825 ;
      RECT 82.63 1.405 82.8 1.575 ;
      RECT 82.29 3.445 82.46 3.615 ;
      RECT 82.21 0.215 82.38 0.385 ;
      RECT 82.21 1.745 82.38 1.915 ;
      RECT 82.21 2.935 82.38 3.105 ;
      RECT 82.21 5.655 82.38 5.825 ;
      RECT 81.75 0.215 81.92 0.385 ;
      RECT 81.75 2.935 81.92 3.105 ;
      RECT 81.75 5.655 81.92 5.825 ;
      RECT 81.61 4.465 81.78 4.635 ;
      RECT 81.29 0.215 81.46 0.385 ;
      RECT 81.29 2.935 81.46 3.105 ;
      RECT 81.29 5.655 81.46 5.825 ;
      RECT 81.27 0.725 81.44 0.895 ;
      RECT 80.93 4.465 81.1 4.635 ;
      RECT 80.83 0.215 81 0.385 ;
      RECT 80.83 2.935 81 3.105 ;
      RECT 80.83 5.655 81 5.825 ;
      RECT 80.475 0.725 80.645 0.895 ;
      RECT 80.37 0.215 80.54 0.385 ;
      RECT 80.37 2.935 80.54 3.105 ;
      RECT 80.37 5.655 80.54 5.825 ;
      RECT 80.25 2.425 80.42 2.595 ;
      RECT 80.25 4.465 80.42 4.635 ;
      RECT 79.91 0.215 80.08 0.385 ;
      RECT 79.91 2.935 80.08 3.105 ;
      RECT 79.91 5.655 80.08 5.825 ;
      RECT 79.74 4.465 79.91 4.635 ;
      RECT 79.57 1.065 79.74 1.235 ;
      RECT 79.45 0.215 79.62 0.385 ;
      RECT 79.45 2.935 79.62 3.105 ;
      RECT 79.45 5.655 79.62 5.825 ;
      RECT 78.99 0.215 79.16 0.385 ;
      RECT 78.99 2.935 79.16 3.105 ;
      RECT 78.99 5.655 79.16 5.825 ;
      RECT 78.55 4.465 78.72 4.635 ;
      RECT 78.53 0.215 78.7 0.385 ;
      RECT 78.53 2.935 78.7 3.105 ;
      RECT 78.53 5.655 78.7 5.825 ;
      RECT 78.21 1.065 78.38 1.235 ;
      RECT 78.07 0.215 78.24 0.385 ;
      RECT 78.07 2.935 78.24 3.105 ;
      RECT 78.07 5.655 78.24 5.825 ;
      RECT 78.04 2.425 78.21 2.595 ;
      RECT 77.61 0.215 77.78 0.385 ;
      RECT 77.61 2.935 77.78 3.105 ;
      RECT 77.61 5.655 77.78 5.825 ;
      RECT 77.53 4.465 77.7 4.635 ;
      RECT 77.15 0.215 77.32 0.385 ;
      RECT 77.15 2.935 77.32 3.105 ;
      RECT 77.15 5.655 77.32 5.825 ;
      RECT 76.85 3.445 77.02 3.615 ;
      RECT 76.69 0.215 76.86 0.385 ;
      RECT 76.69 2.935 76.86 3.105 ;
      RECT 76.69 5.655 76.86 5.825 ;
      RECT 76.23 0.215 76.4 0.385 ;
      RECT 76.23 2.935 76.4 3.105 ;
      RECT 76.23 5.655 76.4 5.825 ;
      RECT 76.175 1.405 76.345 1.575 ;
      RECT 75.83 4.485 76 4.655 ;
      RECT 75.77 2.935 75.94 3.105 ;
      RECT 75.77 5.655 75.94 5.825 ;
      RECT 75.31 2.935 75.48 3.105 ;
      RECT 75.31 5.655 75.48 5.825 ;
      RECT 74.85 2.935 75.02 3.105 ;
      RECT 74.85 5.655 75.02 5.825 ;
      RECT 74.39 2.935 74.56 3.105 ;
      RECT 74.39 5.655 74.56 5.825 ;
      RECT 74.3 3.98 74.47 4.15 ;
      RECT 73.93 2.935 74.1 3.105 ;
      RECT 73.93 5.655 74.1 5.825 ;
      RECT 73.47 2.935 73.64 3.105 ;
      RECT 73.47 5.655 73.64 5.825 ;
      RECT 73.01 2.935 73.18 3.105 ;
      RECT 73.01 5.655 73.18 5.825 ;
      RECT 72.62 4.11 72.79 4.28 ;
      RECT 72.55 2.935 72.72 3.105 ;
      RECT 72.55 5.655 72.72 5.825 ;
      RECT 72.09 2.935 72.26 3.105 ;
      RECT 72.09 5.655 72.26 5.825 ;
      RECT 71.63 0.215 71.8 0.385 ;
      RECT 71.63 2.935 71.8 3.105 ;
      RECT 71.63 5.655 71.8 5.825 ;
      RECT 71.365 3.655 71.535 3.825 ;
      RECT 71.17 0.215 71.34 0.385 ;
      RECT 71.17 2.935 71.34 3.105 ;
      RECT 71.17 5.655 71.34 5.825 ;
      RECT 70.71 0.215 70.88 0.385 ;
      RECT 70.71 2.935 70.88 3.105 ;
      RECT 70.71 5.655 70.88 5.825 ;
      RECT 70.25 0.215 70.42 0.385 ;
      RECT 70.25 2.935 70.42 3.105 ;
      RECT 70.25 5.655 70.42 5.825 ;
      RECT 69.79 0.215 69.96 0.385 ;
      RECT 69.79 2.935 69.96 3.105 ;
      RECT 69.79 5.655 69.96 5.825 ;
      RECT 69.585 4.495 69.755 4.665 ;
      RECT 69.565 1.375 69.735 1.545 ;
      RECT 69.33 0.215 69.5 0.385 ;
      RECT 69.33 2.935 69.5 3.105 ;
      RECT 69.33 5.655 69.5 5.825 ;
      RECT 68.87 0.215 69.04 0.385 ;
      RECT 68.87 2.935 69.04 3.105 ;
      RECT 68.87 5.655 69.04 5.825 ;
      RECT 68.41 0.215 68.58 0.385 ;
      RECT 68.41 2.935 68.58 3.105 ;
      RECT 68.41 5.655 68.58 5.825 ;
      RECT 67.95 0.215 68.12 0.385 ;
      RECT 67.95 2.935 68.12 3.105 ;
      RECT 67.95 5.655 68.12 5.825 ;
      RECT 67.5 1.76 67.67 1.93 ;
      RECT 67.5 4.11 67.67 4.28 ;
      RECT 67.49 0.215 67.66 0.385 ;
      RECT 67.49 2.935 67.66 3.105 ;
      RECT 67.49 5.655 67.66 5.825 ;
      RECT 67.14 1.195 67.31 1.365 ;
      RECT 67.14 4.675 67.31 4.845 ;
      RECT 67.03 0.215 67.2 0.385 ;
      RECT 67.03 2.935 67.2 3.105 ;
      RECT 67.03 5.655 67.2 5.825 ;
      RECT 66.57 0.215 66.74 0.385 ;
      RECT 66.57 2.935 66.74 3.105 ;
      RECT 66.57 5.655 66.74 5.825 ;
      RECT 66.11 0.215 66.28 0.385 ;
      RECT 66.11 2.935 66.28 3.105 ;
      RECT 66.11 5.655 66.28 5.825 ;
      RECT 65.955 1.375 66.125 1.545 ;
      RECT 65.955 4.495 66.125 4.665 ;
      RECT 65.65 0.215 65.82 0.385 ;
      RECT 65.65 2.935 65.82 3.105 ;
      RECT 65.65 5.655 65.82 5.825 ;
      RECT 65.22 5.03 65.39 5.2 ;
      RECT 65.19 0.215 65.36 0.385 ;
      RECT 65.19 2.935 65.36 3.105 ;
      RECT 65.19 5.655 65.36 5.825 ;
      RECT 65.185 0.85 65.355 1.02 ;
      RECT 64.73 0.215 64.9 0.385 ;
      RECT 64.73 2.935 64.9 3.105 ;
      RECT 64.73 5.655 64.9 5.825 ;
      RECT 64.69 1.405 64.86 1.575 ;
      RECT 64.35 3.445 64.52 3.615 ;
      RECT 64.27 0.215 64.44 0.385 ;
      RECT 64.27 1.745 64.44 1.915 ;
      RECT 64.27 2.935 64.44 3.105 ;
      RECT 64.27 5.655 64.44 5.825 ;
      RECT 63.81 0.215 63.98 0.385 ;
      RECT 63.81 2.935 63.98 3.105 ;
      RECT 63.81 5.655 63.98 5.825 ;
      RECT 63.67 4.465 63.84 4.635 ;
      RECT 63.35 0.215 63.52 0.385 ;
      RECT 63.35 2.935 63.52 3.105 ;
      RECT 63.35 5.655 63.52 5.825 ;
      RECT 63.33 0.725 63.5 0.895 ;
      RECT 62.99 4.465 63.16 4.635 ;
      RECT 62.89 0.215 63.06 0.385 ;
      RECT 62.89 2.935 63.06 3.105 ;
      RECT 62.89 5.655 63.06 5.825 ;
      RECT 62.535 0.725 62.705 0.895 ;
      RECT 62.43 0.215 62.6 0.385 ;
      RECT 62.43 2.935 62.6 3.105 ;
      RECT 62.43 5.655 62.6 5.825 ;
      RECT 62.31 2.425 62.48 2.595 ;
      RECT 62.31 4.465 62.48 4.635 ;
      RECT 61.97 0.215 62.14 0.385 ;
      RECT 61.97 2.935 62.14 3.105 ;
      RECT 61.97 5.655 62.14 5.825 ;
      RECT 61.8 4.465 61.97 4.635 ;
      RECT 61.63 1.065 61.8 1.235 ;
      RECT 61.51 0.215 61.68 0.385 ;
      RECT 61.51 2.935 61.68 3.105 ;
      RECT 61.51 5.655 61.68 5.825 ;
      RECT 61.05 0.215 61.22 0.385 ;
      RECT 61.05 2.935 61.22 3.105 ;
      RECT 61.05 5.655 61.22 5.825 ;
      RECT 60.61 4.465 60.78 4.635 ;
      RECT 60.59 0.215 60.76 0.385 ;
      RECT 60.59 2.935 60.76 3.105 ;
      RECT 60.59 5.655 60.76 5.825 ;
      RECT 60.27 1.065 60.44 1.235 ;
      RECT 60.13 0.215 60.3 0.385 ;
      RECT 60.13 2.935 60.3 3.105 ;
      RECT 60.13 5.655 60.3 5.825 ;
      RECT 60.1 2.425 60.27 2.595 ;
      RECT 59.67 0.215 59.84 0.385 ;
      RECT 59.67 2.935 59.84 3.105 ;
      RECT 59.67 5.655 59.84 5.825 ;
      RECT 59.59 4.465 59.76 4.635 ;
      RECT 59.21 0.215 59.38 0.385 ;
      RECT 59.21 2.935 59.38 3.105 ;
      RECT 59.21 5.655 59.38 5.825 ;
      RECT 58.91 3.445 59.08 3.615 ;
      RECT 58.75 0.215 58.92 0.385 ;
      RECT 58.75 2.935 58.92 3.105 ;
      RECT 58.75 5.655 58.92 5.825 ;
      RECT 58.29 0.215 58.46 0.385 ;
      RECT 58.29 2.935 58.46 3.105 ;
      RECT 58.29 5.655 58.46 5.825 ;
      RECT 58.235 1.405 58.405 1.575 ;
      RECT 57.89 4.485 58.06 4.655 ;
      RECT 57.83 2.935 58 3.105 ;
      RECT 57.83 5.655 58 5.825 ;
      RECT 57.37 2.935 57.54 3.105 ;
      RECT 57.37 5.655 57.54 5.825 ;
      RECT 56.91 2.935 57.08 3.105 ;
      RECT 56.91 5.655 57.08 5.825 ;
      RECT 56.45 2.935 56.62 3.105 ;
      RECT 56.45 5.655 56.62 5.825 ;
      RECT 56.36 3.98 56.53 4.15 ;
      RECT 55.99 2.935 56.16 3.105 ;
      RECT 55.99 5.655 56.16 5.825 ;
      RECT 55.53 2.935 55.7 3.105 ;
      RECT 55.53 5.655 55.7 5.825 ;
      RECT 55.07 2.935 55.24 3.105 ;
      RECT 55.07 5.655 55.24 5.825 ;
      RECT 54.68 4.11 54.85 4.28 ;
      RECT 54.61 2.935 54.78 3.105 ;
      RECT 54.61 5.655 54.78 5.825 ;
      RECT 54.15 2.935 54.32 3.105 ;
      RECT 54.15 5.655 54.32 5.825 ;
      RECT 53.695 0.215 53.865 0.385 ;
      RECT 53.695 2.935 53.865 3.105 ;
      RECT 53.695 5.655 53.865 5.825 ;
      RECT 53.43 3.655 53.6 3.825 ;
      RECT 53.235 0.215 53.405 0.385 ;
      RECT 53.235 2.935 53.405 3.105 ;
      RECT 53.235 5.655 53.405 5.825 ;
      RECT 52.775 0.215 52.945 0.385 ;
      RECT 52.775 2.935 52.945 3.105 ;
      RECT 52.775 5.655 52.945 5.825 ;
      RECT 52.315 0.215 52.485 0.385 ;
      RECT 52.315 2.935 52.485 3.105 ;
      RECT 52.315 5.655 52.485 5.825 ;
      RECT 51.855 0.215 52.025 0.385 ;
      RECT 51.855 2.935 52.025 3.105 ;
      RECT 51.855 5.655 52.025 5.825 ;
      RECT 51.65 4.495 51.82 4.665 ;
      RECT 51.63 1.375 51.8 1.545 ;
      RECT 51.395 0.215 51.565 0.385 ;
      RECT 51.395 2.935 51.565 3.105 ;
      RECT 51.395 5.655 51.565 5.825 ;
      RECT 50.935 0.215 51.105 0.385 ;
      RECT 50.935 2.935 51.105 3.105 ;
      RECT 50.935 5.655 51.105 5.825 ;
      RECT 50.475 0.215 50.645 0.385 ;
      RECT 50.475 2.935 50.645 3.105 ;
      RECT 50.475 5.655 50.645 5.825 ;
      RECT 50.015 0.215 50.185 0.385 ;
      RECT 50.015 2.935 50.185 3.105 ;
      RECT 50.015 5.655 50.185 5.825 ;
      RECT 49.565 1.76 49.735 1.93 ;
      RECT 49.565 4.11 49.735 4.28 ;
      RECT 49.555 0.215 49.725 0.385 ;
      RECT 49.555 2.935 49.725 3.105 ;
      RECT 49.555 5.655 49.725 5.825 ;
      RECT 49.205 1.195 49.375 1.365 ;
      RECT 49.205 4.675 49.375 4.845 ;
      RECT 49.095 0.215 49.265 0.385 ;
      RECT 49.095 2.935 49.265 3.105 ;
      RECT 49.095 5.655 49.265 5.825 ;
      RECT 48.635 0.215 48.805 0.385 ;
      RECT 48.635 2.935 48.805 3.105 ;
      RECT 48.635 5.655 48.805 5.825 ;
      RECT 48.175 0.215 48.345 0.385 ;
      RECT 48.175 2.935 48.345 3.105 ;
      RECT 48.175 5.655 48.345 5.825 ;
      RECT 48.02 1.375 48.19 1.545 ;
      RECT 48.02 4.495 48.19 4.665 ;
      RECT 47.715 0.215 47.885 0.385 ;
      RECT 47.715 2.935 47.885 3.105 ;
      RECT 47.715 5.655 47.885 5.825 ;
      RECT 47.285 5.03 47.455 5.2 ;
      RECT 47.255 0.215 47.425 0.385 ;
      RECT 47.255 2.935 47.425 3.105 ;
      RECT 47.255 5.655 47.425 5.825 ;
      RECT 47.25 0.85 47.42 1.02 ;
      RECT 46.795 0.215 46.965 0.385 ;
      RECT 46.795 2.935 46.965 3.105 ;
      RECT 46.795 5.655 46.965 5.825 ;
      RECT 46.755 1.405 46.925 1.575 ;
      RECT 46.415 3.445 46.585 3.615 ;
      RECT 46.335 0.215 46.505 0.385 ;
      RECT 46.335 1.745 46.505 1.915 ;
      RECT 46.335 2.935 46.505 3.105 ;
      RECT 46.335 5.655 46.505 5.825 ;
      RECT 45.875 0.215 46.045 0.385 ;
      RECT 45.875 2.935 46.045 3.105 ;
      RECT 45.875 5.655 46.045 5.825 ;
      RECT 45.735 4.465 45.905 4.635 ;
      RECT 45.415 0.215 45.585 0.385 ;
      RECT 45.415 2.935 45.585 3.105 ;
      RECT 45.415 5.655 45.585 5.825 ;
      RECT 45.395 0.725 45.565 0.895 ;
      RECT 45.055 4.465 45.225 4.635 ;
      RECT 44.955 0.215 45.125 0.385 ;
      RECT 44.955 2.935 45.125 3.105 ;
      RECT 44.955 5.655 45.125 5.825 ;
      RECT 44.6 0.725 44.77 0.895 ;
      RECT 44.495 0.215 44.665 0.385 ;
      RECT 44.495 2.935 44.665 3.105 ;
      RECT 44.495 5.655 44.665 5.825 ;
      RECT 44.375 2.425 44.545 2.595 ;
      RECT 44.375 4.465 44.545 4.635 ;
      RECT 44.035 0.215 44.205 0.385 ;
      RECT 44.035 2.935 44.205 3.105 ;
      RECT 44.035 5.655 44.205 5.825 ;
      RECT 43.865 4.465 44.035 4.635 ;
      RECT 43.695 1.065 43.865 1.235 ;
      RECT 43.575 0.215 43.745 0.385 ;
      RECT 43.575 2.935 43.745 3.105 ;
      RECT 43.575 5.655 43.745 5.825 ;
      RECT 43.115 0.215 43.285 0.385 ;
      RECT 43.115 2.935 43.285 3.105 ;
      RECT 43.115 5.655 43.285 5.825 ;
      RECT 42.675 4.465 42.845 4.635 ;
      RECT 42.655 0.215 42.825 0.385 ;
      RECT 42.655 2.935 42.825 3.105 ;
      RECT 42.655 5.655 42.825 5.825 ;
      RECT 42.335 1.065 42.505 1.235 ;
      RECT 42.195 0.215 42.365 0.385 ;
      RECT 42.195 2.935 42.365 3.105 ;
      RECT 42.195 5.655 42.365 5.825 ;
      RECT 42.165 2.425 42.335 2.595 ;
      RECT 41.735 0.215 41.905 0.385 ;
      RECT 41.735 2.935 41.905 3.105 ;
      RECT 41.735 5.655 41.905 5.825 ;
      RECT 41.655 4.465 41.825 4.635 ;
      RECT 41.275 0.215 41.445 0.385 ;
      RECT 41.275 2.935 41.445 3.105 ;
      RECT 41.275 5.655 41.445 5.825 ;
      RECT 40.975 3.445 41.145 3.615 ;
      RECT 40.815 0.215 40.985 0.385 ;
      RECT 40.815 2.935 40.985 3.105 ;
      RECT 40.815 5.655 40.985 5.825 ;
      RECT 40.355 0.215 40.525 0.385 ;
      RECT 40.355 2.935 40.525 3.105 ;
      RECT 40.355 5.655 40.525 5.825 ;
      RECT 40.3 1.405 40.47 1.575 ;
      RECT 39.955 4.485 40.125 4.655 ;
      RECT 39.895 2.935 40.065 3.105 ;
      RECT 39.895 5.655 40.065 5.825 ;
      RECT 39.435 2.935 39.605 3.105 ;
      RECT 39.435 5.655 39.605 5.825 ;
      RECT 38.975 2.935 39.145 3.105 ;
      RECT 38.975 5.655 39.145 5.825 ;
      RECT 38.515 2.935 38.685 3.105 ;
      RECT 38.515 5.655 38.685 5.825 ;
      RECT 38.425 3.98 38.595 4.15 ;
      RECT 38.055 2.935 38.225 3.105 ;
      RECT 38.055 5.655 38.225 5.825 ;
      RECT 37.595 2.935 37.765 3.105 ;
      RECT 37.595 5.655 37.765 5.825 ;
      RECT 37.135 2.935 37.305 3.105 ;
      RECT 37.135 5.655 37.305 5.825 ;
      RECT 36.745 4.11 36.915 4.28 ;
      RECT 36.675 2.935 36.845 3.105 ;
      RECT 36.675 5.655 36.845 5.825 ;
      RECT 36.215 2.935 36.385 3.105 ;
      RECT 36.215 5.655 36.385 5.825 ;
      RECT 35.755 0.215 35.925 0.385 ;
      RECT 35.755 2.935 35.925 3.105 ;
      RECT 35.755 5.655 35.925 5.825 ;
      RECT 35.49 3.655 35.66 3.825 ;
      RECT 35.295 0.215 35.465 0.385 ;
      RECT 35.295 2.935 35.465 3.105 ;
      RECT 35.295 5.655 35.465 5.825 ;
      RECT 34.835 0.215 35.005 0.385 ;
      RECT 34.835 2.935 35.005 3.105 ;
      RECT 34.835 5.655 35.005 5.825 ;
      RECT 34.375 0.215 34.545 0.385 ;
      RECT 34.375 2.935 34.545 3.105 ;
      RECT 34.375 5.655 34.545 5.825 ;
      RECT 33.915 0.215 34.085 0.385 ;
      RECT 33.915 2.935 34.085 3.105 ;
      RECT 33.915 5.655 34.085 5.825 ;
      RECT 33.71 4.495 33.88 4.665 ;
      RECT 33.69 1.375 33.86 1.545 ;
      RECT 33.455 0.215 33.625 0.385 ;
      RECT 33.455 2.935 33.625 3.105 ;
      RECT 33.455 5.655 33.625 5.825 ;
      RECT 32.995 0.215 33.165 0.385 ;
      RECT 32.995 2.935 33.165 3.105 ;
      RECT 32.995 5.655 33.165 5.825 ;
      RECT 32.535 0.215 32.705 0.385 ;
      RECT 32.535 2.935 32.705 3.105 ;
      RECT 32.535 5.655 32.705 5.825 ;
      RECT 32.075 0.215 32.245 0.385 ;
      RECT 32.075 2.935 32.245 3.105 ;
      RECT 32.075 5.655 32.245 5.825 ;
      RECT 31.625 1.76 31.795 1.93 ;
      RECT 31.625 4.11 31.795 4.28 ;
      RECT 31.615 0.215 31.785 0.385 ;
      RECT 31.615 2.935 31.785 3.105 ;
      RECT 31.615 5.655 31.785 5.825 ;
      RECT 31.265 1.195 31.435 1.365 ;
      RECT 31.265 4.675 31.435 4.845 ;
      RECT 31.155 0.215 31.325 0.385 ;
      RECT 31.155 2.935 31.325 3.105 ;
      RECT 31.155 5.655 31.325 5.825 ;
      RECT 30.695 0.215 30.865 0.385 ;
      RECT 30.695 2.935 30.865 3.105 ;
      RECT 30.695 5.655 30.865 5.825 ;
      RECT 30.235 0.215 30.405 0.385 ;
      RECT 30.235 2.935 30.405 3.105 ;
      RECT 30.235 5.655 30.405 5.825 ;
      RECT 30.08 1.375 30.25 1.545 ;
      RECT 30.08 4.495 30.25 4.665 ;
      RECT 29.775 0.215 29.945 0.385 ;
      RECT 29.775 2.935 29.945 3.105 ;
      RECT 29.775 5.655 29.945 5.825 ;
      RECT 29.345 5.03 29.515 5.2 ;
      RECT 29.315 0.215 29.485 0.385 ;
      RECT 29.315 2.935 29.485 3.105 ;
      RECT 29.315 5.655 29.485 5.825 ;
      RECT 29.31 0.85 29.48 1.02 ;
      RECT 28.855 0.215 29.025 0.385 ;
      RECT 28.855 2.935 29.025 3.105 ;
      RECT 28.855 5.655 29.025 5.825 ;
      RECT 28.815 1.405 28.985 1.575 ;
      RECT 28.475 3.445 28.645 3.615 ;
      RECT 28.395 0.215 28.565 0.385 ;
      RECT 28.395 1.745 28.565 1.915 ;
      RECT 28.395 2.935 28.565 3.105 ;
      RECT 28.395 5.655 28.565 5.825 ;
      RECT 27.935 0.215 28.105 0.385 ;
      RECT 27.935 2.935 28.105 3.105 ;
      RECT 27.935 5.655 28.105 5.825 ;
      RECT 27.795 4.465 27.965 4.635 ;
      RECT 27.475 0.215 27.645 0.385 ;
      RECT 27.475 2.935 27.645 3.105 ;
      RECT 27.475 5.655 27.645 5.825 ;
      RECT 27.455 0.725 27.625 0.895 ;
      RECT 27.115 4.465 27.285 4.635 ;
      RECT 27.015 0.215 27.185 0.385 ;
      RECT 27.015 2.935 27.185 3.105 ;
      RECT 27.015 5.655 27.185 5.825 ;
      RECT 26.66 0.725 26.83 0.895 ;
      RECT 26.555 0.215 26.725 0.385 ;
      RECT 26.555 2.935 26.725 3.105 ;
      RECT 26.555 5.655 26.725 5.825 ;
      RECT 26.435 2.425 26.605 2.595 ;
      RECT 26.435 4.465 26.605 4.635 ;
      RECT 26.095 0.215 26.265 0.385 ;
      RECT 26.095 2.935 26.265 3.105 ;
      RECT 26.095 5.655 26.265 5.825 ;
      RECT 25.925 4.465 26.095 4.635 ;
      RECT 25.755 1.065 25.925 1.235 ;
      RECT 25.635 0.215 25.805 0.385 ;
      RECT 25.635 2.935 25.805 3.105 ;
      RECT 25.635 5.655 25.805 5.825 ;
      RECT 25.175 0.215 25.345 0.385 ;
      RECT 25.175 2.935 25.345 3.105 ;
      RECT 25.175 5.655 25.345 5.825 ;
      RECT 24.735 4.465 24.905 4.635 ;
      RECT 24.715 0.215 24.885 0.385 ;
      RECT 24.715 2.935 24.885 3.105 ;
      RECT 24.715 5.655 24.885 5.825 ;
      RECT 24.395 1.065 24.565 1.235 ;
      RECT 24.255 0.215 24.425 0.385 ;
      RECT 24.255 2.935 24.425 3.105 ;
      RECT 24.255 5.655 24.425 5.825 ;
      RECT 24.225 2.425 24.395 2.595 ;
      RECT 23.795 0.215 23.965 0.385 ;
      RECT 23.795 2.935 23.965 3.105 ;
      RECT 23.795 5.655 23.965 5.825 ;
      RECT 23.715 4.465 23.885 4.635 ;
      RECT 23.335 0.215 23.505 0.385 ;
      RECT 23.335 2.935 23.505 3.105 ;
      RECT 23.335 5.655 23.505 5.825 ;
      RECT 23.035 3.445 23.205 3.615 ;
      RECT 22.875 0.215 23.045 0.385 ;
      RECT 22.875 2.935 23.045 3.105 ;
      RECT 22.875 5.655 23.045 5.825 ;
      RECT 22.415 0.215 22.585 0.385 ;
      RECT 22.415 2.935 22.585 3.105 ;
      RECT 22.415 5.655 22.585 5.825 ;
      RECT 22.36 1.405 22.53 1.575 ;
      RECT 22.015 4.485 22.185 4.655 ;
      RECT 21.955 2.935 22.125 3.105 ;
      RECT 21.955 5.655 22.125 5.825 ;
      RECT 21.495 2.935 21.665 3.105 ;
      RECT 21.495 5.655 21.665 5.825 ;
      RECT 21.035 2.935 21.205 3.105 ;
      RECT 21.035 5.655 21.205 5.825 ;
      RECT 20.575 2.935 20.745 3.105 ;
      RECT 20.575 5.655 20.745 5.825 ;
      RECT 20.485 3.98 20.655 4.15 ;
      RECT 20.115 2.935 20.285 3.105 ;
      RECT 20.115 5.655 20.285 5.825 ;
      RECT 19.655 2.935 19.825 3.105 ;
      RECT 19.655 5.655 19.825 5.825 ;
      RECT 19.195 2.935 19.365 3.105 ;
      RECT 19.195 5.655 19.365 5.825 ;
      RECT 18.805 4.11 18.975 4.28 ;
      RECT 18.735 2.935 18.905 3.105 ;
      RECT 18.735 5.655 18.905 5.825 ;
      RECT 18.275 2.935 18.445 3.105 ;
      RECT 18.275 5.655 18.445 5.825 ;
      RECT 17.815 0.215 17.985 0.385 ;
      RECT 17.815 2.935 17.985 3.105 ;
      RECT 17.815 5.655 17.985 5.825 ;
      RECT 17.55 3.655 17.72 3.825 ;
      RECT 17.355 0.215 17.525 0.385 ;
      RECT 17.355 2.935 17.525 3.105 ;
      RECT 17.355 5.655 17.525 5.825 ;
      RECT 16.895 0.215 17.065 0.385 ;
      RECT 16.895 2.935 17.065 3.105 ;
      RECT 16.895 5.655 17.065 5.825 ;
      RECT 16.435 0.215 16.605 0.385 ;
      RECT 16.435 2.935 16.605 3.105 ;
      RECT 16.435 5.655 16.605 5.825 ;
      RECT 15.975 0.215 16.145 0.385 ;
      RECT 15.975 2.935 16.145 3.105 ;
      RECT 15.975 5.655 16.145 5.825 ;
      RECT 15.77 4.495 15.94 4.665 ;
      RECT 15.75 1.375 15.92 1.545 ;
      RECT 15.515 0.215 15.685 0.385 ;
      RECT 15.515 2.935 15.685 3.105 ;
      RECT 15.515 5.655 15.685 5.825 ;
      RECT 15.055 0.215 15.225 0.385 ;
      RECT 15.055 2.935 15.225 3.105 ;
      RECT 15.055 5.655 15.225 5.825 ;
      RECT 14.595 0.215 14.765 0.385 ;
      RECT 14.595 2.935 14.765 3.105 ;
      RECT 14.595 5.655 14.765 5.825 ;
      RECT 14.135 0.215 14.305 0.385 ;
      RECT 14.135 2.935 14.305 3.105 ;
      RECT 14.135 5.655 14.305 5.825 ;
      RECT 13.685 1.76 13.855 1.93 ;
      RECT 13.685 4.11 13.855 4.28 ;
      RECT 13.675 0.215 13.845 0.385 ;
      RECT 13.675 2.935 13.845 3.105 ;
      RECT 13.675 5.655 13.845 5.825 ;
      RECT 13.325 1.195 13.495 1.365 ;
      RECT 13.325 4.675 13.495 4.845 ;
      RECT 13.215 0.215 13.385 0.385 ;
      RECT 13.215 2.935 13.385 3.105 ;
      RECT 13.215 5.655 13.385 5.825 ;
      RECT 12.755 0.215 12.925 0.385 ;
      RECT 12.755 2.935 12.925 3.105 ;
      RECT 12.755 5.655 12.925 5.825 ;
      RECT 12.295 0.215 12.465 0.385 ;
      RECT 12.295 2.935 12.465 3.105 ;
      RECT 12.295 5.655 12.465 5.825 ;
      RECT 12.14 1.375 12.31 1.545 ;
      RECT 12.14 4.495 12.31 4.665 ;
      RECT 11.835 0.215 12.005 0.385 ;
      RECT 11.835 2.935 12.005 3.105 ;
      RECT 11.835 5.655 12.005 5.825 ;
      RECT 11.405 5.03 11.575 5.2 ;
      RECT 11.375 0.215 11.545 0.385 ;
      RECT 11.375 2.935 11.545 3.105 ;
      RECT 11.375 5.655 11.545 5.825 ;
      RECT 11.37 0.85 11.54 1.02 ;
      RECT 10.915 0.215 11.085 0.385 ;
      RECT 10.915 2.935 11.085 3.105 ;
      RECT 10.915 5.655 11.085 5.825 ;
      RECT 10.875 1.405 11.045 1.575 ;
      RECT 10.535 3.445 10.705 3.615 ;
      RECT 10.455 0.215 10.625 0.385 ;
      RECT 10.455 1.745 10.625 1.915 ;
      RECT 10.455 2.935 10.625 3.105 ;
      RECT 10.455 5.655 10.625 5.825 ;
      RECT 9.995 0.215 10.165 0.385 ;
      RECT 9.995 2.935 10.165 3.105 ;
      RECT 9.995 5.655 10.165 5.825 ;
      RECT 9.855 4.465 10.025 4.635 ;
      RECT 9.535 0.215 9.705 0.385 ;
      RECT 9.535 2.935 9.705 3.105 ;
      RECT 9.535 5.655 9.705 5.825 ;
      RECT 9.515 0.725 9.685 0.895 ;
      RECT 9.175 4.465 9.345 4.635 ;
      RECT 9.075 0.215 9.245 0.385 ;
      RECT 9.075 2.935 9.245 3.105 ;
      RECT 9.075 5.655 9.245 5.825 ;
      RECT 8.72 0.725 8.89 0.895 ;
      RECT 8.615 0.215 8.785 0.385 ;
      RECT 8.615 2.935 8.785 3.105 ;
      RECT 8.615 5.655 8.785 5.825 ;
      RECT 8.495 2.425 8.665 2.595 ;
      RECT 8.495 4.465 8.665 4.635 ;
      RECT 8.155 0.215 8.325 0.385 ;
      RECT 8.155 2.935 8.325 3.105 ;
      RECT 8.155 5.655 8.325 5.825 ;
      RECT 7.985 4.465 8.155 4.635 ;
      RECT 7.815 1.065 7.985 1.235 ;
      RECT 7.695 0.215 7.865 0.385 ;
      RECT 7.695 2.935 7.865 3.105 ;
      RECT 7.695 5.655 7.865 5.825 ;
      RECT 7.235 0.215 7.405 0.385 ;
      RECT 7.235 2.935 7.405 3.105 ;
      RECT 7.235 5.655 7.405 5.825 ;
      RECT 6.795 4.465 6.965 4.635 ;
      RECT 6.775 0.215 6.945 0.385 ;
      RECT 6.775 2.935 6.945 3.105 ;
      RECT 6.775 5.655 6.945 5.825 ;
      RECT 6.455 1.065 6.625 1.235 ;
      RECT 6.315 0.215 6.485 0.385 ;
      RECT 6.315 2.935 6.485 3.105 ;
      RECT 6.315 5.655 6.485 5.825 ;
      RECT 6.285 2.425 6.455 2.595 ;
      RECT 5.855 0.215 6.025 0.385 ;
      RECT 5.855 2.935 6.025 3.105 ;
      RECT 5.855 5.655 6.025 5.825 ;
      RECT 5.775 4.465 5.945 4.635 ;
      RECT 5.395 0.215 5.565 0.385 ;
      RECT 5.395 2.935 5.565 3.105 ;
      RECT 5.395 5.655 5.565 5.825 ;
      RECT 5.095 3.445 5.265 3.615 ;
      RECT 4.935 0.215 5.105 0.385 ;
      RECT 4.935 2.935 5.105 3.105 ;
      RECT 4.935 5.655 5.105 5.825 ;
      RECT 4.475 0.215 4.645 0.385 ;
      RECT 4.475 2.935 4.645 3.105 ;
      RECT 4.475 5.655 4.645 5.825 ;
      RECT 4.42 1.405 4.59 1.575 ;
      RECT 4.075 4.485 4.245 4.655 ;
      RECT 4.015 2.935 4.185 3.105 ;
      RECT 4.015 5.655 4.185 5.825 ;
      RECT 3.555 2.935 3.725 3.105 ;
      RECT 3.555 5.655 3.725 5.825 ;
      RECT 3.095 2.935 3.265 3.105 ;
      RECT 3.095 5.655 3.265 5.825 ;
      RECT 2.635 2.935 2.805 3.105 ;
      RECT 2.635 5.655 2.805 5.825 ;
      RECT 2.545 3.98 2.715 4.15 ;
      RECT 2.175 2.935 2.345 3.105 ;
      RECT 2.175 5.655 2.345 5.825 ;
      RECT 1.715 2.935 1.885 3.105 ;
      RECT 1.715 5.655 1.885 5.825 ;
      RECT 1.255 2.935 1.425 3.105 ;
      RECT 1.255 5.655 1.425 5.825 ;
      RECT 0.865 4.11 1.035 4.28 ;
      RECT 0.795 2.935 0.965 3.105 ;
      RECT 0.795 5.655 0.965 5.825 ;
      RECT 0.335 2.935 0.505 3.105 ;
      RECT 0.335 5.655 0.505 5.825 ;
      RECT -0.125 2.935 0.045 3.105 ;
      RECT -0.125 5.655 0.045 5.825 ;
      RECT -0.585 2.935 -0.415 3.105 ;
      RECT -0.585 5.655 -0.415 5.825 ;
      RECT -1.045 2.935 -0.875 3.105 ;
      RECT -1.045 5.655 -0.875 5.825 ;
      RECT -1.495 4.11 -1.325 4.28 ;
      RECT -1.505 2.935 -1.335 3.105 ;
      RECT -1.505 5.655 -1.335 5.825 ;
      RECT -1.855 4.675 -1.685 4.845 ;
      RECT -1.965 2.935 -1.795 3.105 ;
      RECT -1.965 5.655 -1.795 5.825 ;
      RECT -2.425 2.935 -2.255 3.105 ;
      RECT -2.425 5.655 -2.255 5.825 ;
      RECT -2.885 2.935 -2.715 3.105 ;
      RECT -2.885 5.655 -2.715 5.825 ;
      RECT -3.345 2.935 -3.175 3.105 ;
      RECT -3.345 5.655 -3.175 5.825 ;
      RECT -3.775 3.655 -3.605 3.825 ;
      RECT -3.805 2.935 -3.635 3.105 ;
      RECT -3.805 5.655 -3.635 5.825 ;
    LAYER li ;
      RECT 88.825 0.215 89.055 1.205 ;
      RECT 87.445 0.215 87.675 1.205 ;
      RECT 76.17 0.215 76.43 1.205 ;
      RECT 70.885 0.215 71.115 1.205 ;
      RECT 69.505 0.215 69.735 1.205 ;
      RECT 58.23 0.215 58.49 1.205 ;
      RECT 52.95 0.215 53.18 1.205 ;
      RECT 51.57 0.215 51.8 1.205 ;
      RECT 40.295 0.215 40.555 1.205 ;
      RECT 35.01 0.215 35.24 1.205 ;
      RECT 33.63 0.215 33.86 1.205 ;
      RECT 22.355 0.215 22.615 1.205 ;
      RECT 17.07 0.215 17.3 1.205 ;
      RECT 15.69 0.215 15.92 1.205 ;
      RECT 4.415 0.215 4.675 1.205 ;
      RECT 82.62 0.215 82.89 1.195 ;
      RECT 81.71 0.215 81.95 1.195 ;
      RECT 64.68 0.215 64.95 1.195 ;
      RECT 63.77 0.215 64.01 1.195 ;
      RECT 46.745 0.215 47.015 1.195 ;
      RECT 45.835 0.215 46.075 1.195 ;
      RECT 28.805 0.215 29.075 1.195 ;
      RECT 27.895 0.215 28.135 1.195 ;
      RECT 10.865 0.215 11.135 1.195 ;
      RECT 9.955 0.215 10.195 1.195 ;
      RECT 80.84 0.215 81.09 0.925 ;
      RECT 62.9 0.215 63.15 0.925 ;
      RECT 44.965 0.215 45.215 0.925 ;
      RECT 27.025 0.215 27.275 0.925 ;
      RECT 9.085 0.215 9.335 0.925 ;
      RECT 85.79 0.215 86.3 0.92 ;
      RECT 67.85 0.215 68.36 0.92 ;
      RECT 49.915 0.215 50.425 0.92 ;
      RECT 31.975 0.215 32.485 0.92 ;
      RECT 14.035 0.215 14.545 0.92 ;
      RECT 78.46 0.215 78.79 0.845 ;
      RECT 60.52 0.215 60.85 0.845 ;
      RECT 42.585 0.215 42.915 0.845 ;
      RECT 24.645 0.215 24.975 0.845 ;
      RECT 6.705 0.215 7.035 0.845 ;
      RECT 83.5 0.215 83.83 0.785 ;
      RECT 65.56 0.215 65.89 0.785 ;
      RECT 47.625 0.215 47.955 0.785 ;
      RECT 29.685 0.215 30.015 0.785 ;
      RECT 11.745 0.215 12.075 0.785 ;
      RECT 71.945 0.215 72.16 0.39 ;
      RECT 54.005 0.215 54.22 0.39 ;
      RECT 36.07 0.215 36.285 0.39 ;
      RECT 18.13 0.215 18.345 0.39 ;
      RECT -3.95 0.215 0.405 0.39 ;
      RECT -3.95 0.215 89.885 0.385 ;
      RECT 88.845 1.795 89.055 4.245 ;
      RECT 87.465 1.795 87.675 4.245 ;
      RECT 83.58 1.795 83.75 4.245 ;
      RECT 75.32 2.935 75.49 4.245 ;
      RECT 70.905 1.795 71.115 4.245 ;
      RECT 69.525 1.795 69.735 4.245 ;
      RECT 65.64 1.795 65.81 4.245 ;
      RECT 57.38 2.935 57.55 4.245 ;
      RECT 52.97 1.795 53.18 4.245 ;
      RECT 51.59 1.795 51.8 4.245 ;
      RECT 47.705 1.795 47.875 4.245 ;
      RECT 39.445 2.935 39.615 4.245 ;
      RECT 35.03 1.795 35.24 4.245 ;
      RECT 33.65 1.795 33.86 4.245 ;
      RECT 29.765 1.795 29.935 4.245 ;
      RECT 21.505 2.935 21.675 4.245 ;
      RECT 17.09 1.795 17.3 4.245 ;
      RECT 15.71 1.795 15.92 4.245 ;
      RECT 11.825 1.795 11.995 4.245 ;
      RECT 3.565 2.935 3.735 4.245 ;
      RECT -3.355 2.935 -3.185 4.245 ;
      RECT 79.44 2.28 79.705 3.885 ;
      RECT 61.5 2.28 61.765 3.885 ;
      RECT 43.565 2.28 43.83 3.885 ;
      RECT 25.625 2.28 25.89 3.885 ;
      RECT 7.685 2.28 7.95 3.885 ;
      RECT 86.12 2.175 86.29 3.865 ;
      RECT 72.78 2.935 72.95 3.865 ;
      RECT 68.18 2.175 68.35 3.865 ;
      RECT 54.84 2.935 55.01 3.865 ;
      RECT 50.245 2.175 50.415 3.865 ;
      RECT 36.905 2.935 37.075 3.865 ;
      RECT 32.305 2.175 32.475 3.865 ;
      RECT 18.965 2.935 19.135 3.865 ;
      RECT 14.365 2.175 14.535 3.865 ;
      RECT 1.025 2.935 1.195 3.865 ;
      RECT -0.815 2.935 -0.645 3.865 ;
      RECT 77.28 2.43 77.61 3.825 ;
      RECT 59.34 2.43 59.67 3.825 ;
      RECT 41.405 2.43 41.735 3.825 ;
      RECT 23.465 2.43 23.795 3.825 ;
      RECT 5.525 2.43 5.855 3.825 ;
      RECT 78.28 2.935 78.56 3.775 ;
      RECT 60.34 2.935 60.62 3.775 ;
      RECT 42.405 2.935 42.685 3.775 ;
      RECT 24.465 2.935 24.745 3.775 ;
      RECT 6.525 2.935 6.805 3.775 ;
      RECT 80.255 2.935 80.63 3.485 ;
      RECT 62.315 2.935 62.69 3.485 ;
      RECT 44.38 2.935 44.755 3.485 ;
      RECT 26.44 2.935 26.815 3.485 ;
      RECT 8.5 2.935 8.875 3.485 ;
      RECT -3.95 2.935 89.885 3.105 ;
      RECT 82.56 1.795 82.89 3.105 ;
      RECT 80.82 2.39 81.075 3.105 ;
      RECT 79.39 2.28 79.995 3.105 ;
      RECT 78.52 2.39 78.735 3.105 ;
      RECT 77.09 2.43 77.705 3.105 ;
      RECT 77.51 2.065 77.705 3.105 ;
      RECT 76.17 2.425 76.43 3.105 ;
      RECT 64.62 1.795 64.95 3.105 ;
      RECT 62.88 2.39 63.135 3.105 ;
      RECT 61.45 2.28 62.055 3.105 ;
      RECT 60.58 2.39 60.795 3.105 ;
      RECT 59.15 2.43 59.765 3.105 ;
      RECT 59.57 2.065 59.765 3.105 ;
      RECT 58.23 2.425 58.49 3.105 ;
      RECT 46.685 1.795 47.015 3.105 ;
      RECT 44.945 2.39 45.2 3.105 ;
      RECT 43.515 2.28 44.12 3.105 ;
      RECT 42.645 2.39 42.86 3.105 ;
      RECT 41.215 2.43 41.83 3.105 ;
      RECT 41.635 2.065 41.83 3.105 ;
      RECT 40.295 2.425 40.555 3.105 ;
      RECT 28.745 1.795 29.075 3.105 ;
      RECT 27.005 2.39 27.26 3.105 ;
      RECT 25.575 2.28 26.18 3.105 ;
      RECT 24.705 2.39 24.92 3.105 ;
      RECT 23.275 2.43 23.89 3.105 ;
      RECT 23.695 2.065 23.89 3.105 ;
      RECT 22.355 2.425 22.615 3.105 ;
      RECT 10.805 1.795 11.135 3.105 ;
      RECT 9.065 2.39 9.32 3.105 ;
      RECT 7.635 2.28 8.24 3.105 ;
      RECT 6.765 2.39 6.98 3.105 ;
      RECT 5.335 2.43 5.95 3.105 ;
      RECT 5.755 2.065 5.95 3.105 ;
      RECT 4.415 2.425 4.675 3.105 ;
      RECT 79.82 2.01 80.005 2.38 ;
      RECT 61.88 2.01 62.065 2.38 ;
      RECT 43.945 2.01 44.13 2.38 ;
      RECT 26.005 2.01 26.19 2.38 ;
      RECT 8.065 2.01 8.25 2.38 ;
      RECT 79.82 2.01 80.15 2.255 ;
      RECT 77.51 2.065 77.84 2.255 ;
      RECT 61.88 2.01 62.21 2.255 ;
      RECT 59.57 2.065 59.9 2.255 ;
      RECT 43.945 2.01 44.275 2.255 ;
      RECT 41.635 2.065 41.965 2.255 ;
      RECT 26.005 2.01 26.335 2.255 ;
      RECT 23.695 2.065 24.025 2.255 ;
      RECT 8.065 2.01 8.395 2.255 ;
      RECT 5.755 2.065 6.085 2.255 ;
      RECT -3.95 5.655 89.885 5.825 ;
      RECT 88.825 4.835 89.055 5.825 ;
      RECT 87.445 4.835 87.675 5.825 ;
      RECT 85.79 5.12 86.3 5.825 ;
      RECT 83.5 5.255 83.83 5.825 ;
      RECT 81.52 5.145 81.97 5.825 ;
      RECT 79.43 5.255 79.76 5.825 ;
      RECT 77.36 5.195 77.61 5.825 ;
      RECT 75.24 5.255 75.57 5.825 ;
      RECT 73.82 4.325 74.095 5.825 ;
      RECT 72.77 5.12 73.28 5.825 ;
      RECT 70.885 4.835 71.115 5.825 ;
      RECT 69.505 4.835 69.735 5.825 ;
      RECT 67.85 5.12 68.36 5.825 ;
      RECT 65.56 5.255 65.89 5.825 ;
      RECT 63.58 5.145 64.03 5.825 ;
      RECT 61.49 5.255 61.82 5.825 ;
      RECT 59.42 5.195 59.67 5.825 ;
      RECT 57.3 5.255 57.63 5.825 ;
      RECT 55.88 4.325 56.155 5.825 ;
      RECT 54.83 5.12 55.34 5.825 ;
      RECT 52.95 4.835 53.18 5.825 ;
      RECT 51.57 4.835 51.8 5.825 ;
      RECT 49.915 5.12 50.425 5.825 ;
      RECT 47.625 5.255 47.955 5.825 ;
      RECT 45.645 5.145 46.095 5.825 ;
      RECT 43.555 5.255 43.885 5.825 ;
      RECT 41.485 5.195 41.735 5.825 ;
      RECT 39.365 5.255 39.695 5.825 ;
      RECT 37.945 4.325 38.22 5.825 ;
      RECT 36.895 5.12 37.405 5.825 ;
      RECT 35.01 4.835 35.24 5.825 ;
      RECT 33.63 4.835 33.86 5.825 ;
      RECT 31.975 5.12 32.485 5.825 ;
      RECT 29.685 5.255 30.015 5.825 ;
      RECT 27.705 5.145 28.155 5.825 ;
      RECT 25.615 5.255 25.945 5.825 ;
      RECT 23.545 5.195 23.795 5.825 ;
      RECT 21.425 5.255 21.755 5.825 ;
      RECT 20.005 4.325 20.28 5.825 ;
      RECT 18.955 5.12 19.465 5.825 ;
      RECT 17.07 4.835 17.3 5.825 ;
      RECT 15.69 4.835 15.92 5.825 ;
      RECT 14.035 5.12 14.545 5.825 ;
      RECT 11.745 5.255 12.075 5.825 ;
      RECT 9.765 5.145 10.215 5.825 ;
      RECT 7.675 5.255 8.005 5.825 ;
      RECT 5.605 5.195 5.855 5.825 ;
      RECT 3.485 5.255 3.815 5.825 ;
      RECT 2.065 4.325 2.34 5.825 ;
      RECT 1.015 5.12 1.525 5.825 ;
      RECT -1.145 5.12 -0.635 5.825 ;
      RECT -3.435 5.255 -3.105 5.825 ;
      RECT 89.225 1.785 89.555 2.765 ;
      RECT 89.325 0.555 89.555 2.765 ;
      RECT 89.225 0.555 89.555 1.185 ;
      RECT 89.225 4.855 89.555 5.485 ;
      RECT 89.325 3.275 89.555 5.485 ;
      RECT 89.225 3.275 89.555 4.255 ;
      RECT 87.845 1.785 88.175 2.765 ;
      RECT 87.945 0.555 88.175 2.765 ;
      RECT 88.825 1.375 89.155 1.615 ;
      RECT 87.945 1.405 89.155 1.575 ;
      RECT 87.845 0.555 88.175 1.185 ;
      RECT 87.845 4.855 88.175 5.485 ;
      RECT 87.945 3.275 88.175 5.485 ;
      RECT 88.825 4.425 89.155 4.665 ;
      RECT 87.945 4.43 89.155 4.6 ;
      RECT 87.845 3.275 88.175 4.255 ;
      RECT 86.525 2.175 87.04 2.585 ;
      RECT 86.7 1.195 87.04 2.585 ;
      RECT 85.81 1.195 87.04 1.365 ;
      RECT 86.52 0.59 86.765 1.365 ;
      RECT 86.52 4.675 86.765 5.45 ;
      RECT 85.81 4.675 87.04 4.845 ;
      RECT 86.7 3.455 87.04 4.845 ;
      RECT 86.525 3.455 87.04 3.865 ;
      RECT 83.92 2.595 85.95 2.765 ;
      RECT 85.78 1.74 85.95 2.765 ;
      RECT 83.92 1.295 84.09 2.765 ;
      RECT 85.78 1.74 86.53 1.93 ;
      RECT 83.895 1.295 84.09 1.625 ;
      RECT 83.895 4.415 84.09 4.745 ;
      RECT 83.92 3.275 84.09 4.745 ;
      RECT 85.78 4.11 86.53 4.3 ;
      RECT 85.78 3.275 85.95 4.3 ;
      RECT 83.92 3.275 85.95 3.445 ;
      RECT 84.6 1.915 85.61 2.085 ;
      RECT 85.42 0.555 85.61 2.085 ;
      RECT 84.6 1.115 84.77 2.085 ;
      RECT 85.42 3.955 85.61 5.485 ;
      RECT 84.6 3.955 84.77 4.925 ;
      RECT 84.6 3.955 85.61 4.125 ;
      RECT 84.26 2.255 85.385 2.425 ;
      RECT 84.26 0.555 84.43 2.425 ;
      RECT 83.415 1.295 83.67 1.625 ;
      RECT 83.5 0.955 83.67 1.625 ;
      RECT 83.5 0.955 84.43 1.125 ;
      RECT 84.255 0.555 84.43 1.125 ;
      RECT 84.255 0.555 84.785 0.92 ;
      RECT 84.255 5.12 84.785 5.485 ;
      RECT 84.255 4.915 84.43 5.485 ;
      RECT 84.26 3.615 84.43 5.485 ;
      RECT 83.5 4.915 84.43 5.085 ;
      RECT 83.5 4.415 83.67 5.085 ;
      RECT 83.415 4.415 83.67 4.745 ;
      RECT 84.26 3.615 85.385 3.785 ;
      RECT 83.075 1.795 83.41 2.765 ;
      RECT 83.075 0.555 83.245 2.765 ;
      RECT 83.075 0.555 83.33 1.125 ;
      RECT 83.075 4.915 83.33 5.485 ;
      RECT 83.075 3.275 83.245 5.485 ;
      RECT 83.075 3.275 83.41 4.245 ;
      RECT 79.94 5.235 81.245 5.485 ;
      RECT 79.94 4.915 80.12 5.485 ;
      RECT 79.39 4.915 80.12 5.085 ;
      RECT 79.39 4.075 79.56 5.085 ;
      RECT 80.225 4.115 81.97 4.295 ;
      RECT 81.64 3.275 81.97 4.295 ;
      RECT 79.39 4.075 80.45 4.245 ;
      RECT 81.64 3.445 82.46 3.615 ;
      RECT 80.8 3.275 81.13 3.485 ;
      RECT 80.8 3.275 81.97 3.445 ;
      RECT 81.7 1.795 82.03 2.75 ;
      RECT 81.7 1.795 82.38 1.965 ;
      RECT 82.21 0.555 82.38 1.965 ;
      RECT 82.12 0.555 82.45 1.195 ;
      RECT 81.245 2.065 81.52 2.765 ;
      RECT 81.35 0.555 81.52 2.765 ;
      RECT 81.69 1.375 82.04 1.625 ;
      RECT 81.35 1.405 82.04 1.575 ;
      RECT 81.26 0.555 81.52 1.035 ;
      RECT 80.59 3.705 81.47 3.945 ;
      RECT 81.24 3.615 81.47 3.945 ;
      RECT 79.94 3.705 81.47 3.905 ;
      RECT 80.855 3.655 81.47 3.945 ;
      RECT 79.94 3.575 80.11 3.905 ;
      RECT 80.825 4.465 81.075 5.065 ;
      RECT 80.825 4.465 81.3 4.665 ;
      RECT 80.32 1.685 81.075 2.185 ;
      RECT 79.39 1.49 79.65 2.11 ;
      RECT 80.305 1.63 80.32 1.935 ;
      RECT 80.29 1.615 80.31 1.9 ;
      RECT 80.95 1.29 81.18 1.89 ;
      RECT 80.265 1.56 80.285 1.875 ;
      RECT 80.245 1.685 81.18 1.86 ;
      RECT 80.22 1.685 81.18 1.85 ;
      RECT 80.15 1.685 81.18 1.84 ;
      RECT 80.13 1.685 81.18 1.81 ;
      RECT 80.11 0.595 80.28 1.78 ;
      RECT 80.08 1.685 81.18 1.75 ;
      RECT 80.045 1.685 81.18 1.725 ;
      RECT 80.015 1.68 80.405 1.69 ;
      RECT 80.015 1.67 80.38 1.69 ;
      RECT 80.015 1.665 80.365 1.69 ;
      RECT 80.015 1.655 80.35 1.69 ;
      RECT 79.39 1.49 80.28 1.66 ;
      RECT 79.39 1.645 80.34 1.66 ;
      RECT 79.39 1.64 80.33 1.66 ;
      RECT 80.285 1.585 80.295 1.89 ;
      RECT 79.39 1.62 80.315 1.66 ;
      RECT 79.39 1.6 80.3 1.66 ;
      RECT 79.39 0.595 80.28 0.765 ;
      RECT 80.45 1.09 80.78 1.515 ;
      RECT 80.45 0.605 80.67 1.515 ;
      RECT 80.365 4.465 80.575 5.065 ;
      RECT 80.225 4.465 80.575 4.665 ;
      RECT 78.945 2.065 79.22 2.765 ;
      RECT 79.165 0.555 79.22 2.765 ;
      RECT 79.05 1.36 79.22 2.765 ;
      RECT 79.05 0.555 79.22 1.355 ;
      RECT 78.96 0.555 79.22 1.03 ;
      RECT 77.09 1.725 77.34 2.26 ;
      RECT 78.06 1.725 78.775 2.19 ;
      RECT 77.09 1.725 78.88 1.895 ;
      RECT 78.65 1.36 78.88 1.895 ;
      RECT 77.645 0.605 77.9 1.895 ;
      RECT 78.65 1.295 78.71 2.19 ;
      RECT 78.71 1.29 78.88 1.355 ;
      RECT 77.11 0.605 77.9 0.87 ;
      RECT 78.07 4.415 78.745 4.665 ;
      RECT 78.48 4.055 78.745 4.665 ;
      RECT 78.23 4.835 78.56 5.385 ;
      RECT 77.17 4.835 78.56 5.025 ;
      RECT 77.17 3.995 77.34 5.025 ;
      RECT 77.05 4.415 77.34 4.745 ;
      RECT 77.17 3.995 78.11 4.165 ;
      RECT 77.81 3.445 78.11 4.165 ;
      RECT 78.07 1.025 78.48 1.545 ;
      RECT 78.07 0.605 78.27 1.545 ;
      RECT 76.68 0.785 76.85 2.765 ;
      RECT 76.68 1.295 77.475 1.545 ;
      RECT 76.68 0.785 76.93 1.545 ;
      RECT 76.6 0.785 76.93 1.205 ;
      RECT 76.63 5.195 77.19 5.485 ;
      RECT 76.63 3.275 76.88 5.485 ;
      RECT 76.63 3.275 77.09 3.825 ;
      RECT 75.74 4.915 75.995 5.485 ;
      RECT 75.825 3.275 75.995 5.485 ;
      RECT 75.825 4.485 76 4.655 ;
      RECT 75.66 3.275 75.995 4.245 ;
      RECT 74.285 5.12 74.815 5.485 ;
      RECT 74.64 4.915 74.815 5.485 ;
      RECT 74.64 4.915 75.57 5.085 ;
      RECT 75.4 4.415 75.57 5.085 ;
      RECT 74.64 3.615 74.81 5.485 ;
      RECT 75.4 4.415 75.655 4.745 ;
      RECT 73.685 3.615 74.81 3.785 ;
      RECT 74.98 4.415 75.175 4.745 ;
      RECT 74.98 3.275 75.15 4.745 ;
      RECT 72.54 4.11 73.29 4.3 ;
      RECT 73.12 3.275 73.29 4.3 ;
      RECT 73.12 3.275 75.15 3.445 ;
      RECT 73.46 3.955 73.65 5.485 ;
      RECT 74.3 3.955 74.47 4.925 ;
      RECT 74.295 3.955 74.47 4.21 ;
      RECT 73.46 3.955 74.47 4.125 ;
      RECT 72.305 4.675 72.55 5.45 ;
      RECT 72.03 4.675 73.26 4.845 ;
      RECT 72.03 3.455 72.37 4.845 ;
      RECT 72.03 3.455 72.545 3.865 ;
      RECT 71.285 1.785 71.615 2.765 ;
      RECT 71.385 0.555 71.615 2.765 ;
      RECT 71.285 0.555 71.615 1.185 ;
      RECT 71.285 4.855 71.615 5.485 ;
      RECT 71.385 3.275 71.615 5.485 ;
      RECT 71.285 3.275 71.615 4.255 ;
      RECT 69.905 1.785 70.235 2.765 ;
      RECT 70.005 0.555 70.235 2.765 ;
      RECT 70.885 1.375 71.215 1.615 ;
      RECT 70.005 1.405 71.215 1.575 ;
      RECT 69.905 0.555 70.235 1.185 ;
      RECT 69.905 4.855 70.235 5.485 ;
      RECT 70.005 3.275 70.235 5.485 ;
      RECT 70.885 4.425 71.215 4.665 ;
      RECT 70.005 4.43 71.215 4.6 ;
      RECT 69.905 3.275 70.235 4.255 ;
      RECT 68.585 2.175 69.1 2.585 ;
      RECT 68.76 1.195 69.1 2.585 ;
      RECT 67.87 1.195 69.1 1.365 ;
      RECT 68.58 0.59 68.825 1.365 ;
      RECT 68.58 4.675 68.825 5.45 ;
      RECT 67.87 4.675 69.1 4.845 ;
      RECT 68.76 3.455 69.1 4.845 ;
      RECT 68.585 3.455 69.1 3.865 ;
      RECT 65.98 2.595 68.01 2.765 ;
      RECT 67.84 1.74 68.01 2.765 ;
      RECT 65.98 1.295 66.15 2.765 ;
      RECT 67.84 1.74 68.59 1.93 ;
      RECT 65.955 1.295 66.15 1.625 ;
      RECT 65.955 4.415 66.15 4.745 ;
      RECT 65.98 3.275 66.15 4.745 ;
      RECT 67.84 4.11 68.59 4.3 ;
      RECT 67.84 3.275 68.01 4.3 ;
      RECT 65.98 3.275 68.01 3.445 ;
      RECT 66.66 1.915 67.67 2.085 ;
      RECT 67.48 0.555 67.67 2.085 ;
      RECT 66.66 1.115 66.83 2.085 ;
      RECT 67.48 3.955 67.67 5.485 ;
      RECT 66.66 3.955 66.83 4.925 ;
      RECT 66.66 3.955 67.67 4.125 ;
      RECT 66.32 2.255 67.445 2.425 ;
      RECT 66.32 0.555 66.49 2.425 ;
      RECT 65.475 1.295 65.73 1.625 ;
      RECT 65.56 0.955 65.73 1.625 ;
      RECT 65.56 0.955 66.49 1.125 ;
      RECT 66.315 0.555 66.49 1.125 ;
      RECT 66.315 0.555 66.845 0.92 ;
      RECT 66.315 5.12 66.845 5.485 ;
      RECT 66.315 4.915 66.49 5.485 ;
      RECT 66.32 3.615 66.49 5.485 ;
      RECT 65.56 4.915 66.49 5.085 ;
      RECT 65.56 4.415 65.73 5.085 ;
      RECT 65.475 4.415 65.73 4.745 ;
      RECT 66.32 3.615 67.445 3.785 ;
      RECT 65.135 1.795 65.47 2.765 ;
      RECT 65.135 0.555 65.305 2.765 ;
      RECT 65.135 0.555 65.39 1.125 ;
      RECT 65.135 4.915 65.39 5.485 ;
      RECT 65.135 3.275 65.305 5.485 ;
      RECT 65.135 3.275 65.47 4.245 ;
      RECT 62 5.235 63.305 5.485 ;
      RECT 62 4.915 62.18 5.485 ;
      RECT 61.45 4.915 62.18 5.085 ;
      RECT 61.45 4.075 61.62 5.085 ;
      RECT 62.285 4.115 64.03 4.295 ;
      RECT 63.7 3.275 64.03 4.295 ;
      RECT 61.45 4.075 62.51 4.245 ;
      RECT 63.7 3.445 64.52 3.615 ;
      RECT 62.86 3.275 63.19 3.485 ;
      RECT 62.86 3.275 64.03 3.445 ;
      RECT 63.76 1.795 64.09 2.75 ;
      RECT 63.76 1.795 64.44 1.965 ;
      RECT 64.27 0.555 64.44 1.965 ;
      RECT 64.18 0.555 64.51 1.195 ;
      RECT 63.305 2.065 63.58 2.765 ;
      RECT 63.41 0.555 63.58 2.765 ;
      RECT 63.75 1.375 64.1 1.625 ;
      RECT 63.41 1.405 64.1 1.575 ;
      RECT 63.32 0.555 63.58 1.035 ;
      RECT 62.65 3.705 63.53 3.945 ;
      RECT 63.3 3.615 63.53 3.945 ;
      RECT 62 3.705 63.53 3.905 ;
      RECT 62.915 3.655 63.53 3.945 ;
      RECT 62 3.575 62.17 3.905 ;
      RECT 62.885 4.465 63.135 5.065 ;
      RECT 62.885 4.465 63.36 4.665 ;
      RECT 62.38 1.685 63.135 2.185 ;
      RECT 61.45 1.49 61.71 2.11 ;
      RECT 62.365 1.63 62.38 1.935 ;
      RECT 62.35 1.615 62.37 1.9 ;
      RECT 63.01 1.29 63.24 1.89 ;
      RECT 62.325 1.56 62.345 1.875 ;
      RECT 62.305 1.685 63.24 1.86 ;
      RECT 62.28 1.685 63.24 1.85 ;
      RECT 62.21 1.685 63.24 1.84 ;
      RECT 62.19 1.685 63.24 1.81 ;
      RECT 62.17 0.595 62.34 1.78 ;
      RECT 62.14 1.685 63.24 1.75 ;
      RECT 62.105 1.685 63.24 1.725 ;
      RECT 62.075 1.68 62.465 1.69 ;
      RECT 62.075 1.67 62.44 1.69 ;
      RECT 62.075 1.665 62.425 1.69 ;
      RECT 62.075 1.655 62.41 1.69 ;
      RECT 61.45 1.49 62.34 1.66 ;
      RECT 61.45 1.645 62.4 1.66 ;
      RECT 61.45 1.64 62.39 1.66 ;
      RECT 62.345 1.585 62.355 1.89 ;
      RECT 61.45 1.62 62.375 1.66 ;
      RECT 61.45 1.6 62.36 1.66 ;
      RECT 61.45 0.595 62.34 0.765 ;
      RECT 62.51 1.09 62.84 1.515 ;
      RECT 62.51 0.605 62.73 1.515 ;
      RECT 62.425 4.465 62.635 5.065 ;
      RECT 62.285 4.465 62.635 4.665 ;
      RECT 61.005 2.065 61.28 2.765 ;
      RECT 61.225 0.555 61.28 2.765 ;
      RECT 61.11 1.36 61.28 2.765 ;
      RECT 61.11 0.555 61.28 1.355 ;
      RECT 61.02 0.555 61.28 1.03 ;
      RECT 59.15 1.725 59.4 2.26 ;
      RECT 60.12 1.725 60.835 2.19 ;
      RECT 59.15 1.725 60.94 1.895 ;
      RECT 60.71 1.36 60.94 1.895 ;
      RECT 59.705 0.605 59.96 1.895 ;
      RECT 60.71 1.295 60.77 2.19 ;
      RECT 60.77 1.29 60.94 1.355 ;
      RECT 59.17 0.605 59.96 0.87 ;
      RECT 60.13 4.415 60.805 4.665 ;
      RECT 60.54 4.055 60.805 4.665 ;
      RECT 60.29 4.835 60.62 5.385 ;
      RECT 59.23 4.835 60.62 5.025 ;
      RECT 59.23 3.995 59.4 5.025 ;
      RECT 59.11 4.415 59.4 4.745 ;
      RECT 59.23 3.995 60.17 4.165 ;
      RECT 59.87 3.445 60.17 4.165 ;
      RECT 60.13 1.025 60.54 1.545 ;
      RECT 60.13 0.605 60.33 1.545 ;
      RECT 58.74 0.785 58.91 2.765 ;
      RECT 58.74 1.295 59.535 1.545 ;
      RECT 58.74 0.785 58.99 1.545 ;
      RECT 58.66 0.785 58.99 1.205 ;
      RECT 58.69 5.195 59.25 5.485 ;
      RECT 58.69 3.275 58.94 5.485 ;
      RECT 58.69 3.275 59.15 3.825 ;
      RECT 57.8 4.915 58.055 5.485 ;
      RECT 57.885 3.275 58.055 5.485 ;
      RECT 57.885 4.485 58.06 4.655 ;
      RECT 57.72 3.275 58.055 4.245 ;
      RECT 56.345 5.12 56.875 5.485 ;
      RECT 56.7 4.915 56.875 5.485 ;
      RECT 56.7 4.915 57.63 5.085 ;
      RECT 57.46 4.415 57.63 5.085 ;
      RECT 56.7 3.615 56.87 5.485 ;
      RECT 57.46 4.415 57.715 4.745 ;
      RECT 55.745 3.615 56.87 3.785 ;
      RECT 57.04 4.415 57.235 4.745 ;
      RECT 57.04 3.275 57.21 4.745 ;
      RECT 54.6 4.11 55.35 4.3 ;
      RECT 55.18 3.275 55.35 4.3 ;
      RECT 55.18 3.275 57.21 3.445 ;
      RECT 55.52 3.955 55.71 5.485 ;
      RECT 56.36 3.955 56.53 4.925 ;
      RECT 56.355 3.955 56.53 4.21 ;
      RECT 55.52 3.955 56.53 4.125 ;
      RECT 54.365 4.675 54.61 5.45 ;
      RECT 54.09 4.675 55.32 4.845 ;
      RECT 54.09 3.455 54.43 4.845 ;
      RECT 54.09 3.455 54.605 3.865 ;
      RECT 53.35 1.785 53.68 2.765 ;
      RECT 53.45 0.555 53.68 2.765 ;
      RECT 53.35 0.555 53.68 1.185 ;
      RECT 53.35 4.855 53.68 5.485 ;
      RECT 53.45 3.275 53.68 5.485 ;
      RECT 53.35 3.275 53.68 4.255 ;
      RECT 51.97 1.785 52.3 2.765 ;
      RECT 52.07 0.555 52.3 2.765 ;
      RECT 52.95 1.375 53.28 1.615 ;
      RECT 52.07 1.405 53.28 1.575 ;
      RECT 51.97 0.555 52.3 1.185 ;
      RECT 51.97 4.855 52.3 5.485 ;
      RECT 52.07 3.275 52.3 5.485 ;
      RECT 52.95 4.425 53.28 4.665 ;
      RECT 52.07 4.43 53.28 4.6 ;
      RECT 51.97 3.275 52.3 4.255 ;
      RECT 50.65 2.175 51.165 2.585 ;
      RECT 50.825 1.195 51.165 2.585 ;
      RECT 49.935 1.195 51.165 1.365 ;
      RECT 50.645 0.59 50.89 1.365 ;
      RECT 50.645 4.675 50.89 5.45 ;
      RECT 49.935 4.675 51.165 4.845 ;
      RECT 50.825 3.455 51.165 4.845 ;
      RECT 50.65 3.455 51.165 3.865 ;
      RECT 48.045 2.595 50.075 2.765 ;
      RECT 49.905 1.74 50.075 2.765 ;
      RECT 48.045 1.295 48.215 2.765 ;
      RECT 49.905 1.74 50.655 1.93 ;
      RECT 48.02 1.295 48.215 1.625 ;
      RECT 48.02 4.415 48.215 4.745 ;
      RECT 48.045 3.275 48.215 4.745 ;
      RECT 49.905 4.11 50.655 4.3 ;
      RECT 49.905 3.275 50.075 4.3 ;
      RECT 48.045 3.275 50.075 3.445 ;
      RECT 48.725 1.915 49.735 2.085 ;
      RECT 49.545 0.555 49.735 2.085 ;
      RECT 48.725 1.115 48.895 2.085 ;
      RECT 49.545 3.955 49.735 5.485 ;
      RECT 48.725 3.955 48.895 4.925 ;
      RECT 48.725 3.955 49.735 4.125 ;
      RECT 48.385 2.255 49.51 2.425 ;
      RECT 48.385 0.555 48.555 2.425 ;
      RECT 47.54 1.295 47.795 1.625 ;
      RECT 47.625 0.955 47.795 1.625 ;
      RECT 47.625 0.955 48.555 1.125 ;
      RECT 48.38 0.555 48.555 1.125 ;
      RECT 48.38 0.555 48.91 0.92 ;
      RECT 48.38 5.12 48.91 5.485 ;
      RECT 48.38 4.915 48.555 5.485 ;
      RECT 48.385 3.615 48.555 5.485 ;
      RECT 47.625 4.915 48.555 5.085 ;
      RECT 47.625 4.415 47.795 5.085 ;
      RECT 47.54 4.415 47.795 4.745 ;
      RECT 48.385 3.615 49.51 3.785 ;
      RECT 47.2 1.795 47.535 2.765 ;
      RECT 47.2 0.555 47.37 2.765 ;
      RECT 47.2 0.555 47.455 1.125 ;
      RECT 47.2 4.915 47.455 5.485 ;
      RECT 47.2 3.275 47.37 5.485 ;
      RECT 47.2 3.275 47.535 4.245 ;
      RECT 44.065 5.235 45.37 5.485 ;
      RECT 44.065 4.915 44.245 5.485 ;
      RECT 43.515 4.915 44.245 5.085 ;
      RECT 43.515 4.075 43.685 5.085 ;
      RECT 44.35 4.115 46.095 4.295 ;
      RECT 45.765 3.275 46.095 4.295 ;
      RECT 43.515 4.075 44.575 4.245 ;
      RECT 45.765 3.445 46.585 3.615 ;
      RECT 44.925 3.275 45.255 3.485 ;
      RECT 44.925 3.275 46.095 3.445 ;
      RECT 45.825 1.795 46.155 2.75 ;
      RECT 45.825 1.795 46.505 1.965 ;
      RECT 46.335 0.555 46.505 1.965 ;
      RECT 46.245 0.555 46.575 1.195 ;
      RECT 45.37 2.065 45.645 2.765 ;
      RECT 45.475 0.555 45.645 2.765 ;
      RECT 45.815 1.375 46.165 1.625 ;
      RECT 45.475 1.405 46.165 1.575 ;
      RECT 45.385 0.555 45.645 1.035 ;
      RECT 44.715 3.705 45.595 3.945 ;
      RECT 45.365 3.615 45.595 3.945 ;
      RECT 44.065 3.705 45.595 3.905 ;
      RECT 44.98 3.655 45.595 3.945 ;
      RECT 44.065 3.575 44.235 3.905 ;
      RECT 44.95 4.465 45.2 5.065 ;
      RECT 44.95 4.465 45.425 4.665 ;
      RECT 44.445 1.685 45.2 2.185 ;
      RECT 43.515 1.49 43.775 2.11 ;
      RECT 44.43 1.63 44.445 1.935 ;
      RECT 44.415 1.615 44.435 1.9 ;
      RECT 45.075 1.29 45.305 1.89 ;
      RECT 44.39 1.56 44.41 1.875 ;
      RECT 44.37 1.685 45.305 1.86 ;
      RECT 44.345 1.685 45.305 1.85 ;
      RECT 44.275 1.685 45.305 1.84 ;
      RECT 44.255 1.685 45.305 1.81 ;
      RECT 44.235 0.595 44.405 1.78 ;
      RECT 44.205 1.685 45.305 1.75 ;
      RECT 44.17 1.685 45.305 1.725 ;
      RECT 44.14 1.68 44.53 1.69 ;
      RECT 44.14 1.67 44.505 1.69 ;
      RECT 44.14 1.665 44.49 1.69 ;
      RECT 44.14 1.655 44.475 1.69 ;
      RECT 43.515 1.49 44.405 1.66 ;
      RECT 43.515 1.645 44.465 1.66 ;
      RECT 43.515 1.64 44.455 1.66 ;
      RECT 44.41 1.585 44.42 1.89 ;
      RECT 43.515 1.62 44.44 1.66 ;
      RECT 43.515 1.6 44.425 1.66 ;
      RECT 43.515 0.595 44.405 0.765 ;
      RECT 44.575 1.09 44.905 1.515 ;
      RECT 44.575 0.605 44.795 1.515 ;
      RECT 44.49 4.465 44.7 5.065 ;
      RECT 44.35 4.465 44.7 4.665 ;
      RECT 43.07 2.065 43.345 2.765 ;
      RECT 43.29 0.555 43.345 2.765 ;
      RECT 43.175 1.36 43.345 2.765 ;
      RECT 43.175 0.555 43.345 1.355 ;
      RECT 43.085 0.555 43.345 1.03 ;
      RECT 41.215 1.725 41.465 2.26 ;
      RECT 42.185 1.725 42.9 2.19 ;
      RECT 41.215 1.725 43.005 1.895 ;
      RECT 42.775 1.36 43.005 1.895 ;
      RECT 41.77 0.605 42.025 1.895 ;
      RECT 42.775 1.295 42.835 2.19 ;
      RECT 42.835 1.29 43.005 1.355 ;
      RECT 41.235 0.605 42.025 0.87 ;
      RECT 42.195 4.415 42.87 4.665 ;
      RECT 42.605 4.055 42.87 4.665 ;
      RECT 42.355 4.835 42.685 5.385 ;
      RECT 41.295 4.835 42.685 5.025 ;
      RECT 41.295 3.995 41.465 5.025 ;
      RECT 41.175 4.415 41.465 4.745 ;
      RECT 41.295 3.995 42.235 4.165 ;
      RECT 41.935 3.445 42.235 4.165 ;
      RECT 42.195 1.025 42.605 1.545 ;
      RECT 42.195 0.605 42.395 1.545 ;
      RECT 40.805 0.785 40.975 2.765 ;
      RECT 40.805 1.295 41.6 1.545 ;
      RECT 40.805 0.785 41.055 1.545 ;
      RECT 40.725 0.785 41.055 1.205 ;
      RECT 40.755 5.195 41.315 5.485 ;
      RECT 40.755 3.275 41.005 5.485 ;
      RECT 40.755 3.275 41.215 3.825 ;
      RECT 39.865 4.915 40.12 5.485 ;
      RECT 39.95 3.275 40.12 5.485 ;
      RECT 39.95 4.485 40.125 4.655 ;
      RECT 39.785 3.275 40.12 4.245 ;
      RECT 38.41 5.12 38.94 5.485 ;
      RECT 38.765 4.915 38.94 5.485 ;
      RECT 38.765 4.915 39.695 5.085 ;
      RECT 39.525 4.415 39.695 5.085 ;
      RECT 38.765 3.615 38.935 5.485 ;
      RECT 39.525 4.415 39.78 4.745 ;
      RECT 37.81 3.615 38.935 3.785 ;
      RECT 39.105 4.415 39.3 4.745 ;
      RECT 39.105 3.275 39.275 4.745 ;
      RECT 36.665 4.11 37.415 4.3 ;
      RECT 37.245 3.275 37.415 4.3 ;
      RECT 37.245 3.275 39.275 3.445 ;
      RECT 37.585 3.955 37.775 5.485 ;
      RECT 38.425 3.955 38.595 4.925 ;
      RECT 38.42 3.955 38.595 4.21 ;
      RECT 37.585 3.955 38.595 4.125 ;
      RECT 36.43 4.675 36.675 5.45 ;
      RECT 36.155 4.675 37.385 4.845 ;
      RECT 36.155 3.455 36.495 4.845 ;
      RECT 36.155 3.455 36.67 3.865 ;
      RECT 35.41 1.785 35.74 2.765 ;
      RECT 35.51 0.555 35.74 2.765 ;
      RECT 35.41 0.555 35.74 1.185 ;
      RECT 35.41 4.855 35.74 5.485 ;
      RECT 35.51 3.275 35.74 5.485 ;
      RECT 35.41 3.275 35.74 4.255 ;
      RECT 34.03 1.785 34.36 2.765 ;
      RECT 34.13 0.555 34.36 2.765 ;
      RECT 35.01 1.375 35.34 1.615 ;
      RECT 34.13 1.405 35.34 1.575 ;
      RECT 34.03 0.555 34.36 1.185 ;
      RECT 34.03 4.855 34.36 5.485 ;
      RECT 34.13 3.275 34.36 5.485 ;
      RECT 35.01 4.425 35.34 4.665 ;
      RECT 34.13 4.43 35.34 4.6 ;
      RECT 34.03 3.275 34.36 4.255 ;
      RECT 32.71 2.175 33.225 2.585 ;
      RECT 32.885 1.195 33.225 2.585 ;
      RECT 31.995 1.195 33.225 1.365 ;
      RECT 32.705 0.59 32.95 1.365 ;
      RECT 32.705 4.675 32.95 5.45 ;
      RECT 31.995 4.675 33.225 4.845 ;
      RECT 32.885 3.455 33.225 4.845 ;
      RECT 32.71 3.455 33.225 3.865 ;
      RECT 30.105 2.595 32.135 2.765 ;
      RECT 31.965 1.74 32.135 2.765 ;
      RECT 30.105 1.295 30.275 2.765 ;
      RECT 31.965 1.74 32.715 1.93 ;
      RECT 30.08 1.295 30.275 1.625 ;
      RECT 30.08 4.415 30.275 4.745 ;
      RECT 30.105 3.275 30.275 4.745 ;
      RECT 31.965 4.11 32.715 4.3 ;
      RECT 31.965 3.275 32.135 4.3 ;
      RECT 30.105 3.275 32.135 3.445 ;
      RECT 30.785 1.915 31.795 2.085 ;
      RECT 31.605 0.555 31.795 2.085 ;
      RECT 30.785 1.115 30.955 2.085 ;
      RECT 31.605 3.955 31.795 5.485 ;
      RECT 30.785 3.955 30.955 4.925 ;
      RECT 30.785 3.955 31.795 4.125 ;
      RECT 30.445 2.255 31.57 2.425 ;
      RECT 30.445 0.555 30.615 2.425 ;
      RECT 29.6 1.295 29.855 1.625 ;
      RECT 29.685 0.955 29.855 1.625 ;
      RECT 29.685 0.955 30.615 1.125 ;
      RECT 30.44 0.555 30.615 1.125 ;
      RECT 30.44 0.555 30.97 0.92 ;
      RECT 30.44 5.12 30.97 5.485 ;
      RECT 30.44 4.915 30.615 5.485 ;
      RECT 30.445 3.615 30.615 5.485 ;
      RECT 29.685 4.915 30.615 5.085 ;
      RECT 29.685 4.415 29.855 5.085 ;
      RECT 29.6 4.415 29.855 4.745 ;
      RECT 30.445 3.615 31.57 3.785 ;
      RECT 29.26 1.795 29.595 2.765 ;
      RECT 29.26 0.555 29.43 2.765 ;
      RECT 29.26 0.555 29.515 1.125 ;
      RECT 29.26 4.915 29.515 5.485 ;
      RECT 29.26 3.275 29.43 5.485 ;
      RECT 29.26 3.275 29.595 4.245 ;
      RECT 26.125 5.235 27.43 5.485 ;
      RECT 26.125 4.915 26.305 5.485 ;
      RECT 25.575 4.915 26.305 5.085 ;
      RECT 25.575 4.075 25.745 5.085 ;
      RECT 26.41 4.115 28.155 4.295 ;
      RECT 27.825 3.275 28.155 4.295 ;
      RECT 25.575 4.075 26.635 4.245 ;
      RECT 27.825 3.445 28.645 3.615 ;
      RECT 26.985 3.275 27.315 3.485 ;
      RECT 26.985 3.275 28.155 3.445 ;
      RECT 27.885 1.795 28.215 2.75 ;
      RECT 27.885 1.795 28.565 1.965 ;
      RECT 28.395 0.555 28.565 1.965 ;
      RECT 28.305 0.555 28.635 1.195 ;
      RECT 27.43 2.065 27.705 2.765 ;
      RECT 27.535 0.555 27.705 2.765 ;
      RECT 27.875 1.375 28.225 1.625 ;
      RECT 27.535 1.405 28.225 1.575 ;
      RECT 27.445 0.555 27.705 1.035 ;
      RECT 26.775 3.705 27.655 3.945 ;
      RECT 27.425 3.615 27.655 3.945 ;
      RECT 26.125 3.705 27.655 3.905 ;
      RECT 27.04 3.655 27.655 3.945 ;
      RECT 26.125 3.575 26.295 3.905 ;
      RECT 27.01 4.465 27.26 5.065 ;
      RECT 27.01 4.465 27.485 4.665 ;
      RECT 26.505 1.685 27.26 2.185 ;
      RECT 25.575 1.49 25.835 2.11 ;
      RECT 26.49 1.63 26.505 1.935 ;
      RECT 26.475 1.615 26.495 1.9 ;
      RECT 27.135 1.29 27.365 1.89 ;
      RECT 26.45 1.56 26.47 1.875 ;
      RECT 26.43 1.685 27.365 1.86 ;
      RECT 26.405 1.685 27.365 1.85 ;
      RECT 26.335 1.685 27.365 1.84 ;
      RECT 26.315 1.685 27.365 1.81 ;
      RECT 26.295 0.595 26.465 1.78 ;
      RECT 26.265 1.685 27.365 1.75 ;
      RECT 26.23 1.685 27.365 1.725 ;
      RECT 26.2 1.68 26.59 1.69 ;
      RECT 26.2 1.67 26.565 1.69 ;
      RECT 26.2 1.665 26.55 1.69 ;
      RECT 26.2 1.655 26.535 1.69 ;
      RECT 25.575 1.49 26.465 1.66 ;
      RECT 25.575 1.645 26.525 1.66 ;
      RECT 25.575 1.64 26.515 1.66 ;
      RECT 26.47 1.585 26.48 1.89 ;
      RECT 25.575 1.62 26.5 1.66 ;
      RECT 25.575 1.6 26.485 1.66 ;
      RECT 25.575 0.595 26.465 0.765 ;
      RECT 26.635 1.09 26.965 1.515 ;
      RECT 26.635 0.605 26.855 1.515 ;
      RECT 26.55 4.465 26.76 5.065 ;
      RECT 26.41 4.465 26.76 4.665 ;
      RECT 25.13 2.065 25.405 2.765 ;
      RECT 25.35 0.555 25.405 2.765 ;
      RECT 25.235 1.36 25.405 2.765 ;
      RECT 25.235 0.555 25.405 1.355 ;
      RECT 25.145 0.555 25.405 1.03 ;
      RECT 23.275 1.725 23.525 2.26 ;
      RECT 24.245 1.725 24.96 2.19 ;
      RECT 23.275 1.725 25.065 1.895 ;
      RECT 24.835 1.36 25.065 1.895 ;
      RECT 23.83 0.605 24.085 1.895 ;
      RECT 24.835 1.295 24.895 2.19 ;
      RECT 24.895 1.29 25.065 1.355 ;
      RECT 23.295 0.605 24.085 0.87 ;
      RECT 24.255 4.415 24.93 4.665 ;
      RECT 24.665 4.055 24.93 4.665 ;
      RECT 24.415 4.835 24.745 5.385 ;
      RECT 23.355 4.835 24.745 5.025 ;
      RECT 23.355 3.995 23.525 5.025 ;
      RECT 23.235 4.415 23.525 4.745 ;
      RECT 23.355 3.995 24.295 4.165 ;
      RECT 23.995 3.445 24.295 4.165 ;
      RECT 24.255 1.025 24.665 1.545 ;
      RECT 24.255 0.605 24.455 1.545 ;
      RECT 22.865 0.785 23.035 2.765 ;
      RECT 22.865 1.295 23.66 1.545 ;
      RECT 22.865 0.785 23.115 1.545 ;
      RECT 22.785 0.785 23.115 1.205 ;
      RECT 22.815 5.195 23.375 5.485 ;
      RECT 22.815 3.275 23.065 5.485 ;
      RECT 22.815 3.275 23.275 3.825 ;
      RECT 21.925 4.915 22.18 5.485 ;
      RECT 22.01 3.275 22.18 5.485 ;
      RECT 22.01 4.485 22.185 4.655 ;
      RECT 21.845 3.275 22.18 4.245 ;
      RECT 20.47 5.12 21 5.485 ;
      RECT 20.825 4.915 21 5.485 ;
      RECT 20.825 4.915 21.755 5.085 ;
      RECT 21.585 4.415 21.755 5.085 ;
      RECT 20.825 3.615 20.995 5.485 ;
      RECT 21.585 4.415 21.84 4.745 ;
      RECT 19.87 3.615 20.995 3.785 ;
      RECT 21.165 4.415 21.36 4.745 ;
      RECT 21.165 3.275 21.335 4.745 ;
      RECT 18.725 4.11 19.475 4.3 ;
      RECT 19.305 3.275 19.475 4.3 ;
      RECT 19.305 3.275 21.335 3.445 ;
      RECT 19.645 3.955 19.835 5.485 ;
      RECT 20.485 3.955 20.655 4.925 ;
      RECT 20.48 3.955 20.655 4.21 ;
      RECT 19.645 3.955 20.655 4.125 ;
      RECT 18.49 4.675 18.735 5.45 ;
      RECT 18.215 4.675 19.445 4.845 ;
      RECT 18.215 3.455 18.555 4.845 ;
      RECT 18.215 3.455 18.73 3.865 ;
      RECT 17.47 1.785 17.8 2.765 ;
      RECT 17.57 0.555 17.8 2.765 ;
      RECT 17.47 0.555 17.8 1.185 ;
      RECT 17.47 4.855 17.8 5.485 ;
      RECT 17.57 3.275 17.8 5.485 ;
      RECT 17.47 3.275 17.8 4.255 ;
      RECT 16.09 1.785 16.42 2.765 ;
      RECT 16.19 0.555 16.42 2.765 ;
      RECT 17.07 1.375 17.4 1.615 ;
      RECT 16.19 1.405 17.4 1.575 ;
      RECT 16.09 0.555 16.42 1.185 ;
      RECT 16.09 4.855 16.42 5.485 ;
      RECT 16.19 3.275 16.42 5.485 ;
      RECT 17.07 4.425 17.4 4.665 ;
      RECT 16.19 4.43 17.4 4.6 ;
      RECT 16.09 3.275 16.42 4.255 ;
      RECT 14.77 2.175 15.285 2.585 ;
      RECT 14.945 1.195 15.285 2.585 ;
      RECT 14.055 1.195 15.285 1.365 ;
      RECT 14.765 0.59 15.01 1.365 ;
      RECT 14.765 4.675 15.01 5.45 ;
      RECT 14.055 4.675 15.285 4.845 ;
      RECT 14.945 3.455 15.285 4.845 ;
      RECT 14.77 3.455 15.285 3.865 ;
      RECT 12.165 2.595 14.195 2.765 ;
      RECT 14.025 1.74 14.195 2.765 ;
      RECT 12.165 1.295 12.335 2.765 ;
      RECT 14.025 1.74 14.775 1.93 ;
      RECT 12.14 1.295 12.335 1.625 ;
      RECT 12.14 4.415 12.335 4.745 ;
      RECT 12.165 3.275 12.335 4.745 ;
      RECT 14.025 4.11 14.775 4.3 ;
      RECT 14.025 3.275 14.195 4.3 ;
      RECT 12.165 3.275 14.195 3.445 ;
      RECT 12.845 1.915 13.855 2.085 ;
      RECT 13.665 0.555 13.855 2.085 ;
      RECT 12.845 1.115 13.015 2.085 ;
      RECT 13.665 3.955 13.855 5.485 ;
      RECT 12.845 3.955 13.015 4.925 ;
      RECT 12.845 3.955 13.855 4.125 ;
      RECT 12.505 2.255 13.63 2.425 ;
      RECT 12.505 0.555 12.675 2.425 ;
      RECT 11.66 1.295 11.915 1.625 ;
      RECT 11.745 0.955 11.915 1.625 ;
      RECT 11.745 0.955 12.675 1.125 ;
      RECT 12.5 0.555 12.675 1.125 ;
      RECT 12.5 0.555 13.03 0.92 ;
      RECT 12.5 5.12 13.03 5.485 ;
      RECT 12.5 4.915 12.675 5.485 ;
      RECT 12.505 3.615 12.675 5.485 ;
      RECT 11.745 4.915 12.675 5.085 ;
      RECT 11.745 4.415 11.915 5.085 ;
      RECT 11.66 4.415 11.915 4.745 ;
      RECT 12.505 3.615 13.63 3.785 ;
      RECT 11.32 1.795 11.655 2.765 ;
      RECT 11.32 0.555 11.49 2.765 ;
      RECT 11.32 0.555 11.575 1.125 ;
      RECT 11.32 4.915 11.575 5.485 ;
      RECT 11.32 3.275 11.49 5.485 ;
      RECT 11.32 3.275 11.655 4.245 ;
      RECT 8.185 5.235 9.49 5.485 ;
      RECT 8.185 4.915 8.365 5.485 ;
      RECT 7.635 4.915 8.365 5.085 ;
      RECT 7.635 4.075 7.805 5.085 ;
      RECT 8.47 4.115 10.215 4.295 ;
      RECT 9.885 3.275 10.215 4.295 ;
      RECT 7.635 4.075 8.695 4.245 ;
      RECT 9.885 3.445 10.705 3.615 ;
      RECT 9.045 3.275 9.375 3.485 ;
      RECT 9.045 3.275 10.215 3.445 ;
      RECT 9.945 1.795 10.275 2.75 ;
      RECT 9.945 1.795 10.625 1.965 ;
      RECT 10.455 0.555 10.625 1.965 ;
      RECT 10.365 0.555 10.695 1.195 ;
      RECT 9.49 2.065 9.765 2.765 ;
      RECT 9.595 0.555 9.765 2.765 ;
      RECT 9.935 1.375 10.285 1.625 ;
      RECT 9.595 1.405 10.285 1.575 ;
      RECT 9.505 0.555 9.765 1.035 ;
      RECT 8.835 3.705 9.715 3.945 ;
      RECT 9.485 3.615 9.715 3.945 ;
      RECT 8.185 3.705 9.715 3.905 ;
      RECT 9.1 3.655 9.715 3.945 ;
      RECT 8.185 3.575 8.355 3.905 ;
      RECT 9.07 4.465 9.32 5.065 ;
      RECT 9.07 4.465 9.545 4.665 ;
      RECT 8.565 1.685 9.32 2.185 ;
      RECT 7.635 1.49 7.895 2.11 ;
      RECT 8.55 1.63 8.565 1.935 ;
      RECT 8.535 1.615 8.555 1.9 ;
      RECT 9.195 1.29 9.425 1.89 ;
      RECT 8.51 1.56 8.53 1.875 ;
      RECT 8.49 1.685 9.425 1.86 ;
      RECT 8.465 1.685 9.425 1.85 ;
      RECT 8.395 1.685 9.425 1.84 ;
      RECT 8.375 1.685 9.425 1.81 ;
      RECT 8.355 0.595 8.525 1.78 ;
      RECT 8.325 1.685 9.425 1.75 ;
      RECT 8.29 1.685 9.425 1.725 ;
      RECT 8.26 1.68 8.65 1.69 ;
      RECT 8.26 1.67 8.625 1.69 ;
      RECT 8.26 1.665 8.61 1.69 ;
      RECT 8.26 1.655 8.595 1.69 ;
      RECT 7.635 1.49 8.525 1.66 ;
      RECT 7.635 1.645 8.585 1.66 ;
      RECT 7.635 1.64 8.575 1.66 ;
      RECT 8.53 1.585 8.54 1.89 ;
      RECT 7.635 1.62 8.56 1.66 ;
      RECT 7.635 1.6 8.545 1.66 ;
      RECT 7.635 0.595 8.525 0.765 ;
      RECT 8.695 1.09 9.025 1.515 ;
      RECT 8.695 0.605 8.915 1.515 ;
      RECT 8.61 4.465 8.82 5.065 ;
      RECT 8.47 4.465 8.82 4.665 ;
      RECT 7.19 2.065 7.465 2.765 ;
      RECT 7.41 0.555 7.465 2.765 ;
      RECT 7.295 1.36 7.465 2.765 ;
      RECT 7.295 0.555 7.465 1.355 ;
      RECT 7.205 0.555 7.465 1.03 ;
      RECT 5.335 1.725 5.585 2.26 ;
      RECT 6.305 1.725 7.02 2.19 ;
      RECT 5.335 1.725 7.125 1.895 ;
      RECT 6.895 1.36 7.125 1.895 ;
      RECT 5.89 0.605 6.145 1.895 ;
      RECT 6.895 1.295 6.955 2.19 ;
      RECT 6.955 1.29 7.125 1.355 ;
      RECT 5.355 0.605 6.145 0.87 ;
      RECT 6.315 4.415 6.99 4.665 ;
      RECT 6.725 4.055 6.99 4.665 ;
      RECT 6.475 4.835 6.805 5.385 ;
      RECT 5.415 4.835 6.805 5.025 ;
      RECT 5.415 3.995 5.585 5.025 ;
      RECT 5.295 4.415 5.585 4.745 ;
      RECT 5.415 3.995 6.355 4.165 ;
      RECT 6.055 3.445 6.355 4.165 ;
      RECT 6.315 1.025 6.725 1.545 ;
      RECT 6.315 0.605 6.515 1.545 ;
      RECT 4.925 0.785 5.095 2.765 ;
      RECT 4.925 1.295 5.72 1.545 ;
      RECT 4.925 0.785 5.175 1.545 ;
      RECT 4.845 0.785 5.175 1.205 ;
      RECT 4.875 5.195 5.435 5.485 ;
      RECT 4.875 3.275 5.125 5.485 ;
      RECT 4.875 3.275 5.335 3.825 ;
      RECT 3.985 4.915 4.24 5.485 ;
      RECT 4.07 3.275 4.24 5.485 ;
      RECT 4.07 4.485 4.245 4.655 ;
      RECT 3.905 3.275 4.24 4.245 ;
      RECT 2.53 5.12 3.06 5.485 ;
      RECT 2.885 4.915 3.06 5.485 ;
      RECT 2.885 4.915 3.815 5.085 ;
      RECT 3.645 4.415 3.815 5.085 ;
      RECT 2.885 3.615 3.055 5.485 ;
      RECT 3.645 4.415 3.9 4.745 ;
      RECT 1.93 3.615 3.055 3.785 ;
      RECT 3.225 4.415 3.42 4.745 ;
      RECT 3.225 3.275 3.395 4.745 ;
      RECT 0.785 4.11 1.535 4.3 ;
      RECT 1.365 3.275 1.535 4.3 ;
      RECT 1.365 3.275 3.395 3.445 ;
      RECT 1.705 3.955 1.895 5.485 ;
      RECT 2.545 3.955 2.715 4.925 ;
      RECT 2.54 3.955 2.715 4.21 ;
      RECT 1.705 3.955 2.715 4.125 ;
      RECT 0.55 4.675 0.795 5.45 ;
      RECT 0.275 4.675 1.505 4.845 ;
      RECT 0.275 3.455 0.615 4.845 ;
      RECT 0.275 3.455 0.79 3.865 ;
      RECT -0.415 4.675 -0.17 5.45 ;
      RECT -1.125 4.675 0.105 4.845 ;
      RECT -0.235 3.455 0.105 4.845 ;
      RECT -0.41 3.455 0.105 3.865 ;
      RECT -3.04 4.415 -2.845 4.745 ;
      RECT -3.015 3.275 -2.845 4.745 ;
      RECT -1.155 4.11 -0.405 4.3 ;
      RECT -1.155 3.275 -0.985 4.3 ;
      RECT -3.015 3.275 -0.985 3.445 ;
      RECT -1.515 3.955 -1.325 5.485 ;
      RECT -2.335 3.955 -2.165 4.925 ;
      RECT -2.335 3.955 -1.325 4.125 ;
      RECT -2.68 5.12 -2.15 5.485 ;
      RECT -2.68 4.915 -2.505 5.485 ;
      RECT -2.675 3.615 -2.505 5.485 ;
      RECT -3.435 4.915 -2.505 5.085 ;
      RECT -3.435 4.415 -3.265 5.085 ;
      RECT -3.52 4.415 -3.265 4.745 ;
      RECT -2.675 3.615 -1.55 3.785 ;
      RECT -3.86 4.915 -3.605 5.485 ;
      RECT -3.86 3.275 -3.69 5.485 ;
      RECT -3.86 3.275 -3.525 4.245 ;
      RECT 87.445 1.375 87.775 1.615 ;
      RECT 87.445 4.425 87.775 4.665 ;
      RECT 84.975 0.555 85.25 1.715 ;
      RECT 84.975 4.325 85.25 5.485 ;
      RECT 82.55 1.375 82.9 1.625 ;
      RECT 81.49 4.465 81.94 4.975 ;
      RECT 80.17 2.425 80.65 2.765 ;
      RECT 79.73 4.415 80.055 4.745 ;
      RECT 79.39 0.935 79.94 1.32 ;
      RECT 77.875 2.425 78.35 2.765 ;
      RECT 77.51 4.415 77.85 4.665 ;
      RECT 76.17 1.375 76.51 2.255 ;
      RECT 69.505 1.375 69.835 1.615 ;
      RECT 69.505 4.425 69.835 4.665 ;
      RECT 67.035 0.555 67.31 1.715 ;
      RECT 67.035 4.325 67.31 5.485 ;
      RECT 64.61 1.375 64.96 1.625 ;
      RECT 63.55 4.465 64 4.975 ;
      RECT 62.23 2.425 62.71 2.765 ;
      RECT 61.79 4.415 62.115 4.745 ;
      RECT 61.45 0.935 62 1.32 ;
      RECT 59.935 2.425 60.41 2.765 ;
      RECT 59.57 4.415 59.91 4.665 ;
      RECT 58.23 1.375 58.57 2.255 ;
      RECT 51.57 1.375 51.9 1.615 ;
      RECT 51.57 4.425 51.9 4.665 ;
      RECT 49.1 0.555 49.375 1.715 ;
      RECT 49.1 4.325 49.375 5.485 ;
      RECT 46.675 1.375 47.025 1.625 ;
      RECT 45.615 4.465 46.065 4.975 ;
      RECT 44.295 2.425 44.775 2.765 ;
      RECT 43.855 4.415 44.18 4.745 ;
      RECT 43.515 0.935 44.065 1.32 ;
      RECT 42 2.425 42.475 2.765 ;
      RECT 41.635 4.415 41.975 4.665 ;
      RECT 40.295 1.375 40.635 2.255 ;
      RECT 33.63 1.375 33.96 1.615 ;
      RECT 33.63 4.425 33.96 4.665 ;
      RECT 31.16 0.555 31.435 1.715 ;
      RECT 31.16 4.325 31.435 5.485 ;
      RECT 28.735 1.375 29.085 1.625 ;
      RECT 27.675 4.465 28.125 4.975 ;
      RECT 26.355 2.425 26.835 2.765 ;
      RECT 25.915 4.415 26.24 4.745 ;
      RECT 25.575 0.935 26.125 1.32 ;
      RECT 24.06 2.425 24.535 2.765 ;
      RECT 23.695 4.415 24.035 4.665 ;
      RECT 22.355 1.375 22.695 2.255 ;
      RECT 15.69 1.375 16.02 1.615 ;
      RECT 15.69 4.425 16.02 4.665 ;
      RECT 13.22 0.555 13.495 1.715 ;
      RECT 13.22 4.325 13.495 5.485 ;
      RECT 10.795 1.375 11.145 1.625 ;
      RECT 9.735 4.465 10.185 4.975 ;
      RECT 8.415 2.425 8.895 2.765 ;
      RECT 7.975 4.415 8.3 4.745 ;
      RECT 7.635 0.935 8.185 1.32 ;
      RECT 6.12 2.425 6.595 2.765 ;
      RECT 5.755 4.415 6.095 4.665 ;
      RECT 4.415 1.375 4.755 2.255 ;
      RECT -1.96 4.325 -1.685 5.485 ;
  END
END sky130_osu_ring_oscillator_mpr2ca_8_b0r1

END LIBRARY
