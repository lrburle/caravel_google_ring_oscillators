VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO b0r1_aa
  CLASS BLOCK ;
  FOREIGN b0r1_aa ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 50.000 ;
  PIN X1_Y1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 5.480 150.000 6.080 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 15.000 150.000 15.600 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 24.520 150.000 25.120 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 34.040 150.000 34.640 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 43.560 150.000 44.160 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 14.810 46.000 15.090 50.000 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 44.710 46.000 44.990 50.000 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 74.610 46.000 74.890 50.000 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 104.510 46.000 104.790 50.000 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 134.410 46.000 134.690 50.000 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.085 10.640 23.685 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.815 10.640 58.415 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.545 10.640 93.145 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.275 10.640 127.875 38.320 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.450 10.640 41.050 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.180 10.640 75.780 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.910 10.640 110.510 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 143.640 10.640 145.240 38.320 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 144.440 38.165 ;
      LAYER met1 ;
        RECT 4.670 10.640 145.240 38.320 ;
      LAYER met2 ;
        RECT 4.690 45.720 14.530 46.650 ;
        RECT 15.370 45.720 44.430 46.650 ;
        RECT 45.270 45.720 74.330 46.650 ;
        RECT 75.170 45.720 104.230 46.650 ;
        RECT 105.070 45.720 134.130 46.650 ;
        RECT 134.970 45.720 145.210 46.650 ;
        RECT 4.690 5.595 145.210 45.720 ;
      LAYER met3 ;
        RECT 4.000 43.160 145.600 44.025 ;
        RECT 4.000 35.040 146.000 43.160 ;
        RECT 4.000 33.640 145.600 35.040 ;
        RECT 4.000 25.520 146.000 33.640 ;
        RECT 4.400 24.120 145.600 25.520 ;
        RECT 4.000 16.000 146.000 24.120 ;
        RECT 4.000 14.600 145.600 16.000 ;
        RECT 4.000 6.480 146.000 14.600 ;
        RECT 4.000 5.615 145.600 6.480 ;
  END
END b0r1_aa
END LIBRARY

