magic
tech sky130A
magscale 1 2
timestamp 1698721842
<< obsli1 >>
rect 1104 2159 138828 85425
<< obsm1 >>
rect 1104 2128 139090 85456
<< obsm2 >>
rect 1582 2139 139086 85445
<< metal3 >>
rect 139200 85144 140000 85264
rect 139200 80792 140000 80912
rect 139200 76440 140000 76560
rect 139200 72088 140000 72208
rect 139200 67736 140000 67856
rect 139200 63384 140000 63504
rect 139200 59032 140000 59152
rect 139200 54680 140000 54800
rect 139200 50328 140000 50448
rect 139200 45976 140000 46096
rect 0 43800 800 43920
rect 139200 41624 140000 41744
rect 139200 37272 140000 37392
rect 139200 32920 140000 33040
rect 139200 28568 140000 28688
rect 139200 24216 140000 24336
rect 139200 19864 140000 19984
rect 139200 15512 140000 15632
rect 139200 11160 140000 11280
rect 139200 6808 140000 6928
rect 139200 2456 140000 2576
<< obsm3 >>
rect 798 85344 139200 85441
rect 798 85064 139120 85344
rect 798 80992 139200 85064
rect 798 80712 139120 80992
rect 798 76640 139200 80712
rect 798 76360 139120 76640
rect 798 72288 139200 76360
rect 798 72008 139120 72288
rect 798 67936 139200 72008
rect 798 67656 139120 67936
rect 798 63584 139200 67656
rect 798 63304 139120 63584
rect 798 59232 139200 63304
rect 798 58952 139120 59232
rect 798 54880 139200 58952
rect 798 54600 139120 54880
rect 798 50528 139200 54600
rect 798 50248 139120 50528
rect 798 46176 139200 50248
rect 798 45896 139120 46176
rect 798 44000 139200 45896
rect 880 43720 139200 44000
rect 798 41824 139200 43720
rect 798 41544 139120 41824
rect 798 37472 139200 41544
rect 798 37192 139120 37472
rect 798 33120 139200 37192
rect 798 32840 139120 33120
rect 798 28768 139200 32840
rect 798 28488 139120 28768
rect 798 24416 139200 28488
rect 798 24136 139120 24416
rect 798 20064 139200 24136
rect 798 19784 139120 20064
rect 798 15712 139200 19784
rect 798 15432 139120 15712
rect 798 11360 139200 15432
rect 798 11080 139120 11360
rect 798 7008 139200 11080
rect 798 6728 139120 7008
rect 798 2656 139200 6728
rect 798 2376 139120 2656
rect 798 2143 139200 2376
<< metal4 >>
rect 4208 2128 4528 85456
rect 19568 2128 19888 85456
rect 34928 2128 35248 85456
rect 50288 2128 50608 85456
rect 65648 2128 65968 85456
rect 81008 2128 81328 85456
rect 96368 2128 96688 85456
rect 111728 2128 112048 85456
rect 127088 2128 127408 85456
<< labels >>
rlabel metal3 s 139200 2456 140000 2576 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 139200 45976 140000 46096 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 139200 50328 140000 50448 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 139200 54680 140000 54800 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 139200 59032 140000 59152 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 139200 63384 140000 63504 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 139200 67736 140000 67856 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 139200 72088 140000 72208 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 139200 76440 140000 76560 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 139200 80792 140000 80912 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 139200 85144 140000 85264 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 139200 6808 140000 6928 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 139200 11160 140000 11280 6 io_in[2]
port 13 nsew signal input
rlabel metal3 s 139200 15512 140000 15632 6 io_in[3]
port 14 nsew signal input
rlabel metal3 s 139200 19864 140000 19984 6 io_in[4]
port 15 nsew signal input
rlabel metal3 s 139200 24216 140000 24336 6 io_in[5]
port 16 nsew signal input
rlabel metal3 s 139200 28568 140000 28688 6 io_in[6]
port 17 nsew signal input
rlabel metal3 s 139200 32920 140000 33040 6 io_in[7]
port 18 nsew signal input
rlabel metal3 s 139200 37272 140000 37392 6 io_in[8]
port 19 nsew signal input
rlabel metal3 s 139200 41624 140000 41744 6 io_in[9]
port 20 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 io_out
port 21 nsew signal output
rlabel metal4 s 4208 2128 4528 85456 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 85456 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 85456 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 85456 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 85456 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 85456 6 vssd1
port 23 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 85456 6 vssd1
port 23 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 85456 6 vssd1
port 23 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 85456 6 vssd1
port 23 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 140000 88000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3247952
string GDS_FILE /home/lburleson/OSU/google_ring_oscillator/caravel/openlane/mux16x1_project/runs/23_10_30_22_09/results/signoff/mux16x1_project.magic.gds
string GDS_START 140006
<< end >>

