VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_osu_ring_oscillator_mpr2ca_8_b0r1
  CLASS BLOCK ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ca_8_b0r1 ;
  ORIGIN 0.025 0.000 ;
  SIZE 85.755 BY 8.880 ;
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 3.445 5.945 3.615 7.220 ;
        RECT 14.670 5.945 14.840 7.220 ;
        RECT 14.670 1.660 14.840 2.935 ;
      LAYER mcon ;
        RECT 14.670 2.765 14.840 2.935 ;
      LAYER met1 ;
        RECT 3.385 6.115 3.675 6.145 ;
        RECT 5.665 6.115 6.005 6.170 ;
        RECT 3.385 5.945 6.005 6.115 ;
        RECT 3.385 5.915 3.675 5.945 ;
        RECT 5.665 5.890 6.005 5.945 ;
        RECT 14.595 6.115 14.920 6.190 ;
        RECT 14.595 5.945 15.070 6.115 ;
        RECT 14.595 5.865 14.920 5.945 ;
        RECT 14.590 3.635 14.915 3.960 ;
        RECT 14.665 2.965 14.845 3.635 ;
        RECT 14.610 2.935 14.900 2.965 ;
        RECT 14.610 2.765 15.070 2.935 ;
        RECT 14.610 2.735 14.900 2.765 ;
      LAYER via ;
        RECT 5.695 5.890 5.975 6.170 ;
        RECT 14.630 5.895 14.890 6.155 ;
        RECT 14.625 3.665 14.885 3.925 ;
      LAYER met2 ;
        RECT 5.750 7.885 14.835 8.055 ;
        RECT 5.750 6.200 5.920 7.885 ;
        RECT 5.695 5.860 5.975 6.200 ;
        RECT 14.660 6.190 14.835 7.885 ;
        RECT 14.595 5.865 14.920 6.190 ;
        RECT 14.660 3.960 14.835 5.865 ;
        RECT 14.590 3.635 14.915 3.960 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 20.030 5.945 20.200 7.220 ;
        RECT 31.255 5.945 31.425 7.220 ;
        RECT 31.255 1.660 31.425 2.935 ;
      LAYER mcon ;
        RECT 31.255 2.765 31.425 2.935 ;
      LAYER met1 ;
        RECT 19.970 6.115 20.260 6.145 ;
        RECT 22.250 6.115 22.590 6.170 ;
        RECT 19.970 5.945 22.590 6.115 ;
        RECT 19.970 5.915 20.260 5.945 ;
        RECT 22.250 5.890 22.590 5.945 ;
        RECT 31.180 6.115 31.505 6.190 ;
        RECT 31.180 5.945 31.655 6.115 ;
        RECT 31.180 5.865 31.505 5.945 ;
        RECT 31.175 3.635 31.500 3.960 ;
        RECT 31.250 2.965 31.430 3.635 ;
        RECT 31.195 2.935 31.485 2.965 ;
        RECT 31.195 2.765 31.655 2.935 ;
        RECT 31.195 2.735 31.485 2.765 ;
      LAYER via ;
        RECT 22.280 5.890 22.560 6.170 ;
        RECT 31.215 5.895 31.475 6.155 ;
        RECT 31.210 3.665 31.470 3.925 ;
      LAYER met2 ;
        RECT 22.335 7.885 31.420 8.055 ;
        RECT 22.335 6.200 22.505 7.885 ;
        RECT 22.280 5.860 22.560 6.200 ;
        RECT 31.245 6.190 31.420 7.885 ;
        RECT 31.180 5.865 31.505 6.190 ;
        RECT 31.245 3.960 31.420 5.865 ;
        RECT 31.175 3.635 31.500 3.960 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 36.615 5.945 36.785 7.220 ;
        RECT 47.840 5.945 48.010 7.220 ;
        RECT 47.840 1.660 48.010 2.935 ;
      LAYER mcon ;
        RECT 47.840 2.765 48.010 2.935 ;
      LAYER met1 ;
        RECT 36.555 6.115 36.845 6.145 ;
        RECT 38.835 6.115 39.175 6.170 ;
        RECT 36.555 5.945 39.175 6.115 ;
        RECT 36.555 5.915 36.845 5.945 ;
        RECT 38.835 5.890 39.175 5.945 ;
        RECT 47.765 6.115 48.090 6.190 ;
        RECT 47.765 5.945 48.240 6.115 ;
        RECT 47.765 5.865 48.090 5.945 ;
        RECT 47.760 3.635 48.085 3.960 ;
        RECT 47.835 2.965 48.015 3.635 ;
        RECT 47.780 2.935 48.070 2.965 ;
        RECT 47.780 2.765 48.240 2.935 ;
        RECT 47.780 2.735 48.070 2.765 ;
      LAYER via ;
        RECT 38.865 5.890 39.145 6.170 ;
        RECT 47.800 5.895 48.060 6.155 ;
        RECT 47.795 3.665 48.055 3.925 ;
      LAYER met2 ;
        RECT 38.920 7.885 48.005 8.055 ;
        RECT 38.920 6.200 39.090 7.885 ;
        RECT 38.865 5.860 39.145 6.200 ;
        RECT 47.830 6.190 48.005 7.885 ;
        RECT 47.765 5.865 48.090 6.190 ;
        RECT 47.830 3.960 48.005 5.865 ;
        RECT 47.760 3.635 48.085 3.960 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 53.200 5.945 53.370 7.220 ;
        RECT 64.425 5.945 64.595 7.220 ;
        RECT 64.425 1.660 64.595 2.935 ;
      LAYER mcon ;
        RECT 64.425 2.765 64.595 2.935 ;
      LAYER met1 ;
        RECT 53.140 6.115 53.430 6.145 ;
        RECT 55.420 6.115 55.760 6.170 ;
        RECT 53.140 5.945 55.760 6.115 ;
        RECT 53.140 5.915 53.430 5.945 ;
        RECT 55.420 5.890 55.760 5.945 ;
        RECT 64.350 6.115 64.675 6.190 ;
        RECT 64.350 5.945 64.825 6.115 ;
        RECT 64.350 5.865 64.675 5.945 ;
        RECT 64.345 3.635 64.670 3.960 ;
        RECT 64.420 2.965 64.600 3.635 ;
        RECT 64.365 2.935 64.655 2.965 ;
        RECT 64.365 2.765 64.825 2.935 ;
        RECT 64.365 2.735 64.655 2.765 ;
      LAYER via ;
        RECT 55.450 5.890 55.730 6.170 ;
        RECT 64.385 5.895 64.645 6.155 ;
        RECT 64.380 3.665 64.640 3.925 ;
      LAYER met2 ;
        RECT 55.505 7.885 64.590 8.055 ;
        RECT 55.505 6.200 55.675 7.885 ;
        RECT 55.450 5.860 55.730 6.200 ;
        RECT 64.415 6.190 64.590 7.885 ;
        RECT 64.350 5.865 64.675 6.190 ;
        RECT 64.415 3.960 64.590 5.865 ;
        RECT 64.345 3.635 64.670 3.960 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629000 ;
    PORT
      LAYER li1 ;
        RECT 69.780 5.945 69.950 7.220 ;
        RECT 81.005 5.945 81.175 7.220 ;
        RECT 81.005 1.660 81.175 2.935 ;
      LAYER mcon ;
        RECT 81.005 2.765 81.175 2.935 ;
      LAYER met1 ;
        RECT 69.720 6.115 70.010 6.145 ;
        RECT 72.000 6.115 72.340 6.170 ;
        RECT 69.720 5.945 72.340 6.115 ;
        RECT 69.720 5.915 70.010 5.945 ;
        RECT 72.000 5.890 72.340 5.945 ;
        RECT 80.930 6.115 81.255 6.190 ;
        RECT 80.930 5.945 81.405 6.115 ;
        RECT 80.930 5.865 81.255 5.945 ;
        RECT 80.925 3.635 81.250 3.960 ;
        RECT 81.000 2.965 81.180 3.635 ;
        RECT 80.945 2.935 81.235 2.965 ;
        RECT 80.945 2.765 81.405 2.935 ;
        RECT 80.945 2.735 81.235 2.765 ;
      LAYER via ;
        RECT 72.030 5.890 72.310 6.170 ;
        RECT 80.965 5.895 81.225 6.155 ;
        RECT 80.960 3.665 81.220 3.925 ;
      LAYER met2 ;
        RECT 72.085 7.885 81.170 8.055 ;
        RECT 72.085 6.200 72.255 7.885 ;
        RECT 72.030 5.860 72.310 6.200 ;
        RECT 80.995 6.190 81.170 7.885 ;
        RECT 80.930 5.865 81.255 6.190 ;
        RECT 80.995 3.960 81.170 5.865 ;
        RECT 80.925 3.635 81.250 3.960 ;
    END
  END s5
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 85.160 2.395 85.330 3.865 ;
        RECT 85.160 0.575 85.330 1.085 ;
      LAYER mcon ;
        RECT 85.160 0.915 85.330 1.085 ;
      LAYER met1 ;
        RECT 85.100 2.365 85.390 2.595 ;
        RECT 85.160 1.115 85.330 2.365 ;
        RECT 85.100 0.885 85.390 1.115 ;
    END
  END X5_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 68.580 2.395 68.750 3.865 ;
        RECT 68.580 0.575 68.750 1.085 ;
      LAYER mcon ;
        RECT 68.580 0.915 68.750 1.085 ;
      LAYER met1 ;
        RECT 68.520 2.365 68.810 2.595 ;
        RECT 68.580 1.115 68.750 2.365 ;
        RECT 68.520 0.885 68.810 1.115 ;
    END
  END X4_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 51.995 2.395 52.165 3.865 ;
        RECT 51.995 0.575 52.165 1.085 ;
      LAYER mcon ;
        RECT 51.995 0.915 52.165 1.085 ;
      LAYER met1 ;
        RECT 51.935 2.365 52.225 2.595 ;
        RECT 51.995 1.115 52.165 2.365 ;
        RECT 51.935 0.885 52.225 1.115 ;
    END
  END X3_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 35.410 2.395 35.580 3.865 ;
        RECT 35.410 0.575 35.580 1.085 ;
      LAYER mcon ;
        RECT 35.410 0.915 35.580 1.085 ;
      LAYER met1 ;
        RECT 35.350 2.365 35.640 2.595 ;
        RECT 35.410 1.115 35.580 2.365 ;
        RECT 35.350 0.885 35.640 1.115 ;
    END
  END X2_Y1
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.479650 ;
    PORT
      LAYER li1 ;
        RECT 18.825 2.395 18.995 3.865 ;
        RECT 18.825 0.575 18.995 1.085 ;
      LAYER mcon ;
        RECT 18.825 0.915 18.995 1.085 ;
      LAYER met1 ;
        RECT 18.765 2.365 19.055 2.595 ;
        RECT 18.825 1.115 18.995 2.365 ;
        RECT 18.765 0.885 19.055 1.115 ;
    END
  END X1_Y1
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543000 ;
    PORT
      LAYER li1 ;
        RECT 0.215 5.945 0.385 7.220 ;
      LAYER met1 ;
        RECT 0.155 6.115 0.445 6.145 ;
        RECT 0.155 5.945 0.615 6.115 ;
        RECT 0.155 5.915 0.445 5.945 ;
    END
  END start
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.025 8.570 85.730 8.880 ;
        RECT 0.205 7.945 0.375 8.570 ;
        RECT 3.435 7.945 3.605 8.570 ;
        RECT 4.385 8.025 4.555 8.305 ;
        RECT 4.385 7.855 4.610 8.025 ;
        RECT 4.440 6.245 4.610 7.855 ;
        RECT 6.200 7.180 13.400 8.570 ;
        RECT 14.660 7.945 14.830 8.570 ;
        RECT 17.405 7.945 17.575 8.570 ;
        RECT 18.395 7.945 18.565 8.570 ;
        RECT 20.020 7.945 20.190 8.570 ;
        RECT 20.970 8.025 21.140 8.305 ;
        RECT 20.970 7.855 21.195 8.025 ;
        RECT 6.495 7.065 13.395 7.180 ;
        RECT 7.770 6.605 8.020 7.065 ;
        RECT 9.840 6.665 10.170 7.065 ;
        RECT 11.930 6.555 12.380 7.065 ;
        RECT 21.025 6.245 21.195 7.855 ;
        RECT 22.785 7.180 29.985 8.570 ;
        RECT 31.245 7.945 31.415 8.570 ;
        RECT 33.990 7.945 34.160 8.570 ;
        RECT 34.980 7.945 35.150 8.570 ;
        RECT 36.605 7.945 36.775 8.570 ;
        RECT 37.555 8.025 37.725 8.305 ;
        RECT 37.555 7.855 37.780 8.025 ;
        RECT 23.080 7.065 29.980 7.180 ;
        RECT 24.355 6.605 24.605 7.065 ;
        RECT 26.425 6.665 26.755 7.065 ;
        RECT 28.515 6.555 28.965 7.065 ;
        RECT 37.610 6.245 37.780 7.855 ;
        RECT 39.370 7.180 46.570 8.570 ;
        RECT 47.830 7.945 48.000 8.570 ;
        RECT 50.575 7.945 50.745 8.570 ;
        RECT 51.565 7.945 51.735 8.570 ;
        RECT 53.190 7.945 53.360 8.570 ;
        RECT 54.140 8.025 54.310 8.305 ;
        RECT 54.140 7.855 54.365 8.025 ;
        RECT 39.665 7.065 46.565 7.180 ;
        RECT 40.940 6.605 41.190 7.065 ;
        RECT 43.010 6.665 43.340 7.065 ;
        RECT 45.100 6.555 45.550 7.065 ;
        RECT 54.195 6.245 54.365 7.855 ;
        RECT 55.955 7.180 63.155 8.570 ;
        RECT 64.415 7.945 64.585 8.570 ;
        RECT 67.160 7.945 67.330 8.570 ;
        RECT 68.150 7.945 68.320 8.570 ;
        RECT 69.770 7.945 69.940 8.570 ;
        RECT 70.720 8.025 70.890 8.305 ;
        RECT 70.720 7.855 70.945 8.025 ;
        RECT 56.250 7.065 63.150 7.180 ;
        RECT 57.525 6.605 57.775 7.065 ;
        RECT 59.595 6.665 59.925 7.065 ;
        RECT 61.685 6.555 62.135 7.065 ;
        RECT 70.775 6.245 70.945 7.855 ;
        RECT 72.535 7.180 79.735 8.570 ;
        RECT 80.995 7.945 81.165 8.570 ;
        RECT 83.740 7.945 83.910 8.570 ;
        RECT 84.730 7.945 84.900 8.570 ;
        RECT 72.830 7.065 79.730 7.180 ;
        RECT 74.105 6.605 74.355 7.065 ;
        RECT 76.175 6.665 76.505 7.065 ;
        RECT 78.265 6.555 78.715 7.065 ;
        RECT 4.385 6.075 4.610 6.245 ;
        RECT 4.385 5.015 4.555 6.075 ;
        RECT 7.920 5.825 8.260 6.075 ;
        RECT 10.140 5.825 10.465 6.155 ;
        RECT 20.970 6.075 21.195 6.245 ;
        RECT 20.970 5.015 21.140 6.075 ;
        RECT 24.505 5.825 24.845 6.075 ;
        RECT 26.725 5.825 27.050 6.155 ;
        RECT 37.555 6.075 37.780 6.245 ;
        RECT 37.555 5.015 37.725 6.075 ;
        RECT 41.090 5.825 41.430 6.075 ;
        RECT 43.310 5.825 43.635 6.155 ;
        RECT 54.140 6.075 54.365 6.245 ;
        RECT 54.140 5.015 54.310 6.075 ;
        RECT 57.675 5.825 58.015 6.075 ;
        RECT 59.895 5.825 60.220 6.155 ;
        RECT 70.720 6.075 70.945 6.245 ;
        RECT 70.720 5.015 70.890 6.075 ;
        RECT 74.255 5.825 74.595 6.075 ;
        RECT 76.475 5.825 76.800 6.155 ;
      LAYER mcon ;
        RECT 0.285 8.605 0.455 8.775 ;
        RECT 0.965 8.605 1.135 8.775 ;
        RECT 1.645 8.605 1.815 8.775 ;
        RECT 2.325 8.605 2.495 8.775 ;
        RECT 3.515 8.605 3.685 8.775 ;
        RECT 4.195 8.605 4.365 8.775 ;
        RECT 4.875 8.605 5.045 8.775 ;
        RECT 5.555 8.605 5.725 8.775 ;
        RECT 14.740 8.605 14.910 8.775 ;
        RECT 15.420 8.605 15.590 8.775 ;
        RECT 16.100 8.605 16.270 8.775 ;
        RECT 16.780 8.605 16.950 8.775 ;
        RECT 17.485 8.605 17.655 8.775 ;
        RECT 18.475 8.605 18.645 8.775 ;
        RECT 20.100 8.605 20.270 8.775 ;
        RECT 20.780 8.605 20.950 8.775 ;
        RECT 21.460 8.605 21.630 8.775 ;
        RECT 22.140 8.605 22.310 8.775 ;
        RECT 31.325 8.605 31.495 8.775 ;
        RECT 32.005 8.605 32.175 8.775 ;
        RECT 32.685 8.605 32.855 8.775 ;
        RECT 33.365 8.605 33.535 8.775 ;
        RECT 34.070 8.605 34.240 8.775 ;
        RECT 35.060 8.605 35.230 8.775 ;
        RECT 36.685 8.605 36.855 8.775 ;
        RECT 37.365 8.605 37.535 8.775 ;
        RECT 38.045 8.605 38.215 8.775 ;
        RECT 38.725 8.605 38.895 8.775 ;
        RECT 47.910 8.605 48.080 8.775 ;
        RECT 48.590 8.605 48.760 8.775 ;
        RECT 49.270 8.605 49.440 8.775 ;
        RECT 49.950 8.605 50.120 8.775 ;
        RECT 50.655 8.605 50.825 8.775 ;
        RECT 51.645 8.605 51.815 8.775 ;
        RECT 53.270 8.605 53.440 8.775 ;
        RECT 53.950 8.605 54.120 8.775 ;
        RECT 54.630 8.605 54.800 8.775 ;
        RECT 55.310 8.605 55.480 8.775 ;
        RECT 64.495 8.605 64.665 8.775 ;
        RECT 65.175 8.605 65.345 8.775 ;
        RECT 65.855 8.605 66.025 8.775 ;
        RECT 66.535 8.605 66.705 8.775 ;
        RECT 67.240 8.605 67.410 8.775 ;
        RECT 68.230 8.605 68.400 8.775 ;
        RECT 69.850 8.605 70.020 8.775 ;
        RECT 70.530 8.605 70.700 8.775 ;
        RECT 71.210 8.605 71.380 8.775 ;
        RECT 71.890 8.605 72.060 8.775 ;
        RECT 81.075 8.605 81.245 8.775 ;
        RECT 81.755 8.605 81.925 8.775 ;
        RECT 82.435 8.605 82.605 8.775 ;
        RECT 83.115 8.605 83.285 8.775 ;
        RECT 83.820 8.605 83.990 8.775 ;
        RECT 84.810 8.605 84.980 8.775 ;
        RECT 6.640 7.065 6.810 7.235 ;
        RECT 7.100 7.065 7.270 7.235 ;
        RECT 7.560 7.065 7.730 7.235 ;
        RECT 8.020 7.065 8.190 7.235 ;
        RECT 8.480 7.065 8.650 7.235 ;
        RECT 8.940 7.065 9.110 7.235 ;
        RECT 9.400 7.065 9.570 7.235 ;
        RECT 9.860 7.065 10.030 7.235 ;
        RECT 10.320 7.065 10.490 7.235 ;
        RECT 10.780 7.065 10.950 7.235 ;
        RECT 11.240 7.065 11.410 7.235 ;
        RECT 11.700 7.065 11.870 7.235 ;
        RECT 12.160 7.065 12.330 7.235 ;
        RECT 12.620 7.065 12.790 7.235 ;
        RECT 13.080 7.065 13.250 7.235 ;
        RECT 4.440 6.315 4.610 6.485 ;
        RECT 23.225 7.065 23.395 7.235 ;
        RECT 23.685 7.065 23.855 7.235 ;
        RECT 24.145 7.065 24.315 7.235 ;
        RECT 24.605 7.065 24.775 7.235 ;
        RECT 25.065 7.065 25.235 7.235 ;
        RECT 25.525 7.065 25.695 7.235 ;
        RECT 25.985 7.065 26.155 7.235 ;
        RECT 26.445 7.065 26.615 7.235 ;
        RECT 26.905 7.065 27.075 7.235 ;
        RECT 27.365 7.065 27.535 7.235 ;
        RECT 27.825 7.065 27.995 7.235 ;
        RECT 28.285 7.065 28.455 7.235 ;
        RECT 28.745 7.065 28.915 7.235 ;
        RECT 29.205 7.065 29.375 7.235 ;
        RECT 29.665 7.065 29.835 7.235 ;
        RECT 21.025 6.315 21.195 6.485 ;
        RECT 39.810 7.065 39.980 7.235 ;
        RECT 40.270 7.065 40.440 7.235 ;
        RECT 40.730 7.065 40.900 7.235 ;
        RECT 41.190 7.065 41.360 7.235 ;
        RECT 41.650 7.065 41.820 7.235 ;
        RECT 42.110 7.065 42.280 7.235 ;
        RECT 42.570 7.065 42.740 7.235 ;
        RECT 43.030 7.065 43.200 7.235 ;
        RECT 43.490 7.065 43.660 7.235 ;
        RECT 43.950 7.065 44.120 7.235 ;
        RECT 44.410 7.065 44.580 7.235 ;
        RECT 44.870 7.065 45.040 7.235 ;
        RECT 45.330 7.065 45.500 7.235 ;
        RECT 45.790 7.065 45.960 7.235 ;
        RECT 46.250 7.065 46.420 7.235 ;
        RECT 37.610 6.315 37.780 6.485 ;
        RECT 56.395 7.065 56.565 7.235 ;
        RECT 56.855 7.065 57.025 7.235 ;
        RECT 57.315 7.065 57.485 7.235 ;
        RECT 57.775 7.065 57.945 7.235 ;
        RECT 58.235 7.065 58.405 7.235 ;
        RECT 58.695 7.065 58.865 7.235 ;
        RECT 59.155 7.065 59.325 7.235 ;
        RECT 59.615 7.065 59.785 7.235 ;
        RECT 60.075 7.065 60.245 7.235 ;
        RECT 60.535 7.065 60.705 7.235 ;
        RECT 60.995 7.065 61.165 7.235 ;
        RECT 61.455 7.065 61.625 7.235 ;
        RECT 61.915 7.065 62.085 7.235 ;
        RECT 62.375 7.065 62.545 7.235 ;
        RECT 62.835 7.065 63.005 7.235 ;
        RECT 54.195 6.315 54.365 6.485 ;
        RECT 72.975 7.065 73.145 7.235 ;
        RECT 73.435 7.065 73.605 7.235 ;
        RECT 73.895 7.065 74.065 7.235 ;
        RECT 74.355 7.065 74.525 7.235 ;
        RECT 74.815 7.065 74.985 7.235 ;
        RECT 75.275 7.065 75.445 7.235 ;
        RECT 75.735 7.065 75.905 7.235 ;
        RECT 76.195 7.065 76.365 7.235 ;
        RECT 76.655 7.065 76.825 7.235 ;
        RECT 77.115 7.065 77.285 7.235 ;
        RECT 77.575 7.065 77.745 7.235 ;
        RECT 78.035 7.065 78.205 7.235 ;
        RECT 78.495 7.065 78.665 7.235 ;
        RECT 78.955 7.065 79.125 7.235 ;
        RECT 79.415 7.065 79.585 7.235 ;
        RECT 70.775 6.315 70.945 6.485 ;
        RECT 7.940 5.875 8.110 6.045 ;
        RECT 10.150 5.875 10.320 6.045 ;
        RECT 24.525 5.875 24.695 6.045 ;
        RECT 26.735 5.875 26.905 6.045 ;
        RECT 41.110 5.875 41.280 6.045 ;
        RECT 43.320 5.875 43.490 6.045 ;
        RECT 57.695 5.875 57.865 6.045 ;
        RECT 59.905 5.875 60.075 6.045 ;
        RECT 74.275 5.875 74.445 6.045 ;
        RECT 76.485 5.875 76.655 6.045 ;
      LAYER met1 ;
        RECT 0.025 8.570 85.730 8.880 ;
        RECT 4.220 6.515 4.390 8.570 ;
        RECT 6.200 7.180 13.400 8.570 ;
        RECT 6.495 6.910 13.395 7.180 ;
        RECT 8.920 6.770 9.175 6.910 ;
        RECT 8.885 6.710 9.205 6.770 ;
        RECT 7.955 6.570 10.305 6.710 ;
        RECT 4.220 6.485 4.670 6.515 ;
        RECT 4.210 6.315 4.670 6.485 ;
        RECT 4.380 6.285 4.670 6.315 ;
        RECT 7.955 6.075 8.095 6.570 ;
        RECT 8.885 6.510 9.205 6.570 ;
        RECT 10.165 6.075 10.305 6.570 ;
        RECT 20.805 6.515 20.975 8.570 ;
        RECT 22.785 7.180 29.985 8.570 ;
        RECT 23.080 6.910 29.980 7.180 ;
        RECT 25.505 6.770 25.760 6.910 ;
        RECT 25.470 6.710 25.790 6.770 ;
        RECT 24.540 6.570 26.890 6.710 ;
        RECT 20.805 6.485 21.255 6.515 ;
        RECT 20.795 6.315 21.255 6.485 ;
        RECT 20.965 6.285 21.255 6.315 ;
        RECT 24.540 6.075 24.680 6.570 ;
        RECT 25.470 6.510 25.790 6.570 ;
        RECT 26.750 6.075 26.890 6.570 ;
        RECT 37.390 6.515 37.560 8.570 ;
        RECT 39.370 7.180 46.570 8.570 ;
        RECT 39.665 6.910 46.565 7.180 ;
        RECT 42.090 6.770 42.345 6.910 ;
        RECT 42.055 6.710 42.375 6.770 ;
        RECT 41.125 6.570 43.475 6.710 ;
        RECT 37.390 6.485 37.840 6.515 ;
        RECT 37.380 6.315 37.840 6.485 ;
        RECT 37.550 6.285 37.840 6.315 ;
        RECT 41.125 6.075 41.265 6.570 ;
        RECT 42.055 6.510 42.375 6.570 ;
        RECT 43.335 6.075 43.475 6.570 ;
        RECT 53.975 6.515 54.145 8.570 ;
        RECT 55.955 7.180 63.155 8.570 ;
        RECT 56.250 6.910 63.150 7.180 ;
        RECT 58.675 6.770 58.930 6.910 ;
        RECT 58.640 6.710 58.960 6.770 ;
        RECT 57.710 6.570 60.060 6.710 ;
        RECT 53.975 6.485 54.425 6.515 ;
        RECT 53.965 6.315 54.425 6.485 ;
        RECT 54.135 6.285 54.425 6.315 ;
        RECT 57.710 6.075 57.850 6.570 ;
        RECT 58.640 6.510 58.960 6.570 ;
        RECT 59.920 6.075 60.060 6.570 ;
        RECT 70.555 6.515 70.725 8.570 ;
        RECT 72.535 7.180 79.735 8.570 ;
        RECT 72.830 6.910 79.730 7.180 ;
        RECT 75.255 6.770 75.510 6.910 ;
        RECT 75.220 6.710 75.540 6.770 ;
        RECT 74.290 6.570 76.640 6.710 ;
        RECT 70.555 6.485 71.005 6.515 ;
        RECT 70.545 6.315 71.005 6.485 ;
        RECT 70.715 6.285 71.005 6.315 ;
        RECT 74.290 6.075 74.430 6.570 ;
        RECT 75.220 6.510 75.540 6.570 ;
        RECT 76.500 6.075 76.640 6.570 ;
        RECT 7.880 5.845 8.170 6.075 ;
        RECT 10.090 5.845 10.380 6.075 ;
        RECT 24.465 5.845 24.755 6.075 ;
        RECT 26.675 5.845 26.965 6.075 ;
        RECT 41.050 5.845 41.340 6.075 ;
        RECT 43.260 5.845 43.550 6.075 ;
        RECT 57.635 5.845 57.925 6.075 ;
        RECT 59.845 5.845 60.135 6.075 ;
        RECT 74.215 5.845 74.505 6.075 ;
        RECT 76.425 5.845 76.715 6.075 ;
      LAYER via ;
        RECT 8.915 6.510 9.175 6.770 ;
        RECT 25.500 6.510 25.760 6.770 ;
        RECT 42.085 6.510 42.345 6.770 ;
        RECT 58.670 6.510 58.930 6.770 ;
        RECT 75.250 6.510 75.510 6.770 ;
      LAYER met2 ;
        RECT 8.895 6.455 9.175 6.825 ;
        RECT 25.480 6.455 25.760 6.825 ;
        RECT 42.065 6.455 42.345 6.825 ;
        RECT 58.650 6.455 58.930 6.825 ;
        RECT 75.230 6.455 75.510 6.825 ;
      LAYER via2 ;
        RECT 8.895 6.500 9.175 6.780 ;
        RECT 25.480 6.500 25.760 6.780 ;
        RECT 42.065 6.500 42.345 6.780 ;
        RECT 58.650 6.500 58.930 6.780 ;
        RECT 75.230 6.500 75.510 6.780 ;
      LAYER met3 ;
        RECT 8.840 6.805 9.140 6.905 ;
        RECT 25.425 6.805 25.725 6.905 ;
        RECT 42.010 6.805 42.310 6.905 ;
        RECT 58.595 6.805 58.895 6.905 ;
        RECT 75.175 6.805 75.475 6.905 ;
        RECT 8.840 6.790 9.200 6.805 ;
        RECT 25.425 6.790 25.785 6.805 ;
        RECT 42.010 6.790 42.370 6.805 ;
        RECT 58.595 6.790 58.955 6.805 ;
        RECT 75.175 6.790 75.535 6.805 ;
        RECT 8.400 6.490 9.200 6.790 ;
        RECT 24.985 6.490 25.785 6.790 ;
        RECT 41.570 6.490 42.370 6.790 ;
        RECT 58.155 6.490 58.955 6.790 ;
        RECT 74.735 6.490 75.535 6.790 ;
        RECT 8.870 6.475 9.200 6.490 ;
        RECT 25.455 6.475 25.785 6.490 ;
        RECT 42.040 6.475 42.370 6.490 ;
        RECT 58.625 6.475 58.955 6.490 ;
        RECT 75.205 6.475 75.535 6.490 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.580 1.795 6.840 2.615 ;
        RECT 8.870 1.795 9.200 2.255 ;
        RECT 11.250 1.795 11.500 2.335 ;
        RECT 12.120 1.795 12.360 2.605 ;
        RECT 13.030 1.795 13.300 2.605 ;
        RECT 23.165 1.795 23.425 2.615 ;
        RECT 25.455 1.795 25.785 2.255 ;
        RECT 27.835 1.795 28.085 2.335 ;
        RECT 28.705 1.795 28.945 2.605 ;
        RECT 29.615 1.795 29.885 2.605 ;
        RECT 39.750 1.795 40.010 2.615 ;
        RECT 42.040 1.795 42.370 2.255 ;
        RECT 44.420 1.795 44.670 2.335 ;
        RECT 45.290 1.795 45.530 2.605 ;
        RECT 46.200 1.795 46.470 2.605 ;
        RECT 56.335 1.795 56.595 2.615 ;
        RECT 58.625 1.795 58.955 2.255 ;
        RECT 61.005 1.795 61.255 2.335 ;
        RECT 61.875 1.795 62.115 2.605 ;
        RECT 62.785 1.795 63.055 2.605 ;
        RECT 72.915 1.795 73.175 2.615 ;
        RECT 75.205 1.795 75.535 2.255 ;
        RECT 77.585 1.795 77.835 2.335 ;
        RECT 78.455 1.795 78.695 2.605 ;
        RECT 79.365 1.795 79.635 2.605 ;
        RECT 6.495 1.655 13.585 1.795 ;
        RECT 23.080 1.655 30.170 1.795 ;
        RECT 39.665 1.655 46.755 1.795 ;
        RECT 56.250 1.655 63.340 1.795 ;
        RECT 72.830 1.655 79.920 1.795 ;
        RECT 6.240 0.310 13.585 1.655 ;
        RECT 14.660 0.310 14.830 0.935 ;
        RECT 17.405 0.310 17.575 0.935 ;
        RECT 18.395 0.310 18.565 0.935 ;
        RECT 22.825 0.310 30.170 1.655 ;
        RECT 31.245 0.310 31.415 0.935 ;
        RECT 33.990 0.310 34.160 0.935 ;
        RECT 34.980 0.310 35.150 0.935 ;
        RECT 39.410 0.310 46.755 1.655 ;
        RECT 47.830 0.310 48.000 0.935 ;
        RECT 50.575 0.310 50.745 0.935 ;
        RECT 51.565 0.310 51.735 0.935 ;
        RECT 55.995 0.310 63.340 1.655 ;
        RECT 64.415 0.310 64.585 0.935 ;
        RECT 67.160 0.310 67.330 0.935 ;
        RECT 68.150 0.310 68.320 0.935 ;
        RECT 72.575 0.310 79.920 1.655 ;
        RECT 80.995 0.310 81.165 0.935 ;
        RECT 83.740 0.310 83.910 0.935 ;
        RECT 84.730 0.310 84.900 0.935 ;
        RECT 0.000 0.000 85.705 0.310 ;
      LAYER mcon ;
        RECT 6.640 1.625 6.810 1.795 ;
        RECT 7.100 1.625 7.270 1.795 ;
        RECT 7.560 1.625 7.730 1.795 ;
        RECT 8.020 1.625 8.190 1.795 ;
        RECT 8.480 1.625 8.650 1.795 ;
        RECT 8.940 1.625 9.110 1.795 ;
        RECT 9.400 1.625 9.570 1.795 ;
        RECT 9.860 1.625 10.030 1.795 ;
        RECT 10.320 1.625 10.490 1.795 ;
        RECT 10.780 1.625 10.950 1.795 ;
        RECT 11.240 1.625 11.410 1.795 ;
        RECT 11.700 1.625 11.870 1.795 ;
        RECT 12.160 1.625 12.330 1.795 ;
        RECT 12.620 1.625 12.790 1.795 ;
        RECT 13.080 1.625 13.250 1.795 ;
        RECT 23.225 1.625 23.395 1.795 ;
        RECT 23.685 1.625 23.855 1.795 ;
        RECT 24.145 1.625 24.315 1.795 ;
        RECT 24.605 1.625 24.775 1.795 ;
        RECT 25.065 1.625 25.235 1.795 ;
        RECT 25.525 1.625 25.695 1.795 ;
        RECT 25.985 1.625 26.155 1.795 ;
        RECT 26.445 1.625 26.615 1.795 ;
        RECT 26.905 1.625 27.075 1.795 ;
        RECT 27.365 1.625 27.535 1.795 ;
        RECT 27.825 1.625 27.995 1.795 ;
        RECT 28.285 1.625 28.455 1.795 ;
        RECT 28.745 1.625 28.915 1.795 ;
        RECT 29.205 1.625 29.375 1.795 ;
        RECT 29.665 1.625 29.835 1.795 ;
        RECT 39.810 1.625 39.980 1.795 ;
        RECT 40.270 1.625 40.440 1.795 ;
        RECT 40.730 1.625 40.900 1.795 ;
        RECT 41.190 1.625 41.360 1.795 ;
        RECT 41.650 1.625 41.820 1.795 ;
        RECT 42.110 1.625 42.280 1.795 ;
        RECT 42.570 1.625 42.740 1.795 ;
        RECT 43.030 1.625 43.200 1.795 ;
        RECT 43.490 1.625 43.660 1.795 ;
        RECT 43.950 1.625 44.120 1.795 ;
        RECT 44.410 1.625 44.580 1.795 ;
        RECT 44.870 1.625 45.040 1.795 ;
        RECT 45.330 1.625 45.500 1.795 ;
        RECT 45.790 1.625 45.960 1.795 ;
        RECT 46.250 1.625 46.420 1.795 ;
        RECT 56.395 1.625 56.565 1.795 ;
        RECT 56.855 1.625 57.025 1.795 ;
        RECT 57.315 1.625 57.485 1.795 ;
        RECT 57.775 1.625 57.945 1.795 ;
        RECT 58.235 1.625 58.405 1.795 ;
        RECT 58.695 1.625 58.865 1.795 ;
        RECT 59.155 1.625 59.325 1.795 ;
        RECT 59.615 1.625 59.785 1.795 ;
        RECT 60.075 1.625 60.245 1.795 ;
        RECT 60.535 1.625 60.705 1.795 ;
        RECT 60.995 1.625 61.165 1.795 ;
        RECT 61.455 1.625 61.625 1.795 ;
        RECT 61.915 1.625 62.085 1.795 ;
        RECT 62.375 1.625 62.545 1.795 ;
        RECT 62.835 1.625 63.005 1.795 ;
        RECT 72.975 1.625 73.145 1.795 ;
        RECT 73.435 1.625 73.605 1.795 ;
        RECT 73.895 1.625 74.065 1.795 ;
        RECT 74.355 1.625 74.525 1.795 ;
        RECT 74.815 1.625 74.985 1.795 ;
        RECT 75.275 1.625 75.445 1.795 ;
        RECT 75.735 1.625 75.905 1.795 ;
        RECT 76.195 1.625 76.365 1.795 ;
        RECT 76.655 1.625 76.825 1.795 ;
        RECT 77.115 1.625 77.285 1.795 ;
        RECT 77.575 1.625 77.745 1.795 ;
        RECT 78.035 1.625 78.205 1.795 ;
        RECT 78.495 1.625 78.665 1.795 ;
        RECT 78.955 1.625 79.125 1.795 ;
        RECT 79.415 1.625 79.585 1.795 ;
        RECT 14.740 0.105 14.910 0.275 ;
        RECT 15.420 0.105 15.590 0.275 ;
        RECT 16.100 0.105 16.270 0.275 ;
        RECT 16.780 0.105 16.950 0.275 ;
        RECT 17.485 0.105 17.655 0.275 ;
        RECT 18.475 0.105 18.645 0.275 ;
        RECT 31.325 0.105 31.495 0.275 ;
        RECT 32.005 0.105 32.175 0.275 ;
        RECT 32.685 0.105 32.855 0.275 ;
        RECT 33.365 0.105 33.535 0.275 ;
        RECT 34.070 0.105 34.240 0.275 ;
        RECT 35.060 0.105 35.230 0.275 ;
        RECT 47.910 0.105 48.080 0.275 ;
        RECT 48.590 0.105 48.760 0.275 ;
        RECT 49.270 0.105 49.440 0.275 ;
        RECT 49.950 0.105 50.120 0.275 ;
        RECT 50.655 0.105 50.825 0.275 ;
        RECT 51.645 0.105 51.815 0.275 ;
        RECT 64.495 0.105 64.665 0.275 ;
        RECT 65.175 0.105 65.345 0.275 ;
        RECT 65.855 0.105 66.025 0.275 ;
        RECT 66.535 0.105 66.705 0.275 ;
        RECT 67.240 0.105 67.410 0.275 ;
        RECT 68.230 0.105 68.400 0.275 ;
        RECT 81.075 0.105 81.245 0.275 ;
        RECT 81.755 0.105 81.925 0.275 ;
        RECT 82.435 0.105 82.605 0.275 ;
        RECT 83.115 0.105 83.285 0.275 ;
        RECT 83.820 0.105 83.990 0.275 ;
        RECT 84.810 0.105 84.980 0.275 ;
      LAYER met1 ;
        RECT 6.495 1.795 13.395 1.950 ;
        RECT 23.080 1.795 29.980 1.950 ;
        RECT 39.665 1.795 46.565 1.950 ;
        RECT 56.250 1.795 63.150 1.950 ;
        RECT 72.830 1.795 79.730 1.950 ;
        RECT 6.495 1.655 13.585 1.795 ;
        RECT 23.080 1.655 30.170 1.795 ;
        RECT 39.665 1.655 46.755 1.795 ;
        RECT 56.250 1.655 63.340 1.795 ;
        RECT 72.830 1.655 79.920 1.795 ;
        RECT 6.240 0.310 13.585 1.655 ;
        RECT 22.825 0.310 30.170 1.655 ;
        RECT 39.410 0.310 46.755 1.655 ;
        RECT 55.995 0.310 63.340 1.655 ;
        RECT 72.575 0.310 79.920 1.655 ;
        RECT 0.000 0.000 85.705 0.310 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT -0.015 5.845 6.285 6.455 ;
        RECT 13.670 5.845 22.870 6.455 ;
        RECT 30.255 5.845 39.455 6.455 ;
        RECT 46.840 5.845 56.040 6.455 ;
        RECT 63.425 5.845 72.620 6.455 ;
        RECT 80.005 5.845 85.700 6.455 ;
        RECT -0.015 4.770 85.700 5.845 ;
        RECT -0.025 3.015 85.700 4.770 ;
        RECT -0.025 2.420 6.290 3.015 ;
        RECT 13.670 2.425 22.875 3.015 ;
        RECT 30.255 2.425 39.460 3.015 ;
        RECT 46.840 2.425 56.045 3.015 ;
        RECT 63.425 2.425 72.625 3.015 ;
        RECT 80.005 2.425 85.700 3.015 ;
        RECT 19.360 2.420 22.875 2.425 ;
        RECT 35.945 2.420 39.460 2.425 ;
        RECT 52.530 2.420 56.045 2.425 ;
        RECT 69.110 2.420 72.625 2.425 ;
        RECT 2.775 2.415 5.750 2.420 ;
        RECT 19.360 2.415 22.335 2.420 ;
        RECT 35.945 2.415 38.920 2.420 ;
        RECT 52.530 2.415 55.505 2.420 ;
        RECT 69.110 2.415 72.085 2.420 ;
      LAYER li1 ;
        RECT 0.205 4.745 0.375 5.475 ;
        RECT 2.015 4.745 2.185 8.305 ;
        RECT 3.435 4.745 3.605 5.475 ;
        RECT 0.030 4.740 2.780 4.745 ;
        RECT 3.260 4.740 6.010 4.745 ;
        RECT 0.030 4.515 6.355 4.740 ;
        RECT 7.690 4.515 8.020 5.235 ;
        RECT 8.690 4.515 8.970 5.185 ;
        RECT 9.850 4.515 10.115 5.295 ;
        RECT 10.665 4.515 11.040 4.895 ;
        RECT 14.660 4.745 14.830 5.475 ;
        RECT 17.405 4.745 17.575 5.475 ;
        RECT 18.395 4.745 18.565 5.475 ;
        RECT 20.020 4.745 20.190 5.475 ;
        RECT 13.425 4.740 19.365 4.745 ;
        RECT 19.845 4.740 22.595 4.745 ;
        RECT 13.425 4.670 22.940 4.740 ;
        RECT 13.295 4.515 22.940 4.670 ;
        RECT 24.275 4.515 24.605 5.235 ;
        RECT 25.275 4.515 25.555 5.185 ;
        RECT 26.435 4.515 26.700 5.295 ;
        RECT 27.250 4.515 27.625 4.895 ;
        RECT 31.245 4.745 31.415 5.475 ;
        RECT 33.990 4.745 34.160 5.475 ;
        RECT 34.980 4.745 35.150 5.475 ;
        RECT 36.605 4.745 36.775 5.475 ;
        RECT 30.010 4.740 35.950 4.745 ;
        RECT 36.430 4.740 39.180 4.745 ;
        RECT 30.010 4.670 39.525 4.740 ;
        RECT 29.880 4.515 39.525 4.670 ;
        RECT 40.860 4.515 41.190 5.235 ;
        RECT 41.860 4.515 42.140 5.185 ;
        RECT 43.020 4.515 43.285 5.295 ;
        RECT 43.835 4.515 44.210 4.895 ;
        RECT 47.830 4.745 48.000 5.475 ;
        RECT 50.575 4.745 50.745 5.475 ;
        RECT 51.565 4.745 51.735 5.475 ;
        RECT 53.190 4.745 53.360 5.475 ;
        RECT 46.595 4.740 52.535 4.745 ;
        RECT 53.015 4.740 55.765 4.745 ;
        RECT 46.595 4.670 56.110 4.740 ;
        RECT 46.465 4.515 56.110 4.670 ;
        RECT 57.445 4.515 57.775 5.235 ;
        RECT 58.445 4.515 58.725 5.185 ;
        RECT 59.605 4.515 59.870 5.295 ;
        RECT 60.420 4.515 60.795 4.895 ;
        RECT 64.415 4.745 64.585 5.475 ;
        RECT 67.160 4.745 67.330 5.475 ;
        RECT 68.150 4.745 68.320 5.475 ;
        RECT 69.770 4.745 69.940 5.475 ;
        RECT 63.180 4.740 69.120 4.745 ;
        RECT 69.595 4.740 72.345 4.745 ;
        RECT 63.180 4.670 72.690 4.740 ;
        RECT 63.050 4.515 72.690 4.670 ;
        RECT 74.025 4.515 74.355 5.235 ;
        RECT 75.025 4.515 75.305 5.185 ;
        RECT 76.185 4.515 76.450 5.295 ;
        RECT 77.000 4.515 77.375 4.895 ;
        RECT 80.995 4.745 81.165 5.475 ;
        RECT 83.740 4.745 83.910 5.475 ;
        RECT 84.730 4.745 84.900 5.475 ;
        RECT 79.760 4.670 85.700 4.745 ;
        RECT 79.630 4.515 85.700 4.670 ;
        RECT 0.030 4.345 85.700 4.515 ;
        RECT 0.030 4.130 6.355 4.345 ;
        RECT 6.580 3.835 6.840 4.345 ;
        RECT 7.500 3.840 8.115 4.345 ;
        RECT 7.920 3.665 8.115 3.840 ;
        RECT 8.930 3.800 9.145 4.345 ;
        RECT 9.800 3.790 10.405 4.345 ;
        RECT 11.230 3.800 11.485 4.345 ;
        RECT 12.970 4.135 22.940 4.345 ;
        RECT 9.800 3.690 10.415 3.790 ;
        RECT 10.230 3.665 10.415 3.690 ;
        RECT 7.920 3.475 8.250 3.665 ;
        RECT 10.230 3.420 10.560 3.665 ;
        RECT 12.970 3.205 13.300 4.135 ;
        RECT 14.660 3.405 14.830 4.135 ;
        RECT 17.405 3.405 17.575 4.135 ;
        RECT 18.395 3.405 18.565 4.135 ;
        RECT 19.365 4.130 22.940 4.135 ;
        RECT 23.165 3.835 23.425 4.345 ;
        RECT 24.085 3.840 24.700 4.345 ;
        RECT 24.505 3.665 24.700 3.840 ;
        RECT 25.515 3.800 25.730 4.345 ;
        RECT 26.385 3.790 26.990 4.345 ;
        RECT 27.815 3.800 28.070 4.345 ;
        RECT 29.555 4.135 39.525 4.345 ;
        RECT 26.385 3.690 27.000 3.790 ;
        RECT 26.815 3.665 27.000 3.690 ;
        RECT 24.505 3.475 24.835 3.665 ;
        RECT 26.815 3.420 27.145 3.665 ;
        RECT 29.555 3.205 29.885 4.135 ;
        RECT 31.245 3.405 31.415 4.135 ;
        RECT 33.990 3.405 34.160 4.135 ;
        RECT 34.980 3.405 35.150 4.135 ;
        RECT 35.950 4.130 39.525 4.135 ;
        RECT 39.750 3.835 40.010 4.345 ;
        RECT 40.670 3.840 41.285 4.345 ;
        RECT 41.090 3.665 41.285 3.840 ;
        RECT 42.100 3.800 42.315 4.345 ;
        RECT 42.970 3.790 43.575 4.345 ;
        RECT 44.400 3.800 44.655 4.345 ;
        RECT 46.140 4.135 56.110 4.345 ;
        RECT 42.970 3.690 43.585 3.790 ;
        RECT 43.400 3.665 43.585 3.690 ;
        RECT 41.090 3.475 41.420 3.665 ;
        RECT 43.400 3.420 43.730 3.665 ;
        RECT 46.140 3.205 46.470 4.135 ;
        RECT 47.830 3.405 48.000 4.135 ;
        RECT 50.575 3.405 50.745 4.135 ;
        RECT 51.565 3.405 51.735 4.135 ;
        RECT 52.535 4.130 56.110 4.135 ;
        RECT 56.335 3.835 56.595 4.345 ;
        RECT 57.255 3.840 57.870 4.345 ;
        RECT 57.675 3.665 57.870 3.840 ;
        RECT 58.685 3.800 58.900 4.345 ;
        RECT 59.555 3.790 60.160 4.345 ;
        RECT 60.985 3.800 61.240 4.345 ;
        RECT 62.725 4.135 72.690 4.345 ;
        RECT 59.555 3.690 60.170 3.790 ;
        RECT 59.985 3.665 60.170 3.690 ;
        RECT 57.675 3.475 58.005 3.665 ;
        RECT 59.985 3.420 60.315 3.665 ;
        RECT 62.725 3.205 63.055 4.135 ;
        RECT 64.415 3.405 64.585 4.135 ;
        RECT 67.160 3.405 67.330 4.135 ;
        RECT 68.150 3.405 68.320 4.135 ;
        RECT 69.115 4.130 72.690 4.135 ;
        RECT 72.915 3.835 73.175 4.345 ;
        RECT 73.835 3.840 74.450 4.345 ;
        RECT 74.255 3.665 74.450 3.840 ;
        RECT 75.265 3.800 75.480 4.345 ;
        RECT 76.135 3.790 76.740 4.345 ;
        RECT 77.565 3.800 77.820 4.345 ;
        RECT 79.305 4.135 85.700 4.345 ;
        RECT 76.135 3.690 76.750 3.790 ;
        RECT 76.565 3.665 76.750 3.690 ;
        RECT 74.255 3.475 74.585 3.665 ;
        RECT 76.565 3.420 76.895 3.665 ;
        RECT 79.305 3.205 79.635 4.135 ;
        RECT 80.995 3.405 81.165 4.135 ;
        RECT 83.740 3.405 83.910 4.135 ;
        RECT 84.730 3.405 84.900 4.135 ;
      LAYER mcon ;
        RECT 2.015 6.685 2.185 6.855 ;
        RECT 2.325 4.545 2.495 4.715 ;
        RECT 5.555 4.545 5.725 4.715 ;
        RECT 16.780 4.545 16.950 4.715 ;
        RECT 17.485 4.545 17.655 4.715 ;
        RECT 18.475 4.545 18.645 4.715 ;
        RECT 22.140 4.545 22.310 4.715 ;
        RECT 33.365 4.545 33.535 4.715 ;
        RECT 34.070 4.545 34.240 4.715 ;
        RECT 35.060 4.545 35.230 4.715 ;
        RECT 38.725 4.545 38.895 4.715 ;
        RECT 49.950 4.545 50.120 4.715 ;
        RECT 50.655 4.545 50.825 4.715 ;
        RECT 51.645 4.545 51.815 4.715 ;
        RECT 55.310 4.545 55.480 4.715 ;
        RECT 66.535 4.545 66.705 4.715 ;
        RECT 67.240 4.545 67.410 4.715 ;
        RECT 68.230 4.545 68.400 4.715 ;
        RECT 71.890 4.545 72.060 4.715 ;
        RECT 83.115 4.545 83.285 4.715 ;
        RECT 83.820 4.545 83.990 4.715 ;
        RECT 84.810 4.545 84.980 4.715 ;
        RECT 6.640 4.345 6.810 4.515 ;
        RECT 7.100 4.345 7.270 4.515 ;
        RECT 7.560 4.345 7.730 4.515 ;
        RECT 8.020 4.345 8.190 4.515 ;
        RECT 8.480 4.345 8.650 4.515 ;
        RECT 8.940 4.345 9.110 4.515 ;
        RECT 9.400 4.345 9.570 4.515 ;
        RECT 9.860 4.345 10.030 4.515 ;
        RECT 10.320 4.345 10.490 4.515 ;
        RECT 10.780 4.345 10.950 4.515 ;
        RECT 11.240 4.345 11.410 4.515 ;
        RECT 11.700 4.345 11.870 4.515 ;
        RECT 12.160 4.345 12.330 4.515 ;
        RECT 12.620 4.345 12.790 4.515 ;
        RECT 13.080 4.345 13.250 4.515 ;
        RECT 23.225 4.345 23.395 4.515 ;
        RECT 23.685 4.345 23.855 4.515 ;
        RECT 24.145 4.345 24.315 4.515 ;
        RECT 24.605 4.345 24.775 4.515 ;
        RECT 25.065 4.345 25.235 4.515 ;
        RECT 25.525 4.345 25.695 4.515 ;
        RECT 25.985 4.345 26.155 4.515 ;
        RECT 26.445 4.345 26.615 4.515 ;
        RECT 26.905 4.345 27.075 4.515 ;
        RECT 27.365 4.345 27.535 4.515 ;
        RECT 27.825 4.345 27.995 4.515 ;
        RECT 28.285 4.345 28.455 4.515 ;
        RECT 28.745 4.345 28.915 4.515 ;
        RECT 29.205 4.345 29.375 4.515 ;
        RECT 29.665 4.345 29.835 4.515 ;
        RECT 39.810 4.345 39.980 4.515 ;
        RECT 40.270 4.345 40.440 4.515 ;
        RECT 40.730 4.345 40.900 4.515 ;
        RECT 41.190 4.345 41.360 4.515 ;
        RECT 41.650 4.345 41.820 4.515 ;
        RECT 42.110 4.345 42.280 4.515 ;
        RECT 42.570 4.345 42.740 4.515 ;
        RECT 43.030 4.345 43.200 4.515 ;
        RECT 43.490 4.345 43.660 4.515 ;
        RECT 43.950 4.345 44.120 4.515 ;
        RECT 44.410 4.345 44.580 4.515 ;
        RECT 44.870 4.345 45.040 4.515 ;
        RECT 45.330 4.345 45.500 4.515 ;
        RECT 45.790 4.345 45.960 4.515 ;
        RECT 46.250 4.345 46.420 4.515 ;
        RECT 56.395 4.345 56.565 4.515 ;
        RECT 56.855 4.345 57.025 4.515 ;
        RECT 57.315 4.345 57.485 4.515 ;
        RECT 57.775 4.345 57.945 4.515 ;
        RECT 58.235 4.345 58.405 4.515 ;
        RECT 58.695 4.345 58.865 4.515 ;
        RECT 59.155 4.345 59.325 4.515 ;
        RECT 59.615 4.345 59.785 4.515 ;
        RECT 60.075 4.345 60.245 4.515 ;
        RECT 60.535 4.345 60.705 4.515 ;
        RECT 60.995 4.345 61.165 4.515 ;
        RECT 61.455 4.345 61.625 4.515 ;
        RECT 61.915 4.345 62.085 4.515 ;
        RECT 62.375 4.345 62.545 4.515 ;
        RECT 62.835 4.345 63.005 4.515 ;
        RECT 72.975 4.345 73.145 4.515 ;
        RECT 73.435 4.345 73.605 4.515 ;
        RECT 73.895 4.345 74.065 4.515 ;
        RECT 74.355 4.345 74.525 4.515 ;
        RECT 74.815 4.345 74.985 4.515 ;
        RECT 75.275 4.345 75.445 4.515 ;
        RECT 75.735 4.345 75.905 4.515 ;
        RECT 76.195 4.345 76.365 4.515 ;
        RECT 76.655 4.345 76.825 4.515 ;
        RECT 77.115 4.345 77.285 4.515 ;
        RECT 77.575 4.345 77.745 4.515 ;
        RECT 78.035 4.345 78.205 4.515 ;
        RECT 78.495 4.345 78.665 4.515 ;
        RECT 78.955 4.345 79.125 4.515 ;
        RECT 79.415 4.345 79.585 4.515 ;
        RECT 16.780 4.165 16.950 4.335 ;
        RECT 17.485 4.165 17.655 4.335 ;
        RECT 18.475 4.165 18.645 4.335 ;
        RECT 33.365 4.165 33.535 4.335 ;
        RECT 34.070 4.165 34.240 4.335 ;
        RECT 35.060 4.165 35.230 4.335 ;
        RECT 49.950 4.165 50.120 4.335 ;
        RECT 50.655 4.165 50.825 4.335 ;
        RECT 51.645 4.165 51.815 4.335 ;
        RECT 66.535 4.165 66.705 4.335 ;
        RECT 67.240 4.165 67.410 4.335 ;
        RECT 68.230 4.165 68.400 4.335 ;
        RECT 83.115 4.165 83.285 4.335 ;
        RECT 83.820 4.165 83.990 4.335 ;
        RECT 84.810 4.165 84.980 4.335 ;
      LAYER met1 ;
        RECT 1.955 6.855 2.245 6.885 ;
        RECT 1.785 6.685 2.245 6.855 ;
        RECT 1.955 6.655 2.245 6.685 ;
        RECT 0.030 4.740 2.780 4.745 ;
        RECT 3.260 4.740 6.010 4.745 ;
        RECT 13.425 4.740 19.365 4.745 ;
        RECT 19.845 4.740 22.595 4.745 ;
        RECT 30.010 4.740 35.950 4.745 ;
        RECT 36.430 4.740 39.180 4.745 ;
        RECT 46.595 4.740 52.535 4.745 ;
        RECT 53.015 4.740 55.765 4.745 ;
        RECT 63.180 4.740 69.120 4.745 ;
        RECT 69.595 4.740 72.345 4.745 ;
        RECT 0.030 4.670 6.355 4.740 ;
        RECT 13.425 4.670 22.940 4.740 ;
        RECT 30.010 4.670 39.525 4.740 ;
        RECT 46.595 4.670 56.110 4.740 ;
        RECT 63.180 4.670 72.690 4.740 ;
        RECT 79.760 4.670 85.700 4.745 ;
        RECT 0.030 4.190 85.700 4.670 ;
        RECT 0.030 4.130 6.355 4.190 ;
        RECT 13.295 4.150 22.940 4.190 ;
        RECT 29.880 4.150 39.525 4.190 ;
        RECT 46.465 4.150 56.110 4.190 ;
        RECT 63.050 4.150 72.690 4.190 ;
        RECT 79.630 4.150 85.700 4.190 ;
        RECT 13.885 4.135 22.940 4.150 ;
        RECT 30.470 4.135 39.525 4.150 ;
        RECT 47.055 4.135 56.110 4.150 ;
        RECT 63.640 4.135 72.690 4.150 ;
        RECT 80.220 4.135 85.700 4.150 ;
        RECT 19.365 4.130 22.940 4.135 ;
        RECT 35.950 4.130 39.525 4.135 ;
        RECT 52.535 4.130 56.110 4.135 ;
        RECT 69.115 4.130 72.690 4.135 ;
    END
  END vccd1
  OBS
      LAYER pwell ;
        RECT 6.430 7.045 7.030 7.450 ;
        RECT 8.940 7.205 9.110 7.235 ;
        RECT 8.940 7.045 9.515 7.205 ;
        RECT 12.155 7.200 12.325 7.235 ;
        RECT 12.155 7.090 12.790 7.200 ;
        RECT 12.155 7.045 12.470 7.090 ;
        RECT 6.430 6.850 12.470 7.045 ;
        RECT 23.015 7.045 23.615 7.450 ;
        RECT 25.525 7.205 25.695 7.235 ;
        RECT 25.525 7.045 26.100 7.205 ;
        RECT 28.740 7.200 28.910 7.235 ;
        RECT 28.740 7.090 29.375 7.200 ;
        RECT 28.740 7.045 29.055 7.090 ;
        RECT 23.015 6.850 29.055 7.045 ;
        RECT 39.600 7.045 40.200 7.450 ;
        RECT 42.110 7.205 42.280 7.235 ;
        RECT 42.110 7.045 42.685 7.205 ;
        RECT 45.325 7.200 45.495 7.235 ;
        RECT 45.325 7.090 45.960 7.200 ;
        RECT 45.325 7.045 45.640 7.090 ;
        RECT 39.600 6.850 45.640 7.045 ;
        RECT 56.185 7.045 56.785 7.450 ;
        RECT 58.695 7.205 58.865 7.235 ;
        RECT 58.695 7.045 59.270 7.205 ;
        RECT 61.910 7.200 62.080 7.235 ;
        RECT 61.910 7.090 62.545 7.200 ;
        RECT 61.910 7.045 62.225 7.090 ;
        RECT 56.185 6.850 62.225 7.045 ;
        RECT 72.765 7.045 73.365 7.450 ;
        RECT 75.275 7.205 75.445 7.235 ;
        RECT 75.275 7.045 75.850 7.205 ;
        RECT 78.490 7.200 78.660 7.235 ;
        RECT 78.490 7.090 79.125 7.200 ;
        RECT 78.490 7.045 78.805 7.090 ;
        RECT 72.765 6.850 78.805 7.045 ;
        RECT 7.160 6.225 12.470 6.850 ;
        RECT 7.160 6.135 8.110 6.225 ;
        RECT 9.720 6.135 12.470 6.225 ;
        RECT 23.745 6.225 29.055 6.850 ;
        RECT 23.745 6.135 24.695 6.225 ;
        RECT 26.305 6.135 29.055 6.225 ;
        RECT 40.330 6.225 45.640 6.850 ;
        RECT 40.330 6.135 41.280 6.225 ;
        RECT 42.890 6.135 45.640 6.225 ;
        RECT 56.915 6.225 62.225 6.850 ;
        RECT 56.915 6.135 57.865 6.225 ;
        RECT 59.475 6.135 62.225 6.225 ;
        RECT 73.495 6.225 78.805 6.850 ;
        RECT 73.495 6.135 74.445 6.225 ;
        RECT 76.055 6.135 78.805 6.225 ;
        RECT 6.500 2.525 7.430 2.725 ;
        RECT 8.760 2.720 9.120 2.725 ;
        RECT 9.575 2.720 9.710 2.725 ;
        RECT 8.760 2.525 9.710 2.720 ;
        RECT 6.500 2.495 9.710 2.525 ;
        RECT 11.090 2.495 13.370 2.725 ;
        RECT 6.500 2.010 13.370 2.495 ;
        RECT 23.085 2.525 24.015 2.725 ;
        RECT 25.345 2.720 25.705 2.725 ;
        RECT 26.160 2.720 26.295 2.725 ;
        RECT 25.345 2.525 26.295 2.720 ;
        RECT 23.085 2.495 26.295 2.525 ;
        RECT 27.675 2.495 29.955 2.725 ;
        RECT 23.085 2.010 29.955 2.495 ;
        RECT 39.670 2.525 40.600 2.725 ;
        RECT 41.930 2.720 42.290 2.725 ;
        RECT 42.745 2.720 42.880 2.725 ;
        RECT 41.930 2.525 42.880 2.720 ;
        RECT 39.670 2.495 42.880 2.525 ;
        RECT 44.260 2.495 46.540 2.725 ;
        RECT 39.670 2.010 46.540 2.495 ;
        RECT 56.255 2.525 57.185 2.725 ;
        RECT 58.515 2.720 58.875 2.725 ;
        RECT 59.330 2.720 59.465 2.725 ;
        RECT 58.515 2.525 59.465 2.720 ;
        RECT 56.255 2.495 59.465 2.525 ;
        RECT 60.845 2.495 63.125 2.725 ;
        RECT 56.255 2.010 63.125 2.495 ;
        RECT 72.835 2.525 73.765 2.725 ;
        RECT 75.095 2.720 75.455 2.725 ;
        RECT 75.910 2.720 76.045 2.725 ;
        RECT 75.095 2.525 76.045 2.720 ;
        RECT 72.835 2.495 76.045 2.525 ;
        RECT 77.425 2.495 79.705 2.725 ;
        RECT 72.835 2.010 79.705 2.495 ;
        RECT 6.430 1.845 13.370 2.010 ;
        RECT 6.430 1.410 7.030 1.845 ;
        RECT 8.775 1.815 13.370 1.845 ;
        RECT 23.015 1.845 29.955 2.010 ;
        RECT 9.860 1.625 10.030 1.815 ;
        RECT 12.165 1.625 12.335 1.815 ;
        RECT 23.015 1.410 23.615 1.845 ;
        RECT 25.360 1.815 29.955 1.845 ;
        RECT 39.600 1.845 46.540 2.010 ;
        RECT 26.445 1.625 26.615 1.815 ;
        RECT 28.750 1.625 28.920 1.815 ;
        RECT 39.600 1.410 40.200 1.845 ;
        RECT 41.945 1.815 46.540 1.845 ;
        RECT 56.185 1.845 63.125 2.010 ;
        RECT 43.030 1.625 43.200 1.815 ;
        RECT 45.335 1.625 45.505 1.815 ;
        RECT 56.185 1.410 56.785 1.845 ;
        RECT 58.530 1.815 63.125 1.845 ;
        RECT 72.765 1.845 79.705 2.010 ;
        RECT 59.615 1.625 59.785 1.815 ;
        RECT 61.920 1.625 62.090 1.815 ;
        RECT 72.765 1.410 73.365 1.845 ;
        RECT 75.110 1.815 79.705 1.845 ;
        RECT 76.195 1.625 76.365 1.815 ;
        RECT 78.500 1.625 78.670 1.815 ;
      LAYER li1 ;
        RECT 0.635 7.645 0.805 8.305 ;
        RECT 1.155 8.025 1.325 8.305 ;
        RECT 1.155 7.855 1.380 8.025 ;
        RECT 0.635 7.315 1.040 7.645 ;
        RECT 0.635 6.805 0.805 7.315 ;
        RECT 0.635 6.475 1.040 6.805 ;
        RECT 0.635 5.015 0.805 6.475 ;
        RECT 1.210 6.245 1.380 7.855 ;
        RECT 1.585 7.795 1.755 8.305 ;
        RECT 3.865 7.645 4.035 8.305 ;
        RECT 4.815 7.795 4.985 8.305 ;
        RECT 3.865 7.315 4.270 7.645 ;
        RECT 1.155 6.075 1.380 6.245 ;
        RECT 1.155 5.015 1.325 6.075 ;
        RECT 1.585 5.015 1.755 7.225 ;
        RECT 3.865 6.805 4.035 7.315 ;
        RECT 3.865 6.475 4.270 6.805 ;
        RECT 3.865 5.015 4.035 6.475 ;
        RECT 4.815 5.015 4.985 7.225 ;
        RECT 5.245 5.015 5.415 8.305 ;
        RECT 15.090 7.645 15.260 8.305 ;
        RECT 15.610 8.025 15.780 8.305 ;
        RECT 15.610 7.855 15.835 8.025 ;
        RECT 15.090 7.315 15.495 7.645 ;
        RECT 7.040 6.605 7.600 6.895 ;
        RECT 7.040 5.235 7.290 6.605 ;
        RECT 8.640 6.435 8.970 6.795 ;
        RECT 10.350 6.645 11.655 6.895 ;
        RECT 15.090 6.805 15.260 7.315 ;
        RECT 10.350 6.495 10.530 6.645 ;
        RECT 7.580 6.245 8.970 6.435 ;
        RECT 9.800 6.325 10.530 6.495 ;
        RECT 15.090 6.475 15.495 6.805 ;
        RECT 7.580 6.155 7.750 6.245 ;
        RECT 7.460 5.825 7.750 6.155 ;
        RECT 8.480 5.825 9.155 6.075 ;
        RECT 7.580 5.575 7.750 5.825 ;
        RECT 7.580 5.405 8.520 5.575 ;
        RECT 8.890 5.465 9.155 5.825 ;
        RECT 9.800 5.655 9.970 6.325 ;
        RECT 10.775 6.075 10.985 6.475 ;
        RECT 10.635 5.875 10.985 6.075 ;
        RECT 11.235 6.075 11.485 6.475 ;
        RECT 11.235 5.875 11.710 6.075 ;
        RECT 11.900 5.875 12.350 6.385 ;
        RECT 10.635 5.655 12.380 5.705 ;
        RECT 9.800 5.525 12.380 5.655 ;
        RECT 9.800 5.485 10.860 5.525 ;
        RECT 7.040 4.685 7.500 5.235 ;
        RECT 8.220 4.855 8.520 5.405 ;
        RECT 11.000 5.315 11.880 5.355 ;
        RECT 10.350 5.115 11.880 5.315 ;
        RECT 10.350 4.985 10.520 5.115 ;
        RECT 11.265 5.065 11.880 5.115 ;
        RECT 11.650 5.025 11.880 5.065 ;
        RECT 12.050 5.025 12.380 5.525 ;
        RECT 11.210 4.855 11.540 4.895 ;
        RECT 12.050 4.855 12.870 5.025 ;
        RECT 15.090 5.015 15.260 6.475 ;
        RECT 15.665 6.245 15.835 7.855 ;
        RECT 16.040 7.795 16.210 8.305 ;
        RECT 15.610 6.075 15.835 6.245 ;
        RECT 15.610 5.015 15.780 6.075 ;
        RECT 16.040 5.015 16.210 7.225 ;
        RECT 16.470 5.015 16.640 8.305 ;
        RECT 17.835 7.795 18.005 8.305 ;
        RECT 18.825 7.795 18.995 8.305 ;
        RECT 20.450 7.645 20.620 8.305 ;
        RECT 21.400 7.795 21.570 8.305 ;
        RECT 20.450 7.315 20.855 7.645 ;
        RECT 17.465 6.970 17.930 7.140 ;
        RECT 18.455 6.970 18.920 7.140 ;
        RECT 17.465 5.945 17.635 6.970 ;
        RECT 17.835 5.015 18.005 6.485 ;
        RECT 18.455 5.945 18.625 6.970 ;
        RECT 20.450 6.805 20.620 7.315 ;
        RECT 18.825 5.015 18.995 6.485 ;
        RECT 20.450 6.475 20.855 6.805 ;
        RECT 20.450 5.015 20.620 6.475 ;
        RECT 21.400 5.015 21.570 7.225 ;
        RECT 21.830 5.015 22.000 8.305 ;
        RECT 31.675 7.645 31.845 8.305 ;
        RECT 32.195 8.025 32.365 8.305 ;
        RECT 32.195 7.855 32.420 8.025 ;
        RECT 31.675 7.315 32.080 7.645 ;
        RECT 23.625 6.605 24.185 6.895 ;
        RECT 23.625 5.235 23.875 6.605 ;
        RECT 25.225 6.435 25.555 6.795 ;
        RECT 26.935 6.645 28.240 6.895 ;
        RECT 31.675 6.805 31.845 7.315 ;
        RECT 26.935 6.495 27.115 6.645 ;
        RECT 24.165 6.245 25.555 6.435 ;
        RECT 26.385 6.325 27.115 6.495 ;
        RECT 31.675 6.475 32.080 6.805 ;
        RECT 24.165 6.155 24.335 6.245 ;
        RECT 24.045 5.825 24.335 6.155 ;
        RECT 25.065 5.825 25.740 6.075 ;
        RECT 24.165 5.575 24.335 5.825 ;
        RECT 24.165 5.405 25.105 5.575 ;
        RECT 25.475 5.465 25.740 5.825 ;
        RECT 26.385 5.655 26.555 6.325 ;
        RECT 27.360 6.075 27.570 6.475 ;
        RECT 27.220 5.875 27.570 6.075 ;
        RECT 27.820 6.075 28.070 6.475 ;
        RECT 27.820 5.875 28.295 6.075 ;
        RECT 28.485 5.875 28.935 6.385 ;
        RECT 27.220 5.655 28.965 5.705 ;
        RECT 26.385 5.525 28.965 5.655 ;
        RECT 26.385 5.485 27.445 5.525 ;
        RECT 11.210 4.685 12.380 4.855 ;
        RECT 23.625 4.685 24.085 5.235 ;
        RECT 24.805 4.855 25.105 5.405 ;
        RECT 27.585 5.315 28.465 5.355 ;
        RECT 26.935 5.115 28.465 5.315 ;
        RECT 26.935 4.985 27.105 5.115 ;
        RECT 27.850 5.065 28.465 5.115 ;
        RECT 28.235 5.025 28.465 5.065 ;
        RECT 28.635 5.025 28.965 5.525 ;
        RECT 27.795 4.855 28.125 4.895 ;
        RECT 28.635 4.855 29.455 5.025 ;
        RECT 31.675 5.015 31.845 6.475 ;
        RECT 32.250 6.245 32.420 7.855 ;
        RECT 32.625 7.795 32.795 8.305 ;
        RECT 32.195 6.075 32.420 6.245 ;
        RECT 32.195 5.015 32.365 6.075 ;
        RECT 32.625 5.015 32.795 7.225 ;
        RECT 33.055 5.015 33.225 8.305 ;
        RECT 34.420 7.795 34.590 8.305 ;
        RECT 35.410 7.795 35.580 8.305 ;
        RECT 37.035 7.645 37.205 8.305 ;
        RECT 37.985 7.795 38.155 8.305 ;
        RECT 37.035 7.315 37.440 7.645 ;
        RECT 34.050 6.970 34.515 7.140 ;
        RECT 35.040 6.970 35.505 7.140 ;
        RECT 34.050 5.945 34.220 6.970 ;
        RECT 34.420 5.015 34.590 6.485 ;
        RECT 35.040 5.945 35.210 6.970 ;
        RECT 37.035 6.805 37.205 7.315 ;
        RECT 35.410 5.015 35.580 6.485 ;
        RECT 37.035 6.475 37.440 6.805 ;
        RECT 37.035 5.015 37.205 6.475 ;
        RECT 37.985 5.015 38.155 7.225 ;
        RECT 38.415 5.015 38.585 8.305 ;
        RECT 48.260 7.645 48.430 8.305 ;
        RECT 48.780 8.025 48.950 8.305 ;
        RECT 48.780 7.855 49.005 8.025 ;
        RECT 48.260 7.315 48.665 7.645 ;
        RECT 40.210 6.605 40.770 6.895 ;
        RECT 40.210 5.235 40.460 6.605 ;
        RECT 41.810 6.435 42.140 6.795 ;
        RECT 43.520 6.645 44.825 6.895 ;
        RECT 48.260 6.805 48.430 7.315 ;
        RECT 43.520 6.495 43.700 6.645 ;
        RECT 40.750 6.245 42.140 6.435 ;
        RECT 42.970 6.325 43.700 6.495 ;
        RECT 48.260 6.475 48.665 6.805 ;
        RECT 40.750 6.155 40.920 6.245 ;
        RECT 40.630 5.825 40.920 6.155 ;
        RECT 41.650 5.825 42.325 6.075 ;
        RECT 40.750 5.575 40.920 5.825 ;
        RECT 40.750 5.405 41.690 5.575 ;
        RECT 42.060 5.465 42.325 5.825 ;
        RECT 42.970 5.655 43.140 6.325 ;
        RECT 43.945 6.075 44.155 6.475 ;
        RECT 43.805 5.875 44.155 6.075 ;
        RECT 44.405 6.075 44.655 6.475 ;
        RECT 44.405 5.875 44.880 6.075 ;
        RECT 45.070 5.875 45.520 6.385 ;
        RECT 43.805 5.655 45.550 5.705 ;
        RECT 42.970 5.525 45.550 5.655 ;
        RECT 42.970 5.485 44.030 5.525 ;
        RECT 27.795 4.685 28.965 4.855 ;
        RECT 40.210 4.685 40.670 5.235 ;
        RECT 41.390 4.855 41.690 5.405 ;
        RECT 44.170 5.315 45.050 5.355 ;
        RECT 43.520 5.115 45.050 5.315 ;
        RECT 43.520 4.985 43.690 5.115 ;
        RECT 44.435 5.065 45.050 5.115 ;
        RECT 44.820 5.025 45.050 5.065 ;
        RECT 45.220 5.025 45.550 5.525 ;
        RECT 44.380 4.855 44.710 4.895 ;
        RECT 45.220 4.855 46.040 5.025 ;
        RECT 48.260 5.015 48.430 6.475 ;
        RECT 48.835 6.245 49.005 7.855 ;
        RECT 49.210 7.795 49.380 8.305 ;
        RECT 48.780 6.075 49.005 6.245 ;
        RECT 48.780 5.015 48.950 6.075 ;
        RECT 49.210 5.015 49.380 7.225 ;
        RECT 49.640 5.015 49.810 8.305 ;
        RECT 51.005 7.795 51.175 8.305 ;
        RECT 51.995 7.795 52.165 8.305 ;
        RECT 53.620 7.645 53.790 8.305 ;
        RECT 54.570 7.795 54.740 8.305 ;
        RECT 53.620 7.315 54.025 7.645 ;
        RECT 50.635 6.970 51.100 7.140 ;
        RECT 51.625 6.970 52.090 7.140 ;
        RECT 50.635 5.945 50.805 6.970 ;
        RECT 51.005 5.015 51.175 6.485 ;
        RECT 51.625 5.945 51.795 6.970 ;
        RECT 53.620 6.805 53.790 7.315 ;
        RECT 51.995 5.015 52.165 6.485 ;
        RECT 53.620 6.475 54.025 6.805 ;
        RECT 53.620 5.015 53.790 6.475 ;
        RECT 54.570 5.015 54.740 7.225 ;
        RECT 55.000 5.015 55.170 8.305 ;
        RECT 64.845 7.645 65.015 8.305 ;
        RECT 65.365 8.025 65.535 8.305 ;
        RECT 65.365 7.855 65.590 8.025 ;
        RECT 64.845 7.315 65.250 7.645 ;
        RECT 56.795 6.605 57.355 6.895 ;
        RECT 56.795 5.235 57.045 6.605 ;
        RECT 58.395 6.435 58.725 6.795 ;
        RECT 60.105 6.645 61.410 6.895 ;
        RECT 64.845 6.805 65.015 7.315 ;
        RECT 60.105 6.495 60.285 6.645 ;
        RECT 57.335 6.245 58.725 6.435 ;
        RECT 59.555 6.325 60.285 6.495 ;
        RECT 64.845 6.475 65.250 6.805 ;
        RECT 57.335 6.155 57.505 6.245 ;
        RECT 57.215 5.825 57.505 6.155 ;
        RECT 58.235 5.825 58.910 6.075 ;
        RECT 57.335 5.575 57.505 5.825 ;
        RECT 57.335 5.405 58.275 5.575 ;
        RECT 58.645 5.465 58.910 5.825 ;
        RECT 59.555 5.655 59.725 6.325 ;
        RECT 60.530 6.075 60.740 6.475 ;
        RECT 60.390 5.875 60.740 6.075 ;
        RECT 60.990 6.075 61.240 6.475 ;
        RECT 60.990 5.875 61.465 6.075 ;
        RECT 61.655 5.875 62.105 6.385 ;
        RECT 60.390 5.655 62.135 5.705 ;
        RECT 59.555 5.525 62.135 5.655 ;
        RECT 59.555 5.485 60.615 5.525 ;
        RECT 44.380 4.685 45.550 4.855 ;
        RECT 56.795 4.685 57.255 5.235 ;
        RECT 57.975 4.855 58.275 5.405 ;
        RECT 60.755 5.315 61.635 5.355 ;
        RECT 60.105 5.115 61.635 5.315 ;
        RECT 60.105 4.985 60.275 5.115 ;
        RECT 61.020 5.065 61.635 5.115 ;
        RECT 61.405 5.025 61.635 5.065 ;
        RECT 61.805 5.025 62.135 5.525 ;
        RECT 60.965 4.855 61.295 4.895 ;
        RECT 61.805 4.855 62.625 5.025 ;
        RECT 64.845 5.015 65.015 6.475 ;
        RECT 65.420 6.245 65.590 7.855 ;
        RECT 65.795 7.795 65.965 8.305 ;
        RECT 65.365 6.075 65.590 6.245 ;
        RECT 65.365 5.015 65.535 6.075 ;
        RECT 65.795 5.015 65.965 7.225 ;
        RECT 66.225 5.015 66.395 8.305 ;
        RECT 67.590 7.795 67.760 8.305 ;
        RECT 68.580 7.795 68.750 8.305 ;
        RECT 70.200 7.645 70.370 8.305 ;
        RECT 71.150 7.795 71.320 8.305 ;
        RECT 70.200 7.315 70.605 7.645 ;
        RECT 67.220 6.970 67.685 7.140 ;
        RECT 68.210 6.970 68.675 7.140 ;
        RECT 67.220 5.945 67.390 6.970 ;
        RECT 67.590 5.015 67.760 6.485 ;
        RECT 68.210 5.945 68.380 6.970 ;
        RECT 70.200 6.805 70.370 7.315 ;
        RECT 68.580 5.015 68.750 6.485 ;
        RECT 70.200 6.475 70.605 6.805 ;
        RECT 70.200 5.015 70.370 6.475 ;
        RECT 71.150 5.015 71.320 7.225 ;
        RECT 71.580 5.015 71.750 8.305 ;
        RECT 81.425 7.645 81.595 8.305 ;
        RECT 81.945 8.025 82.115 8.305 ;
        RECT 81.945 7.855 82.170 8.025 ;
        RECT 81.425 7.315 81.830 7.645 ;
        RECT 73.375 6.605 73.935 6.895 ;
        RECT 73.375 5.235 73.625 6.605 ;
        RECT 74.975 6.435 75.305 6.795 ;
        RECT 76.685 6.645 77.990 6.895 ;
        RECT 81.425 6.805 81.595 7.315 ;
        RECT 76.685 6.495 76.865 6.645 ;
        RECT 73.915 6.245 75.305 6.435 ;
        RECT 76.135 6.325 76.865 6.495 ;
        RECT 81.425 6.475 81.830 6.805 ;
        RECT 73.915 6.155 74.085 6.245 ;
        RECT 73.795 5.825 74.085 6.155 ;
        RECT 74.815 5.825 75.490 6.075 ;
        RECT 73.915 5.575 74.085 5.825 ;
        RECT 73.915 5.405 74.855 5.575 ;
        RECT 75.225 5.465 75.490 5.825 ;
        RECT 76.135 5.655 76.305 6.325 ;
        RECT 77.110 6.075 77.320 6.475 ;
        RECT 76.970 5.875 77.320 6.075 ;
        RECT 77.570 6.075 77.820 6.475 ;
        RECT 77.570 5.875 78.045 6.075 ;
        RECT 78.235 5.875 78.685 6.385 ;
        RECT 76.970 5.655 78.715 5.705 ;
        RECT 76.135 5.525 78.715 5.655 ;
        RECT 76.135 5.485 77.195 5.525 ;
        RECT 60.965 4.685 62.135 4.855 ;
        RECT 73.375 4.685 73.835 5.235 ;
        RECT 74.555 4.855 74.855 5.405 ;
        RECT 77.335 5.315 78.215 5.355 ;
        RECT 76.685 5.115 78.215 5.315 ;
        RECT 76.685 4.985 76.855 5.115 ;
        RECT 77.600 5.065 78.215 5.115 ;
        RECT 77.985 5.025 78.215 5.065 ;
        RECT 78.385 5.025 78.715 5.525 ;
        RECT 77.545 4.855 77.875 4.895 ;
        RECT 78.385 4.855 79.205 5.025 ;
        RECT 81.425 5.015 81.595 6.475 ;
        RECT 82.000 6.245 82.170 7.855 ;
        RECT 82.375 7.795 82.545 8.305 ;
        RECT 81.945 6.075 82.170 6.245 ;
        RECT 81.945 5.015 82.115 6.075 ;
        RECT 82.375 5.015 82.545 7.225 ;
        RECT 82.805 5.015 82.975 8.305 ;
        RECT 84.170 7.795 84.340 8.305 ;
        RECT 85.160 7.795 85.330 8.305 ;
        RECT 83.800 6.970 84.265 7.140 ;
        RECT 84.790 6.970 85.255 7.140 ;
        RECT 83.800 5.945 83.970 6.970 ;
        RECT 84.170 5.015 84.340 6.485 ;
        RECT 84.790 5.945 84.960 6.970 ;
        RECT 85.160 5.015 85.330 6.485 ;
        RECT 77.545 4.685 78.715 4.855 ;
        RECT 6.580 2.785 6.920 3.665 ;
        RECT 7.090 2.955 7.260 4.175 ;
        RECT 8.285 3.835 8.760 4.175 ;
        RECT 7.500 3.305 7.750 3.670 ;
        RECT 8.470 3.305 9.185 3.600 ;
        RECT 9.355 3.475 9.630 4.175 ;
        RECT 10.580 3.835 11.060 4.175 ;
        RECT 7.500 3.135 9.290 3.305 ;
        RECT 7.090 2.705 7.885 2.955 ;
        RECT 7.090 2.615 7.340 2.705 ;
        RECT 7.010 2.195 7.340 2.615 ;
        RECT 8.055 2.280 8.310 3.135 ;
        RECT 7.520 2.015 8.310 2.280 ;
        RECT 8.480 2.435 8.890 2.955 ;
        RECT 9.060 2.770 9.290 3.135 ;
        RECT 9.460 2.770 9.630 3.475 ;
        RECT 9.800 3.070 10.060 3.520 ;
        RECT 10.730 3.345 11.485 3.595 ;
        RECT 11.655 3.475 11.930 4.175 ;
        RECT 10.715 3.310 11.485 3.345 ;
        RECT 10.700 3.300 11.485 3.310 ;
        RECT 10.695 3.285 11.590 3.300 ;
        RECT 10.675 3.270 11.590 3.285 ;
        RECT 10.655 3.260 11.590 3.270 ;
        RECT 10.630 3.250 11.590 3.260 ;
        RECT 10.560 3.220 11.590 3.250 ;
        RECT 10.540 3.190 11.590 3.220 ;
        RECT 10.520 3.160 11.590 3.190 ;
        RECT 10.490 3.135 11.590 3.160 ;
        RECT 10.455 3.100 11.590 3.135 ;
        RECT 10.425 3.095 11.590 3.100 ;
        RECT 10.425 3.090 10.815 3.095 ;
        RECT 10.425 3.080 10.790 3.090 ;
        RECT 10.425 3.075 10.775 3.080 ;
        RECT 10.425 3.070 10.760 3.075 ;
        RECT 9.800 3.065 10.760 3.070 ;
        RECT 9.800 3.055 10.750 3.065 ;
        RECT 9.800 3.050 10.740 3.055 ;
        RECT 9.800 3.040 10.730 3.050 ;
        RECT 9.800 3.030 10.725 3.040 ;
        RECT 9.800 3.025 10.720 3.030 ;
        RECT 9.800 3.010 10.710 3.025 ;
        RECT 9.800 2.995 10.705 3.010 ;
        RECT 9.800 2.970 10.695 2.995 ;
        RECT 9.800 2.900 10.690 2.970 ;
        RECT 9.060 2.765 9.120 2.770 ;
        RECT 9.575 2.765 9.630 2.770 ;
        RECT 9.060 2.705 9.290 2.765 ;
        RECT 9.120 2.700 9.290 2.705 ;
        RECT 9.460 2.440 9.630 2.765 ;
        RECT 8.480 2.015 8.680 2.435 ;
        RECT 9.370 1.965 9.630 2.440 ;
        RECT 9.800 2.345 10.350 2.730 ;
        RECT 10.520 2.175 10.690 2.900 ;
        RECT 9.800 2.005 10.690 2.175 ;
        RECT 10.860 2.500 11.190 2.925 ;
        RECT 11.360 2.700 11.590 3.095 ;
        RECT 11.760 2.985 11.930 3.475 ;
        RECT 12.110 3.375 12.440 4.160 ;
        RECT 12.110 3.205 12.790 3.375 ;
        RECT 12.100 2.985 12.450 3.035 ;
        RECT 11.760 2.815 12.450 2.985 ;
        RECT 10.860 2.015 11.080 2.500 ;
        RECT 11.760 2.445 11.930 2.815 ;
        RECT 12.100 2.785 12.450 2.815 ;
        RECT 12.620 2.605 12.790 3.205 ;
        RECT 12.960 2.785 13.310 3.035 ;
        RECT 11.670 1.965 11.930 2.445 ;
        RECT 12.530 1.965 12.860 2.605 ;
        RECT 15.090 2.405 15.260 3.865 ;
        RECT 15.610 2.805 15.780 3.865 ;
        RECT 15.610 2.635 15.835 2.805 ;
        RECT 15.090 2.075 15.495 2.405 ;
        RECT 15.090 1.565 15.260 2.075 ;
        RECT 15.090 1.235 15.495 1.565 ;
        RECT 15.090 0.575 15.260 1.235 ;
        RECT 15.665 1.025 15.835 2.635 ;
        RECT 16.040 1.655 16.210 3.865 ;
        RECT 15.610 0.855 15.835 1.025 ;
        RECT 15.610 0.575 15.780 0.855 ;
        RECT 16.040 0.575 16.210 1.085 ;
        RECT 16.470 0.575 16.640 3.865 ;
        RECT 17.465 1.910 17.635 2.935 ;
        RECT 17.835 2.395 18.005 3.865 ;
        RECT 18.455 1.910 18.625 2.935 ;
        RECT 23.165 2.785 23.505 3.665 ;
        RECT 23.675 2.955 23.845 4.175 ;
        RECT 24.870 3.835 25.345 4.175 ;
        RECT 24.085 3.305 24.335 3.670 ;
        RECT 25.055 3.305 25.770 3.600 ;
        RECT 25.940 3.475 26.215 4.175 ;
        RECT 27.165 3.835 27.645 4.175 ;
        RECT 24.085 3.135 25.875 3.305 ;
        RECT 23.675 2.705 24.470 2.955 ;
        RECT 23.675 2.615 23.925 2.705 ;
        RECT 23.595 2.195 23.925 2.615 ;
        RECT 24.640 2.280 24.895 3.135 ;
        RECT 24.105 2.015 24.895 2.280 ;
        RECT 25.065 2.435 25.475 2.955 ;
        RECT 25.645 2.770 25.875 3.135 ;
        RECT 26.045 2.770 26.215 3.475 ;
        RECT 26.385 3.070 26.645 3.520 ;
        RECT 27.315 3.345 28.070 3.595 ;
        RECT 28.240 3.475 28.515 4.175 ;
        RECT 27.300 3.310 28.070 3.345 ;
        RECT 27.285 3.300 28.070 3.310 ;
        RECT 27.280 3.285 28.175 3.300 ;
        RECT 27.260 3.270 28.175 3.285 ;
        RECT 27.240 3.260 28.175 3.270 ;
        RECT 27.215 3.250 28.175 3.260 ;
        RECT 27.145 3.220 28.175 3.250 ;
        RECT 27.125 3.190 28.175 3.220 ;
        RECT 27.105 3.160 28.175 3.190 ;
        RECT 27.075 3.135 28.175 3.160 ;
        RECT 27.040 3.100 28.175 3.135 ;
        RECT 27.010 3.095 28.175 3.100 ;
        RECT 27.010 3.090 27.400 3.095 ;
        RECT 27.010 3.080 27.375 3.090 ;
        RECT 27.010 3.075 27.360 3.080 ;
        RECT 27.010 3.070 27.345 3.075 ;
        RECT 26.385 3.065 27.345 3.070 ;
        RECT 26.385 3.055 27.335 3.065 ;
        RECT 26.385 3.050 27.325 3.055 ;
        RECT 26.385 3.040 27.315 3.050 ;
        RECT 26.385 3.030 27.310 3.040 ;
        RECT 26.385 3.025 27.305 3.030 ;
        RECT 26.385 3.010 27.295 3.025 ;
        RECT 26.385 2.995 27.290 3.010 ;
        RECT 26.385 2.970 27.280 2.995 ;
        RECT 26.385 2.900 27.275 2.970 ;
        RECT 25.645 2.765 25.705 2.770 ;
        RECT 26.160 2.765 26.215 2.770 ;
        RECT 25.645 2.705 25.875 2.765 ;
        RECT 25.705 2.700 25.875 2.705 ;
        RECT 26.045 2.440 26.215 2.765 ;
        RECT 25.065 2.015 25.265 2.435 ;
        RECT 25.955 1.965 26.215 2.440 ;
        RECT 26.385 2.345 26.935 2.730 ;
        RECT 27.105 2.175 27.275 2.900 ;
        RECT 26.385 2.005 27.275 2.175 ;
        RECT 27.445 2.500 27.775 2.925 ;
        RECT 27.945 2.700 28.175 3.095 ;
        RECT 28.345 2.985 28.515 3.475 ;
        RECT 28.695 3.375 29.025 4.160 ;
        RECT 28.695 3.205 29.375 3.375 ;
        RECT 28.685 2.985 29.035 3.035 ;
        RECT 28.345 2.815 29.035 2.985 ;
        RECT 27.445 2.015 27.665 2.500 ;
        RECT 28.345 2.445 28.515 2.815 ;
        RECT 28.685 2.785 29.035 2.815 ;
        RECT 29.205 2.605 29.375 3.205 ;
        RECT 29.545 2.785 29.895 3.035 ;
        RECT 28.255 1.965 28.515 2.445 ;
        RECT 29.115 1.965 29.445 2.605 ;
        RECT 31.675 2.405 31.845 3.865 ;
        RECT 32.195 2.805 32.365 3.865 ;
        RECT 32.195 2.635 32.420 2.805 ;
        RECT 31.675 2.075 32.080 2.405 ;
        RECT 17.465 1.740 17.930 1.910 ;
        RECT 18.455 1.740 18.920 1.910 ;
        RECT 31.675 1.565 31.845 2.075 ;
        RECT 31.675 1.235 32.080 1.565 ;
        RECT 17.835 0.575 18.005 1.085 ;
        RECT 31.675 0.575 31.845 1.235 ;
        RECT 32.250 1.025 32.420 2.635 ;
        RECT 32.625 1.655 32.795 3.865 ;
        RECT 32.195 0.855 32.420 1.025 ;
        RECT 32.195 0.575 32.365 0.855 ;
        RECT 32.625 0.575 32.795 1.085 ;
        RECT 33.055 0.575 33.225 3.865 ;
        RECT 34.050 1.910 34.220 2.935 ;
        RECT 34.420 2.395 34.590 3.865 ;
        RECT 35.040 1.910 35.210 2.935 ;
        RECT 39.750 2.785 40.090 3.665 ;
        RECT 40.260 2.955 40.430 4.175 ;
        RECT 41.455 3.835 41.930 4.175 ;
        RECT 40.670 3.305 40.920 3.670 ;
        RECT 41.640 3.305 42.355 3.600 ;
        RECT 42.525 3.475 42.800 4.175 ;
        RECT 43.750 3.835 44.230 4.175 ;
        RECT 40.670 3.135 42.460 3.305 ;
        RECT 40.260 2.705 41.055 2.955 ;
        RECT 40.260 2.615 40.510 2.705 ;
        RECT 40.180 2.195 40.510 2.615 ;
        RECT 41.225 2.280 41.480 3.135 ;
        RECT 40.690 2.015 41.480 2.280 ;
        RECT 41.650 2.435 42.060 2.955 ;
        RECT 42.230 2.770 42.460 3.135 ;
        RECT 42.630 2.770 42.800 3.475 ;
        RECT 42.970 3.070 43.230 3.520 ;
        RECT 43.900 3.345 44.655 3.595 ;
        RECT 44.825 3.475 45.100 4.175 ;
        RECT 43.885 3.310 44.655 3.345 ;
        RECT 43.870 3.300 44.655 3.310 ;
        RECT 43.865 3.285 44.760 3.300 ;
        RECT 43.845 3.270 44.760 3.285 ;
        RECT 43.825 3.260 44.760 3.270 ;
        RECT 43.800 3.250 44.760 3.260 ;
        RECT 43.730 3.220 44.760 3.250 ;
        RECT 43.710 3.190 44.760 3.220 ;
        RECT 43.690 3.160 44.760 3.190 ;
        RECT 43.660 3.135 44.760 3.160 ;
        RECT 43.625 3.100 44.760 3.135 ;
        RECT 43.595 3.095 44.760 3.100 ;
        RECT 43.595 3.090 43.985 3.095 ;
        RECT 43.595 3.080 43.960 3.090 ;
        RECT 43.595 3.075 43.945 3.080 ;
        RECT 43.595 3.070 43.930 3.075 ;
        RECT 42.970 3.065 43.930 3.070 ;
        RECT 42.970 3.055 43.920 3.065 ;
        RECT 42.970 3.050 43.910 3.055 ;
        RECT 42.970 3.040 43.900 3.050 ;
        RECT 42.970 3.030 43.895 3.040 ;
        RECT 42.970 3.025 43.890 3.030 ;
        RECT 42.970 3.010 43.880 3.025 ;
        RECT 42.970 2.995 43.875 3.010 ;
        RECT 42.970 2.970 43.865 2.995 ;
        RECT 42.970 2.900 43.860 2.970 ;
        RECT 42.230 2.765 42.290 2.770 ;
        RECT 42.745 2.765 42.800 2.770 ;
        RECT 42.230 2.705 42.460 2.765 ;
        RECT 42.290 2.700 42.460 2.705 ;
        RECT 42.630 2.440 42.800 2.765 ;
        RECT 41.650 2.015 41.850 2.435 ;
        RECT 42.540 1.965 42.800 2.440 ;
        RECT 42.970 2.345 43.520 2.730 ;
        RECT 43.690 2.175 43.860 2.900 ;
        RECT 42.970 2.005 43.860 2.175 ;
        RECT 44.030 2.500 44.360 2.925 ;
        RECT 44.530 2.700 44.760 3.095 ;
        RECT 44.930 2.985 45.100 3.475 ;
        RECT 45.280 3.375 45.610 4.160 ;
        RECT 45.280 3.205 45.960 3.375 ;
        RECT 45.270 2.985 45.620 3.035 ;
        RECT 44.930 2.815 45.620 2.985 ;
        RECT 44.030 2.015 44.250 2.500 ;
        RECT 44.930 2.445 45.100 2.815 ;
        RECT 45.270 2.785 45.620 2.815 ;
        RECT 45.790 2.605 45.960 3.205 ;
        RECT 46.130 2.785 46.480 3.035 ;
        RECT 44.840 1.965 45.100 2.445 ;
        RECT 45.700 1.965 46.030 2.605 ;
        RECT 48.260 2.405 48.430 3.865 ;
        RECT 48.780 2.805 48.950 3.865 ;
        RECT 48.780 2.635 49.005 2.805 ;
        RECT 48.260 2.075 48.665 2.405 ;
        RECT 34.050 1.740 34.515 1.910 ;
        RECT 35.040 1.740 35.505 1.910 ;
        RECT 48.260 1.565 48.430 2.075 ;
        RECT 48.260 1.235 48.665 1.565 ;
        RECT 34.420 0.575 34.590 1.085 ;
        RECT 48.260 0.575 48.430 1.235 ;
        RECT 48.835 1.025 49.005 2.635 ;
        RECT 49.210 1.655 49.380 3.865 ;
        RECT 48.780 0.855 49.005 1.025 ;
        RECT 48.780 0.575 48.950 0.855 ;
        RECT 49.210 0.575 49.380 1.085 ;
        RECT 49.640 0.575 49.810 3.865 ;
        RECT 50.635 1.910 50.805 2.935 ;
        RECT 51.005 2.395 51.175 3.865 ;
        RECT 51.625 1.910 51.795 2.935 ;
        RECT 56.335 2.785 56.675 3.665 ;
        RECT 56.845 2.955 57.015 4.175 ;
        RECT 58.040 3.835 58.515 4.175 ;
        RECT 57.255 3.305 57.505 3.670 ;
        RECT 58.225 3.305 58.940 3.600 ;
        RECT 59.110 3.475 59.385 4.175 ;
        RECT 60.335 3.835 60.815 4.175 ;
        RECT 57.255 3.135 59.045 3.305 ;
        RECT 56.845 2.705 57.640 2.955 ;
        RECT 56.845 2.615 57.095 2.705 ;
        RECT 56.765 2.195 57.095 2.615 ;
        RECT 57.810 2.280 58.065 3.135 ;
        RECT 57.275 2.015 58.065 2.280 ;
        RECT 58.235 2.435 58.645 2.955 ;
        RECT 58.815 2.770 59.045 3.135 ;
        RECT 59.215 2.770 59.385 3.475 ;
        RECT 59.555 3.070 59.815 3.520 ;
        RECT 60.485 3.345 61.240 3.595 ;
        RECT 61.410 3.475 61.685 4.175 ;
        RECT 60.470 3.310 61.240 3.345 ;
        RECT 60.455 3.300 61.240 3.310 ;
        RECT 60.450 3.285 61.345 3.300 ;
        RECT 60.430 3.270 61.345 3.285 ;
        RECT 60.410 3.260 61.345 3.270 ;
        RECT 60.385 3.250 61.345 3.260 ;
        RECT 60.315 3.220 61.345 3.250 ;
        RECT 60.295 3.190 61.345 3.220 ;
        RECT 60.275 3.160 61.345 3.190 ;
        RECT 60.245 3.135 61.345 3.160 ;
        RECT 60.210 3.100 61.345 3.135 ;
        RECT 60.180 3.095 61.345 3.100 ;
        RECT 60.180 3.090 60.570 3.095 ;
        RECT 60.180 3.080 60.545 3.090 ;
        RECT 60.180 3.075 60.530 3.080 ;
        RECT 60.180 3.070 60.515 3.075 ;
        RECT 59.555 3.065 60.515 3.070 ;
        RECT 59.555 3.055 60.505 3.065 ;
        RECT 59.555 3.050 60.495 3.055 ;
        RECT 59.555 3.040 60.485 3.050 ;
        RECT 59.555 3.030 60.480 3.040 ;
        RECT 59.555 3.025 60.475 3.030 ;
        RECT 59.555 3.010 60.465 3.025 ;
        RECT 59.555 2.995 60.460 3.010 ;
        RECT 59.555 2.970 60.450 2.995 ;
        RECT 59.555 2.900 60.445 2.970 ;
        RECT 58.815 2.765 58.875 2.770 ;
        RECT 59.330 2.765 59.385 2.770 ;
        RECT 58.815 2.705 59.045 2.765 ;
        RECT 58.875 2.700 59.045 2.705 ;
        RECT 59.215 2.440 59.385 2.765 ;
        RECT 58.235 2.015 58.435 2.435 ;
        RECT 59.125 1.965 59.385 2.440 ;
        RECT 59.555 2.345 60.105 2.730 ;
        RECT 60.275 2.175 60.445 2.900 ;
        RECT 59.555 2.005 60.445 2.175 ;
        RECT 60.615 2.500 60.945 2.925 ;
        RECT 61.115 2.700 61.345 3.095 ;
        RECT 61.515 2.985 61.685 3.475 ;
        RECT 61.865 3.375 62.195 4.160 ;
        RECT 61.865 3.205 62.545 3.375 ;
        RECT 61.855 2.985 62.205 3.035 ;
        RECT 61.515 2.815 62.205 2.985 ;
        RECT 60.615 2.015 60.835 2.500 ;
        RECT 61.515 2.445 61.685 2.815 ;
        RECT 61.855 2.785 62.205 2.815 ;
        RECT 62.375 2.605 62.545 3.205 ;
        RECT 62.715 2.785 63.065 3.035 ;
        RECT 61.425 1.965 61.685 2.445 ;
        RECT 62.285 1.965 62.615 2.605 ;
        RECT 64.845 2.405 65.015 3.865 ;
        RECT 65.365 2.805 65.535 3.865 ;
        RECT 65.365 2.635 65.590 2.805 ;
        RECT 64.845 2.075 65.250 2.405 ;
        RECT 50.635 1.740 51.100 1.910 ;
        RECT 51.625 1.740 52.090 1.910 ;
        RECT 64.845 1.565 65.015 2.075 ;
        RECT 64.845 1.235 65.250 1.565 ;
        RECT 51.005 0.575 51.175 1.085 ;
        RECT 64.845 0.575 65.015 1.235 ;
        RECT 65.420 1.025 65.590 2.635 ;
        RECT 65.795 1.655 65.965 3.865 ;
        RECT 65.365 0.855 65.590 1.025 ;
        RECT 65.365 0.575 65.535 0.855 ;
        RECT 65.795 0.575 65.965 1.085 ;
        RECT 66.225 0.575 66.395 3.865 ;
        RECT 67.220 1.910 67.390 2.935 ;
        RECT 67.590 2.395 67.760 3.865 ;
        RECT 68.210 1.910 68.380 2.935 ;
        RECT 72.915 2.785 73.255 3.665 ;
        RECT 73.425 2.955 73.595 4.175 ;
        RECT 74.620 3.835 75.095 4.175 ;
        RECT 73.835 3.305 74.085 3.670 ;
        RECT 74.805 3.305 75.520 3.600 ;
        RECT 75.690 3.475 75.965 4.175 ;
        RECT 76.915 3.835 77.395 4.175 ;
        RECT 73.835 3.135 75.625 3.305 ;
        RECT 73.425 2.705 74.220 2.955 ;
        RECT 73.425 2.615 73.675 2.705 ;
        RECT 73.345 2.195 73.675 2.615 ;
        RECT 74.390 2.280 74.645 3.135 ;
        RECT 73.855 2.015 74.645 2.280 ;
        RECT 74.815 2.435 75.225 2.955 ;
        RECT 75.395 2.770 75.625 3.135 ;
        RECT 75.795 2.770 75.965 3.475 ;
        RECT 76.135 3.070 76.395 3.520 ;
        RECT 77.065 3.345 77.820 3.595 ;
        RECT 77.990 3.475 78.265 4.175 ;
        RECT 77.050 3.310 77.820 3.345 ;
        RECT 77.035 3.300 77.820 3.310 ;
        RECT 77.030 3.285 77.925 3.300 ;
        RECT 77.010 3.270 77.925 3.285 ;
        RECT 76.990 3.260 77.925 3.270 ;
        RECT 76.965 3.250 77.925 3.260 ;
        RECT 76.895 3.220 77.925 3.250 ;
        RECT 76.875 3.190 77.925 3.220 ;
        RECT 76.855 3.160 77.925 3.190 ;
        RECT 76.825 3.135 77.925 3.160 ;
        RECT 76.790 3.100 77.925 3.135 ;
        RECT 76.760 3.095 77.925 3.100 ;
        RECT 76.760 3.090 77.150 3.095 ;
        RECT 76.760 3.080 77.125 3.090 ;
        RECT 76.760 3.075 77.110 3.080 ;
        RECT 76.760 3.070 77.095 3.075 ;
        RECT 76.135 3.065 77.095 3.070 ;
        RECT 76.135 3.055 77.085 3.065 ;
        RECT 76.135 3.050 77.075 3.055 ;
        RECT 76.135 3.040 77.065 3.050 ;
        RECT 76.135 3.030 77.060 3.040 ;
        RECT 76.135 3.025 77.055 3.030 ;
        RECT 76.135 3.010 77.045 3.025 ;
        RECT 76.135 2.995 77.040 3.010 ;
        RECT 76.135 2.970 77.030 2.995 ;
        RECT 76.135 2.900 77.025 2.970 ;
        RECT 75.395 2.765 75.455 2.770 ;
        RECT 75.910 2.765 75.965 2.770 ;
        RECT 75.395 2.705 75.625 2.765 ;
        RECT 75.455 2.700 75.625 2.705 ;
        RECT 75.795 2.440 75.965 2.765 ;
        RECT 74.815 2.015 75.015 2.435 ;
        RECT 75.705 1.965 75.965 2.440 ;
        RECT 76.135 2.345 76.685 2.730 ;
        RECT 76.855 2.175 77.025 2.900 ;
        RECT 76.135 2.005 77.025 2.175 ;
        RECT 77.195 2.500 77.525 2.925 ;
        RECT 77.695 2.700 77.925 3.095 ;
        RECT 78.095 2.985 78.265 3.475 ;
        RECT 78.445 3.375 78.775 4.160 ;
        RECT 78.445 3.205 79.125 3.375 ;
        RECT 78.435 2.985 78.785 3.035 ;
        RECT 78.095 2.815 78.785 2.985 ;
        RECT 77.195 2.015 77.415 2.500 ;
        RECT 78.095 2.445 78.265 2.815 ;
        RECT 78.435 2.785 78.785 2.815 ;
        RECT 78.955 2.605 79.125 3.205 ;
        RECT 79.295 2.785 79.645 3.035 ;
        RECT 78.005 1.965 78.265 2.445 ;
        RECT 78.865 1.965 79.195 2.605 ;
        RECT 81.425 2.405 81.595 3.865 ;
        RECT 81.945 2.805 82.115 3.865 ;
        RECT 81.945 2.635 82.170 2.805 ;
        RECT 81.425 2.075 81.830 2.405 ;
        RECT 67.220 1.740 67.685 1.910 ;
        RECT 68.210 1.740 68.675 1.910 ;
        RECT 81.425 1.565 81.595 2.075 ;
        RECT 81.425 1.235 81.830 1.565 ;
        RECT 67.590 0.575 67.760 1.085 ;
        RECT 81.425 0.575 81.595 1.235 ;
        RECT 82.000 1.025 82.170 2.635 ;
        RECT 82.375 1.655 82.545 3.865 ;
        RECT 81.945 0.855 82.170 1.025 ;
        RECT 81.945 0.575 82.115 0.855 ;
        RECT 82.375 0.575 82.545 1.085 ;
        RECT 82.805 0.575 82.975 3.865 ;
        RECT 83.800 1.910 83.970 2.935 ;
        RECT 84.170 2.395 84.340 3.865 ;
        RECT 84.790 1.910 84.960 2.935 ;
        RECT 83.800 1.740 84.265 1.910 ;
        RECT 84.790 1.740 85.255 1.910 ;
        RECT 84.170 0.575 84.340 1.085 ;
      LAYER mcon ;
        RECT 1.210 6.315 1.380 6.485 ;
        RECT 1.585 7.055 1.755 7.225 ;
        RECT 4.815 7.055 4.985 7.225 ;
        RECT 5.245 6.685 5.415 6.855 ;
        RECT 8.960 5.875 9.130 6.045 ;
        RECT 10.660 5.875 10.830 6.045 ;
        RECT 11.340 5.875 11.510 6.045 ;
        RECT 12.020 5.875 12.190 6.045 ;
        RECT 7.260 4.855 7.430 5.025 ;
        RECT 12.700 4.855 12.870 5.025 ;
        RECT 15.665 6.315 15.835 6.485 ;
        RECT 16.040 7.055 16.210 7.225 ;
        RECT 16.470 6.685 16.640 6.855 ;
        RECT 17.835 6.315 18.005 6.485 ;
        RECT 21.400 7.055 21.570 7.225 ;
        RECT 18.825 6.315 18.995 6.485 ;
        RECT 21.830 6.685 22.000 6.855 ;
        RECT 25.545 5.875 25.715 6.045 ;
        RECT 27.245 5.875 27.415 6.045 ;
        RECT 27.925 5.875 28.095 6.045 ;
        RECT 28.605 5.875 28.775 6.045 ;
        RECT 23.845 4.855 24.015 5.025 ;
        RECT 29.285 4.855 29.455 5.025 ;
        RECT 32.250 6.315 32.420 6.485 ;
        RECT 32.625 7.055 32.795 7.225 ;
        RECT 33.055 6.685 33.225 6.855 ;
        RECT 34.420 6.315 34.590 6.485 ;
        RECT 37.985 7.055 38.155 7.225 ;
        RECT 35.410 6.315 35.580 6.485 ;
        RECT 38.415 6.685 38.585 6.855 ;
        RECT 42.130 5.875 42.300 6.045 ;
        RECT 43.830 5.875 44.000 6.045 ;
        RECT 44.510 5.875 44.680 6.045 ;
        RECT 45.190 5.875 45.360 6.045 ;
        RECT 40.430 4.855 40.600 5.025 ;
        RECT 45.870 4.855 46.040 5.025 ;
        RECT 48.835 6.315 49.005 6.485 ;
        RECT 49.210 7.055 49.380 7.225 ;
        RECT 49.640 6.685 49.810 6.855 ;
        RECT 51.005 6.315 51.175 6.485 ;
        RECT 54.570 7.055 54.740 7.225 ;
        RECT 51.995 6.315 52.165 6.485 ;
        RECT 55.000 6.685 55.170 6.855 ;
        RECT 58.715 5.875 58.885 6.045 ;
        RECT 60.415 5.875 60.585 6.045 ;
        RECT 61.095 5.875 61.265 6.045 ;
        RECT 61.775 5.875 61.945 6.045 ;
        RECT 57.015 4.855 57.185 5.025 ;
        RECT 62.455 4.855 62.625 5.025 ;
        RECT 65.420 6.315 65.590 6.485 ;
        RECT 65.795 7.055 65.965 7.225 ;
        RECT 66.225 6.685 66.395 6.855 ;
        RECT 67.590 6.315 67.760 6.485 ;
        RECT 71.150 7.055 71.320 7.225 ;
        RECT 68.580 6.315 68.750 6.485 ;
        RECT 71.580 6.685 71.750 6.855 ;
        RECT 75.295 5.875 75.465 6.045 ;
        RECT 76.995 5.875 77.165 6.045 ;
        RECT 77.675 5.875 77.845 6.045 ;
        RECT 78.355 5.875 78.525 6.045 ;
        RECT 73.595 4.855 73.765 5.025 ;
        RECT 79.035 4.855 79.205 5.025 ;
        RECT 82.000 6.315 82.170 6.485 ;
        RECT 82.375 7.055 82.545 7.225 ;
        RECT 82.805 6.685 82.975 6.855 ;
        RECT 84.170 6.315 84.340 6.485 ;
        RECT 85.160 6.315 85.330 6.485 ;
        RECT 6.585 2.815 6.755 2.985 ;
        RECT 8.450 3.835 8.620 4.005 ;
        RECT 10.660 3.835 10.830 4.005 ;
        RECT 8.620 2.475 8.790 2.645 ;
        RECT 9.575 2.640 9.630 2.645 ;
        RECT 9.460 2.475 9.630 2.640 ;
        RECT 9.460 2.470 9.575 2.475 ;
        RECT 9.980 2.475 10.150 2.645 ;
        RECT 12.620 3.155 12.790 3.325 ;
        RECT 13.040 2.815 13.210 2.985 ;
        RECT 10.885 2.135 11.055 2.305 ;
        RECT 11.680 2.135 11.850 2.305 ;
        RECT 15.665 2.395 15.835 2.565 ;
        RECT 16.470 2.025 16.640 2.195 ;
        RECT 16.040 0.915 16.210 1.085 ;
        RECT 17.465 2.765 17.635 2.935 ;
        RECT 18.455 2.765 18.625 2.935 ;
        RECT 23.170 2.815 23.340 2.985 ;
        RECT 25.035 3.835 25.205 4.005 ;
        RECT 27.245 3.835 27.415 4.005 ;
        RECT 25.205 2.475 25.375 2.645 ;
        RECT 26.160 2.640 26.215 2.645 ;
        RECT 26.045 2.475 26.215 2.640 ;
        RECT 26.045 2.470 26.160 2.475 ;
        RECT 26.565 2.475 26.735 2.645 ;
        RECT 29.205 3.155 29.375 3.325 ;
        RECT 29.625 2.815 29.795 2.985 ;
        RECT 27.470 2.135 27.640 2.305 ;
        RECT 28.265 2.135 28.435 2.305 ;
        RECT 32.250 2.395 32.420 2.565 ;
        RECT 17.835 0.915 18.005 1.085 ;
        RECT 33.055 2.025 33.225 2.195 ;
        RECT 32.625 0.915 32.795 1.085 ;
        RECT 34.050 2.765 34.220 2.935 ;
        RECT 35.040 2.765 35.210 2.935 ;
        RECT 39.755 2.815 39.925 2.985 ;
        RECT 41.620 3.835 41.790 4.005 ;
        RECT 43.830 3.835 44.000 4.005 ;
        RECT 41.790 2.475 41.960 2.645 ;
        RECT 42.745 2.640 42.800 2.645 ;
        RECT 42.630 2.475 42.800 2.640 ;
        RECT 42.630 2.470 42.745 2.475 ;
        RECT 43.150 2.475 43.320 2.645 ;
        RECT 45.790 3.155 45.960 3.325 ;
        RECT 46.210 2.815 46.380 2.985 ;
        RECT 44.055 2.135 44.225 2.305 ;
        RECT 44.850 2.135 45.020 2.305 ;
        RECT 48.835 2.395 49.005 2.565 ;
        RECT 34.420 0.915 34.590 1.085 ;
        RECT 49.640 2.025 49.810 2.195 ;
        RECT 49.210 0.915 49.380 1.085 ;
        RECT 50.635 2.765 50.805 2.935 ;
        RECT 51.625 2.765 51.795 2.935 ;
        RECT 56.340 2.815 56.510 2.985 ;
        RECT 58.205 3.835 58.375 4.005 ;
        RECT 60.415 3.835 60.585 4.005 ;
        RECT 58.375 2.475 58.545 2.645 ;
        RECT 59.330 2.640 59.385 2.645 ;
        RECT 59.215 2.475 59.385 2.640 ;
        RECT 59.215 2.470 59.330 2.475 ;
        RECT 59.735 2.475 59.905 2.645 ;
        RECT 62.375 3.155 62.545 3.325 ;
        RECT 62.795 2.815 62.965 2.985 ;
        RECT 60.640 2.135 60.810 2.305 ;
        RECT 61.435 2.135 61.605 2.305 ;
        RECT 65.420 2.395 65.590 2.565 ;
        RECT 51.005 0.915 51.175 1.085 ;
        RECT 66.225 2.025 66.395 2.195 ;
        RECT 65.795 0.915 65.965 1.085 ;
        RECT 67.220 2.765 67.390 2.935 ;
        RECT 68.210 2.765 68.380 2.935 ;
        RECT 72.920 2.815 73.090 2.985 ;
        RECT 74.785 3.835 74.955 4.005 ;
        RECT 76.995 3.835 77.165 4.005 ;
        RECT 74.955 2.475 75.125 2.645 ;
        RECT 75.910 2.640 75.965 2.645 ;
        RECT 75.795 2.475 75.965 2.640 ;
        RECT 75.795 2.470 75.910 2.475 ;
        RECT 76.315 2.475 76.485 2.645 ;
        RECT 78.955 3.155 79.125 3.325 ;
        RECT 79.375 2.815 79.545 2.985 ;
        RECT 77.220 2.135 77.390 2.305 ;
        RECT 78.015 2.135 78.185 2.305 ;
        RECT 82.000 2.395 82.170 2.565 ;
        RECT 67.590 0.915 67.760 1.085 ;
        RECT 82.805 2.025 82.975 2.195 ;
        RECT 82.375 0.915 82.545 1.085 ;
        RECT 83.800 2.765 83.970 2.935 ;
        RECT 84.790 2.765 84.960 2.935 ;
        RECT 84.170 0.915 84.340 1.085 ;
      LAYER met1 ;
        RECT 1.525 7.765 1.815 7.995 ;
        RECT 4.755 7.765 5.045 7.995 ;
        RECT 15.980 7.765 16.270 7.995 ;
        RECT 17.775 7.765 18.065 7.995 ;
        RECT 18.765 7.765 19.055 7.995 ;
        RECT 21.340 7.765 21.630 7.995 ;
        RECT 32.565 7.765 32.855 7.995 ;
        RECT 34.360 7.765 34.650 7.995 ;
        RECT 35.350 7.765 35.640 7.995 ;
        RECT 37.925 7.765 38.215 7.995 ;
        RECT 49.150 7.765 49.440 7.995 ;
        RECT 50.945 7.765 51.235 7.995 ;
        RECT 51.935 7.765 52.225 7.995 ;
        RECT 54.510 7.765 54.800 7.995 ;
        RECT 65.735 7.765 66.025 7.995 ;
        RECT 67.530 7.765 67.820 7.995 ;
        RECT 68.520 7.765 68.810 7.995 ;
        RECT 71.090 7.765 71.380 7.995 ;
        RECT 82.315 7.765 82.605 7.995 ;
        RECT 84.110 7.765 84.400 7.995 ;
        RECT 85.100 7.765 85.390 7.995 ;
        RECT 1.585 7.305 1.755 7.765 ;
        RECT 4.815 7.365 4.985 7.765 ;
        RECT 1.495 7.025 1.835 7.305 ;
        RECT 4.715 6.995 5.085 7.365 ;
        RECT 16.040 7.290 16.210 7.765 ;
        RECT 16.040 7.255 17.630 7.290 ;
        RECT 15.980 7.120 17.630 7.255 ;
        RECT 15.980 7.025 16.270 7.120 ;
        RECT 5.215 6.885 5.555 6.910 ;
        RECT 16.435 6.885 16.760 6.980 ;
        RECT 5.185 6.855 5.555 6.885 ;
        RECT 16.410 6.855 16.760 6.885 ;
        RECT 5.015 6.685 5.555 6.855 ;
        RECT 16.240 6.685 16.760 6.855 ;
        RECT 5.185 6.655 5.555 6.685 ;
        RECT 16.410 6.655 16.760 6.685 ;
        RECT 5.215 6.630 5.555 6.655 ;
        RECT 1.120 6.485 1.460 6.565 ;
        RECT 15.635 6.515 15.955 6.605 ;
        RECT 15.605 6.485 15.955 6.515 ;
        RECT 0.980 6.315 1.460 6.485 ;
        RECT 15.435 6.315 15.955 6.485 ;
        RECT 1.120 6.285 1.460 6.315 ;
        RECT 15.605 6.285 15.955 6.315 ;
        RECT 15.635 6.280 15.955 6.285 ;
        RECT 17.460 6.145 17.630 7.120 ;
        RECT 17.835 6.515 18.005 7.765 ;
        RECT 18.825 6.980 18.995 7.765 ;
        RECT 21.400 7.365 21.570 7.765 ;
        RECT 21.300 6.995 21.670 7.365 ;
        RECT 32.625 7.290 32.795 7.765 ;
        RECT 32.625 7.255 34.215 7.290 ;
        RECT 32.565 7.120 34.215 7.255 ;
        RECT 32.565 7.025 32.855 7.120 ;
        RECT 18.825 6.655 19.150 6.980 ;
        RECT 21.800 6.885 22.140 6.910 ;
        RECT 33.020 6.885 33.345 6.980 ;
        RECT 21.770 6.855 22.140 6.885 ;
        RECT 32.995 6.855 33.345 6.885 ;
        RECT 21.600 6.685 22.140 6.855 ;
        RECT 32.825 6.685 33.345 6.855 ;
        RECT 21.770 6.655 22.140 6.685 ;
        RECT 32.995 6.655 33.345 6.685 ;
        RECT 18.825 6.515 18.995 6.655 ;
        RECT 21.800 6.630 22.140 6.655 ;
        RECT 32.220 6.515 32.540 6.605 ;
        RECT 17.775 6.485 18.065 6.515 ;
        RECT 17.775 6.325 18.625 6.485 ;
        RECT 17.775 6.320 18.165 6.325 ;
        RECT 17.775 6.285 18.065 6.320 ;
        RECT 18.455 6.145 18.625 6.325 ;
        RECT 18.765 6.285 19.055 6.515 ;
        RECT 32.190 6.485 32.540 6.515 ;
        RECT 32.020 6.315 32.540 6.485 ;
        RECT 32.190 6.285 32.540 6.315 ;
        RECT 32.220 6.280 32.540 6.285 ;
        RECT 34.045 6.145 34.215 7.120 ;
        RECT 34.420 6.515 34.590 7.765 ;
        RECT 35.410 6.980 35.580 7.765 ;
        RECT 37.985 7.365 38.155 7.765 ;
        RECT 37.885 6.995 38.255 7.365 ;
        RECT 49.210 7.290 49.380 7.765 ;
        RECT 49.210 7.255 50.800 7.290 ;
        RECT 49.150 7.120 50.800 7.255 ;
        RECT 49.150 7.025 49.440 7.120 ;
        RECT 35.410 6.655 35.735 6.980 ;
        RECT 38.385 6.885 38.725 6.910 ;
        RECT 49.605 6.885 49.930 6.980 ;
        RECT 38.355 6.855 38.725 6.885 ;
        RECT 49.580 6.855 49.930 6.885 ;
        RECT 38.185 6.685 38.725 6.855 ;
        RECT 49.410 6.685 49.930 6.855 ;
        RECT 38.355 6.655 38.725 6.685 ;
        RECT 49.580 6.655 49.930 6.685 ;
        RECT 35.410 6.515 35.580 6.655 ;
        RECT 38.385 6.630 38.725 6.655 ;
        RECT 48.805 6.515 49.125 6.605 ;
        RECT 34.360 6.485 34.650 6.515 ;
        RECT 34.360 6.325 35.210 6.485 ;
        RECT 34.360 6.320 34.750 6.325 ;
        RECT 34.360 6.285 34.650 6.320 ;
        RECT 35.040 6.145 35.210 6.325 ;
        RECT 35.350 6.285 35.640 6.515 ;
        RECT 48.775 6.485 49.125 6.515 ;
        RECT 48.605 6.315 49.125 6.485 ;
        RECT 48.775 6.285 49.125 6.315 ;
        RECT 48.805 6.280 49.125 6.285 ;
        RECT 50.630 6.145 50.800 7.120 ;
        RECT 51.005 6.515 51.175 7.765 ;
        RECT 51.995 6.980 52.165 7.765 ;
        RECT 54.570 7.365 54.740 7.765 ;
        RECT 54.470 6.995 54.840 7.365 ;
        RECT 65.795 7.290 65.965 7.765 ;
        RECT 65.795 7.255 67.385 7.290 ;
        RECT 65.735 7.120 67.385 7.255 ;
        RECT 65.735 7.025 66.025 7.120 ;
        RECT 51.995 6.655 52.320 6.980 ;
        RECT 54.970 6.885 55.310 6.910 ;
        RECT 66.190 6.885 66.515 6.980 ;
        RECT 54.940 6.855 55.310 6.885 ;
        RECT 66.165 6.855 66.515 6.885 ;
        RECT 54.770 6.685 55.310 6.855 ;
        RECT 65.995 6.685 66.515 6.855 ;
        RECT 54.940 6.655 55.310 6.685 ;
        RECT 66.165 6.655 66.515 6.685 ;
        RECT 51.995 6.515 52.165 6.655 ;
        RECT 54.970 6.630 55.310 6.655 ;
        RECT 65.390 6.515 65.710 6.605 ;
        RECT 50.945 6.485 51.235 6.515 ;
        RECT 50.945 6.325 51.795 6.485 ;
        RECT 50.945 6.320 51.335 6.325 ;
        RECT 50.945 6.285 51.235 6.320 ;
        RECT 51.625 6.145 51.795 6.325 ;
        RECT 51.935 6.285 52.225 6.515 ;
        RECT 65.360 6.485 65.710 6.515 ;
        RECT 65.190 6.315 65.710 6.485 ;
        RECT 65.360 6.285 65.710 6.315 ;
        RECT 65.390 6.280 65.710 6.285 ;
        RECT 67.215 6.145 67.385 7.120 ;
        RECT 67.590 6.515 67.760 7.765 ;
        RECT 68.580 6.980 68.750 7.765 ;
        RECT 71.150 7.365 71.320 7.765 ;
        RECT 71.050 6.995 71.420 7.365 ;
        RECT 82.375 7.290 82.545 7.765 ;
        RECT 82.375 7.255 83.965 7.290 ;
        RECT 82.315 7.120 83.965 7.255 ;
        RECT 82.315 7.025 82.605 7.120 ;
        RECT 68.580 6.655 68.905 6.980 ;
        RECT 71.550 6.885 71.890 6.910 ;
        RECT 82.770 6.885 83.095 6.980 ;
        RECT 71.520 6.855 71.890 6.885 ;
        RECT 82.745 6.855 83.095 6.885 ;
        RECT 71.350 6.685 71.890 6.855 ;
        RECT 82.575 6.685 83.095 6.855 ;
        RECT 71.520 6.655 71.890 6.685 ;
        RECT 82.745 6.655 83.095 6.685 ;
        RECT 68.580 6.515 68.750 6.655 ;
        RECT 71.550 6.630 71.890 6.655 ;
        RECT 81.970 6.515 82.290 6.605 ;
        RECT 67.530 6.485 67.820 6.515 ;
        RECT 67.530 6.325 68.380 6.485 ;
        RECT 67.530 6.320 67.920 6.325 ;
        RECT 67.530 6.285 67.820 6.320 ;
        RECT 68.210 6.145 68.380 6.325 ;
        RECT 68.520 6.285 68.810 6.515 ;
        RECT 81.940 6.485 82.290 6.515 ;
        RECT 81.770 6.315 82.290 6.485 ;
        RECT 81.940 6.285 82.290 6.315 ;
        RECT 81.970 6.280 82.290 6.285 ;
        RECT 83.795 6.145 83.965 7.120 ;
        RECT 84.170 6.515 84.340 7.765 ;
        RECT 85.160 7.625 85.330 7.765 ;
        RECT 85.125 7.300 85.450 7.625 ;
        RECT 85.160 6.515 85.330 7.300 ;
        RECT 84.110 6.485 84.400 6.515 ;
        RECT 84.110 6.325 84.960 6.485 ;
        RECT 84.110 6.320 84.500 6.325 ;
        RECT 84.110 6.285 84.400 6.320 ;
        RECT 84.790 6.145 84.960 6.325 ;
        RECT 85.100 6.285 85.390 6.515 ;
        RECT 17.405 6.115 17.695 6.145 ;
        RECT 18.395 6.115 18.685 6.145 ;
        RECT 33.990 6.115 34.280 6.145 ;
        RECT 34.980 6.115 35.270 6.145 ;
        RECT 50.575 6.115 50.865 6.145 ;
        RECT 51.565 6.115 51.855 6.145 ;
        RECT 67.160 6.115 67.450 6.145 ;
        RECT 68.150 6.115 68.440 6.145 ;
        RECT 83.740 6.115 84.030 6.145 ;
        RECT 84.730 6.115 85.020 6.145 ;
        RECT 8.900 6.030 9.190 6.075 ;
        RECT 9.565 6.030 9.885 6.090 ;
        RECT 8.900 5.890 9.885 6.030 ;
        RECT 8.900 5.845 9.190 5.890 ;
        RECT 9.565 5.830 9.885 5.890 ;
        RECT 10.585 5.830 10.905 6.090 ;
        RECT 11.280 5.845 11.570 6.075 ;
        RECT 11.945 6.030 12.265 6.090 ;
        RECT 11.945 5.890 12.540 6.030 ;
        RECT 17.405 5.945 17.865 6.115 ;
        RECT 18.395 5.945 18.855 6.115 ;
        RECT 25.485 6.030 25.775 6.075 ;
        RECT 26.150 6.030 26.470 6.090 ;
        RECT 17.405 5.915 17.695 5.945 ;
        RECT 18.395 5.915 18.685 5.945 ;
        RECT 25.485 5.890 26.470 6.030 ;
        RECT 9.655 5.690 9.795 5.830 ;
        RECT 11.355 5.690 11.495 5.845 ;
        RECT 11.945 5.830 12.265 5.890 ;
        RECT 25.485 5.845 25.775 5.890 ;
        RECT 26.150 5.830 26.470 5.890 ;
        RECT 27.170 5.830 27.490 6.090 ;
        RECT 27.865 5.845 28.155 6.075 ;
        RECT 28.530 6.030 28.850 6.090 ;
        RECT 28.530 5.890 29.125 6.030 ;
        RECT 33.990 5.945 34.450 6.115 ;
        RECT 34.980 5.945 35.440 6.115 ;
        RECT 42.070 6.030 42.360 6.075 ;
        RECT 42.735 6.030 43.055 6.090 ;
        RECT 33.990 5.915 34.280 5.945 ;
        RECT 34.980 5.915 35.270 5.945 ;
        RECT 42.070 5.890 43.055 6.030 ;
        RECT 9.655 5.550 11.495 5.690 ;
        RECT 26.240 5.690 26.380 5.830 ;
        RECT 27.940 5.690 28.080 5.845 ;
        RECT 28.530 5.830 28.850 5.890 ;
        RECT 42.070 5.845 42.360 5.890 ;
        RECT 42.735 5.830 43.055 5.890 ;
        RECT 43.755 5.830 44.075 6.090 ;
        RECT 44.450 5.845 44.740 6.075 ;
        RECT 45.115 6.030 45.435 6.090 ;
        RECT 45.115 5.890 45.710 6.030 ;
        RECT 50.575 5.945 51.035 6.115 ;
        RECT 51.565 5.945 52.025 6.115 ;
        RECT 58.655 6.030 58.945 6.075 ;
        RECT 59.320 6.030 59.640 6.090 ;
        RECT 50.575 5.915 50.865 5.945 ;
        RECT 51.565 5.915 51.855 5.945 ;
        RECT 58.655 5.890 59.640 6.030 ;
        RECT 26.240 5.550 28.080 5.690 ;
        RECT 42.825 5.690 42.965 5.830 ;
        RECT 44.525 5.690 44.665 5.845 ;
        RECT 45.115 5.830 45.435 5.890 ;
        RECT 58.655 5.845 58.945 5.890 ;
        RECT 59.320 5.830 59.640 5.890 ;
        RECT 60.340 5.830 60.660 6.090 ;
        RECT 61.035 5.845 61.325 6.075 ;
        RECT 61.700 6.030 62.020 6.090 ;
        RECT 61.700 5.890 62.295 6.030 ;
        RECT 67.160 5.945 67.620 6.115 ;
        RECT 68.150 5.945 68.610 6.115 ;
        RECT 75.235 6.030 75.525 6.075 ;
        RECT 75.900 6.030 76.220 6.090 ;
        RECT 67.160 5.915 67.450 5.945 ;
        RECT 68.150 5.915 68.440 5.945 ;
        RECT 75.235 5.890 76.220 6.030 ;
        RECT 42.825 5.550 44.665 5.690 ;
        RECT 59.410 5.690 59.550 5.830 ;
        RECT 61.110 5.690 61.250 5.845 ;
        RECT 61.700 5.830 62.020 5.890 ;
        RECT 75.235 5.845 75.525 5.890 ;
        RECT 75.900 5.830 76.220 5.890 ;
        RECT 76.920 5.830 77.240 6.090 ;
        RECT 77.615 5.845 77.905 6.075 ;
        RECT 78.280 6.030 78.600 6.090 ;
        RECT 78.280 5.890 78.875 6.030 ;
        RECT 83.740 5.945 84.200 6.115 ;
        RECT 84.730 5.945 85.190 6.115 ;
        RECT 83.740 5.915 84.030 5.945 ;
        RECT 84.730 5.915 85.020 5.945 ;
        RECT 59.410 5.550 61.250 5.690 ;
        RECT 75.990 5.690 76.130 5.830 ;
        RECT 77.690 5.690 77.830 5.845 ;
        RECT 78.280 5.830 78.600 5.890 ;
        RECT 75.990 5.550 77.830 5.690 ;
        RECT 7.200 5.010 7.490 5.055 ;
        RECT 9.905 5.010 10.225 5.070 ;
        RECT 7.200 4.870 10.225 5.010 ;
        RECT 7.200 4.825 7.490 4.870 ;
        RECT 9.905 4.810 10.225 4.870 ;
        RECT 12.640 4.810 13.285 5.070 ;
        RECT 23.785 5.010 24.075 5.055 ;
        RECT 26.490 5.010 26.810 5.070 ;
        RECT 23.785 4.870 26.810 5.010 ;
        RECT 23.785 4.825 24.075 4.870 ;
        RECT 26.490 4.810 26.810 4.870 ;
        RECT 29.225 4.810 29.870 5.070 ;
        RECT 40.370 5.010 40.660 5.055 ;
        RECT 43.075 5.010 43.395 5.070 ;
        RECT 40.370 4.870 43.395 5.010 ;
        RECT 40.370 4.825 40.660 4.870 ;
        RECT 43.075 4.810 43.395 4.870 ;
        RECT 45.810 4.810 46.455 5.070 ;
        RECT 56.955 5.010 57.245 5.055 ;
        RECT 59.660 5.010 59.980 5.070 ;
        RECT 56.955 4.870 59.980 5.010 ;
        RECT 56.955 4.825 57.245 4.870 ;
        RECT 59.660 4.810 59.980 4.870 ;
        RECT 62.395 4.810 63.040 5.070 ;
        RECT 73.535 5.010 73.825 5.055 ;
        RECT 76.240 5.010 76.560 5.070 ;
        RECT 73.535 4.870 76.560 5.010 ;
        RECT 73.535 4.825 73.825 4.870 ;
        RECT 76.240 4.810 76.560 4.870 ;
        RECT 78.975 4.810 79.620 5.070 ;
        RECT 8.390 3.990 8.680 4.035 ;
        RECT 10.600 3.990 10.890 4.035 ;
        RECT 11.265 3.990 11.585 4.050 ;
        RECT 8.390 3.850 11.585 3.990 ;
        RECT 8.390 3.805 8.680 3.850 ;
        RECT 10.600 3.805 10.890 3.850 ;
        RECT 11.265 3.790 11.585 3.850 ;
        RECT 24.975 3.990 25.265 4.035 ;
        RECT 27.185 3.990 27.475 4.035 ;
        RECT 27.850 3.990 28.170 4.050 ;
        RECT 24.975 3.850 28.170 3.990 ;
        RECT 24.975 3.805 25.265 3.850 ;
        RECT 27.185 3.805 27.475 3.850 ;
        RECT 27.850 3.790 28.170 3.850 ;
        RECT 41.560 3.990 41.850 4.035 ;
        RECT 43.770 3.990 44.060 4.035 ;
        RECT 44.435 3.990 44.755 4.050 ;
        RECT 41.560 3.850 44.755 3.990 ;
        RECT 41.560 3.805 41.850 3.850 ;
        RECT 43.770 3.805 44.060 3.850 ;
        RECT 44.435 3.790 44.755 3.850 ;
        RECT 58.145 3.990 58.435 4.035 ;
        RECT 60.355 3.990 60.645 4.035 ;
        RECT 61.020 3.990 61.340 4.050 ;
        RECT 58.145 3.850 61.340 3.990 ;
        RECT 58.145 3.805 58.435 3.850 ;
        RECT 60.355 3.805 60.645 3.850 ;
        RECT 61.020 3.790 61.340 3.850 ;
        RECT 74.725 3.990 75.015 4.035 ;
        RECT 76.935 3.990 77.225 4.035 ;
        RECT 77.600 3.990 77.920 4.050 ;
        RECT 74.725 3.850 77.920 3.990 ;
        RECT 74.725 3.805 75.015 3.850 ;
        RECT 76.935 3.805 77.225 3.850 ;
        RECT 77.600 3.790 77.920 3.850 ;
        RECT 10.585 3.310 10.905 3.370 ;
        RECT 12.560 3.310 12.850 3.355 ;
        RECT 13.380 3.325 13.705 3.510 ;
        RECT 13.280 3.310 13.705 3.325 ;
        RECT 10.585 3.185 13.705 3.310 ;
        RECT 27.170 3.310 27.490 3.370 ;
        RECT 29.145 3.310 29.435 3.355 ;
        RECT 29.965 3.325 30.290 3.510 ;
        RECT 29.865 3.310 30.290 3.325 ;
        RECT 27.170 3.185 30.290 3.310 ;
        RECT 43.755 3.310 44.075 3.370 ;
        RECT 45.730 3.310 46.020 3.355 ;
        RECT 46.550 3.325 46.875 3.510 ;
        RECT 46.450 3.310 46.875 3.325 ;
        RECT 43.755 3.185 46.875 3.310 ;
        RECT 60.340 3.310 60.660 3.370 ;
        RECT 62.315 3.310 62.605 3.355 ;
        RECT 63.135 3.325 63.460 3.510 ;
        RECT 63.035 3.310 63.460 3.325 ;
        RECT 60.340 3.185 63.460 3.310 ;
        RECT 76.920 3.310 77.240 3.370 ;
        RECT 78.895 3.310 79.185 3.355 ;
        RECT 79.715 3.325 80.040 3.510 ;
        RECT 79.615 3.310 80.040 3.325 ;
        RECT 76.920 3.185 80.040 3.310 ;
        RECT 10.585 3.170 13.420 3.185 ;
        RECT 27.170 3.170 30.005 3.185 ;
        RECT 43.755 3.170 46.590 3.185 ;
        RECT 60.340 3.170 63.175 3.185 ;
        RECT 76.920 3.170 79.755 3.185 ;
        RECT 10.585 3.110 10.905 3.170 ;
        RECT 12.560 3.125 12.850 3.170 ;
        RECT 27.170 3.110 27.490 3.170 ;
        RECT 29.145 3.125 29.435 3.170 ;
        RECT 43.755 3.110 44.075 3.170 ;
        RECT 45.730 3.125 46.020 3.170 ;
        RECT 60.340 3.110 60.660 3.170 ;
        RECT 62.315 3.125 62.605 3.170 ;
        RECT 76.920 3.110 77.240 3.170 ;
        RECT 78.895 3.125 79.185 3.170 ;
        RECT 6.525 2.970 6.815 3.015 ;
        RECT 11.265 2.970 11.585 3.030 ;
        RECT 12.965 2.970 13.285 3.030 ;
        RECT 6.525 2.830 11.585 2.970 ;
        RECT 12.690 2.830 13.285 2.970 ;
        RECT 23.110 2.970 23.400 3.015 ;
        RECT 27.850 2.970 28.170 3.030 ;
        RECT 29.550 2.970 29.870 3.030 ;
        RECT 6.525 2.785 6.815 2.830 ;
        RECT 11.265 2.770 11.585 2.830 ;
        RECT 12.965 2.770 13.285 2.830 ;
        RECT 17.405 2.935 17.695 2.965 ;
        RECT 18.355 2.935 18.685 2.965 ;
        RECT 8.560 2.445 8.850 2.675 ;
        RECT 9.225 2.670 9.545 2.685 ;
        RECT 9.575 2.670 9.690 2.675 ;
        RECT 9.225 2.630 9.690 2.670 ;
        RECT 9.905 2.630 10.225 2.690 ;
        RECT 11.355 2.630 11.495 2.770 ;
        RECT 17.405 2.765 17.865 2.935 ;
        RECT 18.355 2.765 18.855 2.935 ;
        RECT 23.110 2.830 28.170 2.970 ;
        RECT 29.275 2.830 29.870 2.970 ;
        RECT 39.695 2.970 39.985 3.015 ;
        RECT 44.435 2.970 44.755 3.030 ;
        RECT 46.135 2.970 46.455 3.030 ;
        RECT 23.110 2.785 23.400 2.830 ;
        RECT 27.850 2.770 28.170 2.830 ;
        RECT 29.550 2.770 29.870 2.830 ;
        RECT 33.990 2.935 34.280 2.965 ;
        RECT 34.940 2.935 35.270 2.965 ;
        RECT 17.405 2.735 17.695 2.765 ;
        RECT 18.355 2.735 18.685 2.765 ;
        RECT 9.110 2.625 9.120 2.630 ;
        RECT 9.225 2.625 9.705 2.630 ;
        RECT 9.110 2.490 9.705 2.625 ;
        RECT 9.905 2.490 10.500 2.630 ;
        RECT 11.355 2.490 11.835 2.630 ;
        RECT 15.635 2.595 15.955 2.685 ;
        RECT 15.605 2.565 15.955 2.595 ;
        RECT 9.120 2.485 9.690 2.490 ;
        RECT 9.225 2.445 9.690 2.485 ;
        RECT 8.635 2.290 8.775 2.445 ;
        RECT 9.225 2.440 9.575 2.445 ;
        RECT 9.225 2.425 9.545 2.440 ;
        RECT 9.905 2.430 10.225 2.490 ;
        RECT 10.925 2.335 11.245 2.350 ;
        RECT 11.695 2.335 11.835 2.490 ;
        RECT 15.320 2.395 15.955 2.565 ;
        RECT 15.605 2.365 15.955 2.395 ;
        RECT 10.825 2.290 11.245 2.335 ;
        RECT 8.635 2.150 11.245 2.290 ;
        RECT 10.825 2.105 11.245 2.150 ;
        RECT 11.620 2.105 11.910 2.335 ;
        RECT 13.965 2.195 14.290 2.320 ;
        RECT 16.410 2.195 16.760 2.315 ;
        RECT 10.925 2.090 11.245 2.105 ;
        RECT 13.965 2.025 16.760 2.195 ;
        RECT 13.965 1.995 14.290 2.025 ;
        RECT 16.410 1.965 16.760 2.025 ;
        RECT 15.980 1.825 16.270 1.855 ;
        RECT 17.465 1.825 17.630 2.735 ;
        RECT 17.775 2.565 18.065 2.595 ;
        RECT 18.355 2.565 18.545 2.735 ;
        RECT 17.775 2.395 18.545 2.565 ;
        RECT 25.145 2.445 25.435 2.675 ;
        RECT 25.810 2.670 26.130 2.685 ;
        RECT 26.160 2.670 26.275 2.675 ;
        RECT 25.810 2.630 26.275 2.670 ;
        RECT 26.490 2.630 26.810 2.690 ;
        RECT 27.940 2.630 28.080 2.770 ;
        RECT 33.990 2.765 34.450 2.935 ;
        RECT 34.940 2.765 35.440 2.935 ;
        RECT 39.695 2.830 44.755 2.970 ;
        RECT 45.860 2.830 46.455 2.970 ;
        RECT 56.280 2.970 56.570 3.015 ;
        RECT 61.020 2.970 61.340 3.030 ;
        RECT 62.720 2.970 63.040 3.030 ;
        RECT 39.695 2.785 39.985 2.830 ;
        RECT 44.435 2.770 44.755 2.830 ;
        RECT 46.135 2.770 46.455 2.830 ;
        RECT 50.575 2.935 50.865 2.965 ;
        RECT 51.525 2.935 51.855 2.965 ;
        RECT 33.990 2.735 34.280 2.765 ;
        RECT 34.940 2.735 35.270 2.765 ;
        RECT 25.695 2.625 25.705 2.630 ;
        RECT 25.810 2.625 26.290 2.630 ;
        RECT 25.695 2.490 26.290 2.625 ;
        RECT 26.490 2.490 27.085 2.630 ;
        RECT 27.940 2.490 28.420 2.630 ;
        RECT 32.220 2.595 32.540 2.685 ;
        RECT 32.190 2.565 32.540 2.595 ;
        RECT 25.705 2.485 26.275 2.490 ;
        RECT 25.810 2.445 26.275 2.485 ;
        RECT 17.775 2.365 18.065 2.395 ;
        RECT 15.980 1.655 17.630 1.825 ;
        RECT 15.980 1.625 16.270 1.655 ;
        RECT 16.040 1.115 16.210 1.625 ;
        RECT 17.835 1.115 18.005 2.365 ;
        RECT 25.220 2.290 25.360 2.445 ;
        RECT 25.810 2.440 26.160 2.445 ;
        RECT 25.810 2.425 26.130 2.440 ;
        RECT 26.490 2.430 26.810 2.490 ;
        RECT 27.510 2.335 27.830 2.350 ;
        RECT 28.280 2.335 28.420 2.490 ;
        RECT 31.905 2.395 32.540 2.565 ;
        RECT 32.190 2.365 32.540 2.395 ;
        RECT 27.410 2.290 27.830 2.335 ;
        RECT 25.220 2.150 27.830 2.290 ;
        RECT 27.410 2.105 27.830 2.150 ;
        RECT 28.205 2.105 28.495 2.335 ;
        RECT 30.550 2.195 30.875 2.320 ;
        RECT 32.995 2.195 33.345 2.315 ;
        RECT 27.510 2.090 27.830 2.105 ;
        RECT 30.550 2.025 33.345 2.195 ;
        RECT 30.550 1.995 30.875 2.025 ;
        RECT 32.995 1.965 33.345 2.025 ;
        RECT 32.565 1.825 32.855 1.855 ;
        RECT 34.050 1.825 34.215 2.735 ;
        RECT 34.360 2.565 34.650 2.595 ;
        RECT 34.940 2.565 35.130 2.735 ;
        RECT 34.360 2.395 35.130 2.565 ;
        RECT 41.730 2.445 42.020 2.675 ;
        RECT 42.395 2.670 42.715 2.685 ;
        RECT 42.745 2.670 42.860 2.675 ;
        RECT 42.395 2.630 42.860 2.670 ;
        RECT 43.075 2.630 43.395 2.690 ;
        RECT 44.525 2.630 44.665 2.770 ;
        RECT 50.575 2.765 51.035 2.935 ;
        RECT 51.525 2.765 52.025 2.935 ;
        RECT 56.280 2.830 61.340 2.970 ;
        RECT 62.445 2.830 63.040 2.970 ;
        RECT 72.860 2.970 73.150 3.015 ;
        RECT 77.600 2.970 77.920 3.030 ;
        RECT 79.300 2.970 79.620 3.030 ;
        RECT 56.280 2.785 56.570 2.830 ;
        RECT 61.020 2.770 61.340 2.830 ;
        RECT 62.720 2.770 63.040 2.830 ;
        RECT 67.160 2.935 67.450 2.965 ;
        RECT 68.110 2.935 68.440 2.965 ;
        RECT 50.575 2.735 50.865 2.765 ;
        RECT 51.525 2.735 51.855 2.765 ;
        RECT 42.280 2.625 42.290 2.630 ;
        RECT 42.395 2.625 42.875 2.630 ;
        RECT 42.280 2.490 42.875 2.625 ;
        RECT 43.075 2.490 43.670 2.630 ;
        RECT 44.525 2.490 45.005 2.630 ;
        RECT 48.805 2.595 49.125 2.685 ;
        RECT 48.775 2.565 49.125 2.595 ;
        RECT 42.290 2.485 42.860 2.490 ;
        RECT 42.395 2.445 42.860 2.485 ;
        RECT 34.360 2.365 34.650 2.395 ;
        RECT 32.565 1.655 34.215 1.825 ;
        RECT 32.565 1.625 32.855 1.655 ;
        RECT 32.625 1.115 32.795 1.625 ;
        RECT 34.420 1.115 34.590 2.365 ;
        RECT 41.805 2.290 41.945 2.445 ;
        RECT 42.395 2.440 42.745 2.445 ;
        RECT 42.395 2.425 42.715 2.440 ;
        RECT 43.075 2.430 43.395 2.490 ;
        RECT 44.095 2.335 44.415 2.350 ;
        RECT 44.865 2.335 45.005 2.490 ;
        RECT 48.490 2.395 49.125 2.565 ;
        RECT 48.775 2.365 49.125 2.395 ;
        RECT 43.995 2.290 44.415 2.335 ;
        RECT 41.805 2.150 44.415 2.290 ;
        RECT 43.995 2.105 44.415 2.150 ;
        RECT 44.790 2.105 45.080 2.335 ;
        RECT 47.135 2.195 47.460 2.320 ;
        RECT 49.580 2.195 49.930 2.315 ;
        RECT 44.095 2.090 44.415 2.105 ;
        RECT 47.135 2.025 49.930 2.195 ;
        RECT 47.135 1.995 47.460 2.025 ;
        RECT 49.580 1.965 49.930 2.025 ;
        RECT 49.150 1.825 49.440 1.855 ;
        RECT 50.635 1.825 50.800 2.735 ;
        RECT 50.945 2.565 51.235 2.595 ;
        RECT 51.525 2.565 51.715 2.735 ;
        RECT 50.945 2.395 51.715 2.565 ;
        RECT 58.315 2.445 58.605 2.675 ;
        RECT 58.980 2.670 59.300 2.685 ;
        RECT 59.330 2.670 59.445 2.675 ;
        RECT 58.980 2.630 59.445 2.670 ;
        RECT 59.660 2.630 59.980 2.690 ;
        RECT 61.110 2.630 61.250 2.770 ;
        RECT 67.160 2.765 67.620 2.935 ;
        RECT 68.110 2.765 68.610 2.935 ;
        RECT 72.860 2.830 77.920 2.970 ;
        RECT 79.025 2.830 79.620 2.970 ;
        RECT 72.860 2.785 73.150 2.830 ;
        RECT 77.600 2.770 77.920 2.830 ;
        RECT 79.300 2.770 79.620 2.830 ;
        RECT 83.740 2.935 84.030 2.965 ;
        RECT 84.690 2.935 85.020 2.965 ;
        RECT 67.160 2.735 67.450 2.765 ;
        RECT 68.110 2.735 68.440 2.765 ;
        RECT 58.865 2.625 58.875 2.630 ;
        RECT 58.980 2.625 59.460 2.630 ;
        RECT 58.865 2.490 59.460 2.625 ;
        RECT 59.660 2.490 60.255 2.630 ;
        RECT 61.110 2.490 61.590 2.630 ;
        RECT 65.390 2.595 65.710 2.685 ;
        RECT 65.360 2.565 65.710 2.595 ;
        RECT 58.875 2.485 59.445 2.490 ;
        RECT 58.980 2.445 59.445 2.485 ;
        RECT 50.945 2.365 51.235 2.395 ;
        RECT 49.150 1.655 50.800 1.825 ;
        RECT 49.150 1.625 49.440 1.655 ;
        RECT 49.210 1.115 49.380 1.625 ;
        RECT 51.005 1.115 51.175 2.365 ;
        RECT 58.390 2.290 58.530 2.445 ;
        RECT 58.980 2.440 59.330 2.445 ;
        RECT 58.980 2.425 59.300 2.440 ;
        RECT 59.660 2.430 59.980 2.490 ;
        RECT 60.680 2.335 61.000 2.350 ;
        RECT 61.450 2.335 61.590 2.490 ;
        RECT 65.075 2.395 65.710 2.565 ;
        RECT 65.360 2.365 65.710 2.395 ;
        RECT 60.580 2.290 61.000 2.335 ;
        RECT 58.390 2.150 61.000 2.290 ;
        RECT 60.580 2.105 61.000 2.150 ;
        RECT 61.375 2.105 61.665 2.335 ;
        RECT 63.720 2.195 64.045 2.320 ;
        RECT 66.165 2.195 66.515 2.315 ;
        RECT 60.680 2.090 61.000 2.105 ;
        RECT 63.720 2.025 66.515 2.195 ;
        RECT 63.720 1.995 64.045 2.025 ;
        RECT 66.165 1.965 66.515 2.025 ;
        RECT 65.735 1.825 66.025 1.855 ;
        RECT 67.220 1.825 67.385 2.735 ;
        RECT 67.530 2.565 67.820 2.595 ;
        RECT 68.110 2.565 68.300 2.735 ;
        RECT 67.530 2.395 68.300 2.565 ;
        RECT 74.895 2.445 75.185 2.675 ;
        RECT 75.560 2.670 75.880 2.685 ;
        RECT 75.910 2.670 76.025 2.675 ;
        RECT 75.560 2.630 76.025 2.670 ;
        RECT 76.240 2.630 76.560 2.690 ;
        RECT 77.690 2.630 77.830 2.770 ;
        RECT 83.740 2.765 84.200 2.935 ;
        RECT 84.690 2.765 85.190 2.935 ;
        RECT 83.740 2.735 84.030 2.765 ;
        RECT 84.690 2.735 85.020 2.765 ;
        RECT 75.445 2.625 75.455 2.630 ;
        RECT 75.560 2.625 76.040 2.630 ;
        RECT 75.445 2.490 76.040 2.625 ;
        RECT 76.240 2.490 76.835 2.630 ;
        RECT 77.690 2.490 78.170 2.630 ;
        RECT 81.970 2.595 82.290 2.685 ;
        RECT 81.940 2.565 82.290 2.595 ;
        RECT 75.455 2.485 76.025 2.490 ;
        RECT 75.560 2.445 76.025 2.485 ;
        RECT 67.530 2.365 67.820 2.395 ;
        RECT 65.735 1.655 67.385 1.825 ;
        RECT 65.735 1.625 66.025 1.655 ;
        RECT 65.795 1.115 65.965 1.625 ;
        RECT 67.590 1.115 67.760 2.365 ;
        RECT 74.970 2.290 75.110 2.445 ;
        RECT 75.560 2.440 75.910 2.445 ;
        RECT 75.560 2.425 75.880 2.440 ;
        RECT 76.240 2.430 76.560 2.490 ;
        RECT 77.260 2.335 77.580 2.350 ;
        RECT 78.030 2.335 78.170 2.490 ;
        RECT 81.655 2.395 82.290 2.565 ;
        RECT 81.940 2.365 82.290 2.395 ;
        RECT 77.160 2.290 77.580 2.335 ;
        RECT 74.970 2.150 77.580 2.290 ;
        RECT 77.160 2.105 77.580 2.150 ;
        RECT 77.955 2.105 78.245 2.335 ;
        RECT 80.300 2.195 80.625 2.320 ;
        RECT 82.745 2.195 83.095 2.315 ;
        RECT 77.260 2.090 77.580 2.105 ;
        RECT 80.300 2.025 83.095 2.195 ;
        RECT 80.300 1.995 80.625 2.025 ;
        RECT 82.745 1.965 83.095 2.025 ;
        RECT 82.315 1.825 82.605 1.855 ;
        RECT 83.800 1.825 83.965 2.735 ;
        RECT 84.110 2.565 84.400 2.595 ;
        RECT 84.690 2.565 84.880 2.735 ;
        RECT 84.110 2.395 84.880 2.565 ;
        RECT 84.110 2.365 84.400 2.395 ;
        RECT 82.315 1.655 83.965 1.825 ;
        RECT 82.315 1.625 82.605 1.655 ;
        RECT 82.375 1.115 82.545 1.625 ;
        RECT 84.170 1.115 84.340 2.365 ;
        RECT 15.980 0.885 16.270 1.115 ;
        RECT 17.775 0.885 18.065 1.115 ;
        RECT 32.565 0.885 32.855 1.115 ;
        RECT 34.360 0.885 34.650 1.115 ;
        RECT 49.150 0.885 49.440 1.115 ;
        RECT 50.945 0.885 51.235 1.115 ;
        RECT 65.735 0.885 66.025 1.115 ;
        RECT 67.530 0.885 67.820 1.115 ;
        RECT 82.315 0.885 82.605 1.115 ;
        RECT 84.110 0.885 84.400 1.115 ;
      LAYER via ;
        RECT 1.525 7.025 1.805 7.305 ;
        RECT 4.760 7.040 5.040 7.320 ;
        RECT 5.245 6.630 5.525 6.910 ;
        RECT 16.470 6.685 16.730 6.945 ;
        RECT 1.150 6.285 1.430 6.565 ;
        RECT 15.665 6.315 15.925 6.575 ;
        RECT 21.345 7.040 21.625 7.320 ;
        RECT 18.860 6.685 19.120 6.945 ;
        RECT 21.830 6.630 22.110 6.910 ;
        RECT 33.055 6.685 33.315 6.945 ;
        RECT 32.250 6.315 32.510 6.575 ;
        RECT 37.930 7.040 38.210 7.320 ;
        RECT 35.445 6.685 35.705 6.945 ;
        RECT 38.415 6.630 38.695 6.910 ;
        RECT 49.640 6.685 49.900 6.945 ;
        RECT 48.835 6.315 49.095 6.575 ;
        RECT 54.515 7.040 54.795 7.320 ;
        RECT 52.030 6.685 52.290 6.945 ;
        RECT 55.000 6.630 55.280 6.910 ;
        RECT 66.225 6.685 66.485 6.945 ;
        RECT 65.420 6.315 65.680 6.575 ;
        RECT 71.095 7.040 71.375 7.320 ;
        RECT 68.615 6.685 68.875 6.945 ;
        RECT 71.580 6.630 71.860 6.910 ;
        RECT 82.805 6.685 83.065 6.945 ;
        RECT 82.000 6.315 82.260 6.575 ;
        RECT 85.160 7.330 85.420 7.590 ;
        RECT 9.595 5.830 9.855 6.090 ;
        RECT 10.615 5.830 10.875 6.090 ;
        RECT 11.975 5.830 12.235 6.090 ;
        RECT 26.180 5.830 26.440 6.090 ;
        RECT 27.200 5.830 27.460 6.090 ;
        RECT 28.560 5.830 28.820 6.090 ;
        RECT 42.765 5.830 43.025 6.090 ;
        RECT 43.785 5.830 44.045 6.090 ;
        RECT 45.145 5.830 45.405 6.090 ;
        RECT 59.350 5.830 59.610 6.090 ;
        RECT 60.370 5.830 60.630 6.090 ;
        RECT 61.730 5.830 61.990 6.090 ;
        RECT 75.930 5.830 76.190 6.090 ;
        RECT 76.950 5.830 77.210 6.090 ;
        RECT 78.310 5.830 78.570 6.090 ;
        RECT 9.935 4.810 10.195 5.070 ;
        RECT 12.995 4.810 13.255 5.070 ;
        RECT 26.520 4.810 26.780 5.070 ;
        RECT 29.580 4.810 29.840 5.070 ;
        RECT 43.105 4.810 43.365 5.070 ;
        RECT 46.165 4.810 46.425 5.070 ;
        RECT 59.690 4.810 59.950 5.070 ;
        RECT 62.750 4.810 63.010 5.070 ;
        RECT 76.270 4.810 76.530 5.070 ;
        RECT 79.330 4.810 79.590 5.070 ;
        RECT 11.295 3.790 11.555 4.050 ;
        RECT 27.880 3.790 28.140 4.050 ;
        RECT 44.465 3.790 44.725 4.050 ;
        RECT 61.050 3.790 61.310 4.050 ;
        RECT 77.630 3.790 77.890 4.050 ;
        RECT 10.615 3.110 10.875 3.370 ;
        RECT 13.415 3.215 13.675 3.475 ;
        RECT 27.200 3.110 27.460 3.370 ;
        RECT 30.000 3.215 30.260 3.475 ;
        RECT 43.785 3.110 44.045 3.370 ;
        RECT 46.585 3.215 46.845 3.475 ;
        RECT 60.370 3.110 60.630 3.370 ;
        RECT 63.170 3.215 63.430 3.475 ;
        RECT 76.950 3.110 77.210 3.370 ;
        RECT 79.750 3.215 80.010 3.475 ;
        RECT 11.295 2.770 11.555 3.030 ;
        RECT 12.995 2.770 13.255 3.030 ;
        RECT 9.255 2.425 9.515 2.685 ;
        RECT 9.935 2.430 10.195 2.690 ;
        RECT 27.880 2.770 28.140 3.030 ;
        RECT 29.580 2.770 29.840 3.030 ;
        RECT 10.955 2.090 11.215 2.350 ;
        RECT 15.665 2.395 15.925 2.655 ;
        RECT 14.000 2.025 14.260 2.285 ;
        RECT 16.440 1.995 16.730 2.285 ;
        RECT 25.840 2.425 26.100 2.685 ;
        RECT 26.520 2.430 26.780 2.690 ;
        RECT 44.465 2.770 44.725 3.030 ;
        RECT 46.165 2.770 46.425 3.030 ;
        RECT 27.540 2.090 27.800 2.350 ;
        RECT 32.250 2.395 32.510 2.655 ;
        RECT 30.585 2.025 30.845 2.285 ;
        RECT 33.025 1.995 33.315 2.285 ;
        RECT 42.425 2.425 42.685 2.685 ;
        RECT 43.105 2.430 43.365 2.690 ;
        RECT 61.050 2.770 61.310 3.030 ;
        RECT 62.750 2.770 63.010 3.030 ;
        RECT 44.125 2.090 44.385 2.350 ;
        RECT 48.835 2.395 49.095 2.655 ;
        RECT 47.170 2.025 47.430 2.285 ;
        RECT 49.610 1.995 49.900 2.285 ;
        RECT 59.010 2.425 59.270 2.685 ;
        RECT 59.690 2.430 59.950 2.690 ;
        RECT 77.630 2.770 77.890 3.030 ;
        RECT 79.330 2.770 79.590 3.030 ;
        RECT 60.710 2.090 60.970 2.350 ;
        RECT 65.420 2.395 65.680 2.655 ;
        RECT 63.755 2.025 64.015 2.285 ;
        RECT 66.195 1.995 66.485 2.285 ;
        RECT 75.590 2.425 75.850 2.685 ;
        RECT 76.270 2.430 76.530 2.690 ;
        RECT 77.290 2.090 77.550 2.350 ;
        RECT 82.000 2.395 82.260 2.655 ;
        RECT 80.335 2.025 80.595 2.285 ;
        RECT 82.775 1.995 83.065 2.285 ;
      LAYER met2 ;
        RECT 1.205 8.600 85.330 8.770 ;
        RECT 1.205 6.595 1.375 8.600 ;
        RECT 5.300 8.290 15.480 8.460 ;
        RECT 1.525 7.230 1.805 7.335 ;
        RECT 1.525 7.060 2.690 7.230 ;
        RECT 1.525 6.995 1.805 7.060 ;
        RECT 2.520 6.855 2.690 7.060 ;
        RECT 4.715 6.995 5.085 7.365 ;
        RECT 5.300 6.940 5.470 8.290 ;
        RECT 5.245 6.855 5.525 6.940 ;
        RECT 2.520 6.685 5.525 6.855 ;
        RECT 5.245 6.600 5.525 6.685 ;
        RECT 15.320 6.915 15.480 8.290 ;
        RECT 21.885 8.290 32.065 8.460 ;
        RECT 21.300 6.995 21.670 7.365 ;
        RECT 16.435 6.915 16.760 6.980 ;
        RECT 15.320 6.745 16.760 6.915 ;
        RECT 1.150 6.255 1.430 6.595 ;
        RECT 9.570 6.120 9.850 6.145 ;
        RECT 9.570 5.800 9.855 6.120 ;
        RECT 9.570 5.775 9.850 5.800 ;
        RECT 10.615 5.775 10.895 6.145 ;
        RECT 11.975 6.030 12.235 6.120 ;
        RECT 11.355 5.890 12.235 6.030 ;
        RECT 9.935 4.755 10.215 5.125 ;
        RECT 9.255 2.370 9.535 2.740 ;
        RECT 9.995 2.720 10.135 4.755 ;
        RECT 10.675 3.990 10.815 5.775 ;
        RECT 11.355 4.105 11.495 5.890 ;
        RECT 11.975 5.800 12.235 5.890 ;
        RECT 12.995 4.780 13.255 5.100 ;
        RECT 10.675 3.850 11.155 3.990 ;
        RECT 10.595 3.055 10.875 3.425 ;
        RECT 9.935 2.400 10.195 2.720 ;
        RECT 11.015 2.380 11.155 3.850 ;
        RECT 11.295 3.735 11.575 4.105 ;
        RECT 11.295 2.715 11.575 3.085 ;
        RECT 13.055 3.060 13.195 4.780 ;
        RECT 13.380 3.400 13.705 3.510 ;
        RECT 13.380 3.215 14.210 3.400 ;
        RECT 13.380 3.185 13.705 3.215 ;
        RECT 12.995 2.740 13.255 3.060 ;
        RECT 10.955 2.060 11.215 2.380 ;
        RECT 14.040 2.320 14.210 3.215 ;
        RECT 15.320 2.565 15.480 6.745 ;
        RECT 16.435 6.655 16.760 6.745 ;
        RECT 18.825 6.855 19.150 6.980 ;
        RECT 21.885 6.940 22.055 8.290 ;
        RECT 21.830 6.855 22.110 6.940 ;
        RECT 18.825 6.685 22.110 6.855 ;
        RECT 18.825 6.655 19.150 6.685 ;
        RECT 15.635 6.280 15.955 6.605 ;
        RECT 21.830 6.600 22.110 6.685 ;
        RECT 31.905 6.915 32.065 8.290 ;
        RECT 38.470 8.290 48.650 8.460 ;
        RECT 37.885 6.995 38.255 7.365 ;
        RECT 33.020 6.915 33.345 6.980 ;
        RECT 31.905 6.745 33.345 6.915 ;
        RECT 15.665 6.045 15.835 6.280 ;
        RECT 26.155 6.120 26.435 6.145 ;
        RECT 15.665 5.870 15.840 6.045 ;
        RECT 15.665 5.695 16.640 5.870 ;
        RECT 26.155 5.800 26.440 6.120 ;
        RECT 26.155 5.775 26.435 5.800 ;
        RECT 27.200 5.775 27.480 6.145 ;
        RECT 28.560 6.030 28.820 6.120 ;
        RECT 27.940 5.890 28.820 6.030 ;
        RECT 15.635 2.565 15.955 2.685 ;
        RECT 15.320 2.395 15.955 2.565 ;
        RECT 15.635 2.365 15.955 2.395 ;
        RECT 13.965 1.995 14.290 2.320 ;
        RECT 16.465 2.315 16.640 5.695 ;
        RECT 26.520 4.755 26.800 5.125 ;
        RECT 25.840 2.370 26.120 2.740 ;
        RECT 26.580 2.720 26.720 4.755 ;
        RECT 27.260 3.990 27.400 5.775 ;
        RECT 27.940 4.105 28.080 5.890 ;
        RECT 28.560 5.800 28.820 5.890 ;
        RECT 29.580 4.780 29.840 5.100 ;
        RECT 27.260 3.850 27.740 3.990 ;
        RECT 27.180 3.055 27.460 3.425 ;
        RECT 26.520 2.400 26.780 2.720 ;
        RECT 27.600 2.380 27.740 3.850 ;
        RECT 27.880 3.735 28.160 4.105 ;
        RECT 27.880 2.715 28.160 3.085 ;
        RECT 29.640 3.060 29.780 4.780 ;
        RECT 29.965 3.400 30.290 3.510 ;
        RECT 29.965 3.215 30.795 3.400 ;
        RECT 29.965 3.185 30.290 3.215 ;
        RECT 29.580 2.740 29.840 3.060 ;
        RECT 16.410 1.965 16.760 2.315 ;
        RECT 27.540 2.060 27.800 2.380 ;
        RECT 30.625 2.320 30.795 3.215 ;
        RECT 31.905 2.565 32.065 6.745 ;
        RECT 33.020 6.655 33.345 6.745 ;
        RECT 35.410 6.855 35.735 6.980 ;
        RECT 38.470 6.940 38.640 8.290 ;
        RECT 38.415 6.855 38.695 6.940 ;
        RECT 35.410 6.685 38.695 6.855 ;
        RECT 35.410 6.655 35.735 6.685 ;
        RECT 32.220 6.280 32.540 6.605 ;
        RECT 38.415 6.600 38.695 6.685 ;
        RECT 48.490 6.915 48.650 8.290 ;
        RECT 55.055 8.290 65.235 8.460 ;
        RECT 54.470 6.995 54.840 7.365 ;
        RECT 49.605 6.915 49.930 6.980 ;
        RECT 48.490 6.745 49.930 6.915 ;
        RECT 32.250 6.045 32.420 6.280 ;
        RECT 42.740 6.120 43.020 6.145 ;
        RECT 32.250 5.870 32.425 6.045 ;
        RECT 32.250 5.695 33.225 5.870 ;
        RECT 42.740 5.800 43.025 6.120 ;
        RECT 42.740 5.775 43.020 5.800 ;
        RECT 43.785 5.775 44.065 6.145 ;
        RECT 45.145 6.030 45.405 6.120 ;
        RECT 44.525 5.890 45.405 6.030 ;
        RECT 32.220 2.565 32.540 2.685 ;
        RECT 31.905 2.395 32.540 2.565 ;
        RECT 32.220 2.365 32.540 2.395 ;
        RECT 30.550 1.995 30.875 2.320 ;
        RECT 33.050 2.315 33.225 5.695 ;
        RECT 43.105 4.755 43.385 5.125 ;
        RECT 42.425 2.370 42.705 2.740 ;
        RECT 43.165 2.720 43.305 4.755 ;
        RECT 43.845 3.990 43.985 5.775 ;
        RECT 44.525 4.105 44.665 5.890 ;
        RECT 45.145 5.800 45.405 5.890 ;
        RECT 46.165 4.780 46.425 5.100 ;
        RECT 43.845 3.850 44.325 3.990 ;
        RECT 43.765 3.055 44.045 3.425 ;
        RECT 43.105 2.400 43.365 2.720 ;
        RECT 44.185 2.380 44.325 3.850 ;
        RECT 44.465 3.735 44.745 4.105 ;
        RECT 44.465 2.715 44.745 3.085 ;
        RECT 46.225 3.060 46.365 4.780 ;
        RECT 46.550 3.400 46.875 3.510 ;
        RECT 46.550 3.215 47.380 3.400 ;
        RECT 46.550 3.185 46.875 3.215 ;
        RECT 46.165 2.740 46.425 3.060 ;
        RECT 32.995 1.965 33.345 2.315 ;
        RECT 44.125 2.060 44.385 2.380 ;
        RECT 47.210 2.320 47.380 3.215 ;
        RECT 48.490 2.565 48.650 6.745 ;
        RECT 49.605 6.655 49.930 6.745 ;
        RECT 51.995 6.855 52.320 6.980 ;
        RECT 55.055 6.940 55.225 8.290 ;
        RECT 55.000 6.855 55.280 6.940 ;
        RECT 51.995 6.685 55.280 6.855 ;
        RECT 51.995 6.655 52.320 6.685 ;
        RECT 48.805 6.280 49.125 6.605 ;
        RECT 55.000 6.600 55.280 6.685 ;
        RECT 65.075 6.915 65.235 8.290 ;
        RECT 71.635 8.290 81.815 8.460 ;
        RECT 71.050 7.005 71.420 7.365 ;
        RECT 71.050 6.995 71.425 7.005 ;
        RECT 66.190 6.915 66.515 6.980 ;
        RECT 65.075 6.745 66.515 6.915 ;
        RECT 48.835 6.045 49.005 6.280 ;
        RECT 59.325 6.120 59.605 6.145 ;
        RECT 48.835 5.870 49.010 6.045 ;
        RECT 48.835 5.695 49.810 5.870 ;
        RECT 59.325 5.800 59.610 6.120 ;
        RECT 59.325 5.775 59.605 5.800 ;
        RECT 60.370 5.775 60.650 6.145 ;
        RECT 61.730 6.030 61.990 6.120 ;
        RECT 61.110 5.890 61.990 6.030 ;
        RECT 48.805 2.565 49.125 2.685 ;
        RECT 48.490 2.395 49.125 2.565 ;
        RECT 48.805 2.365 49.125 2.395 ;
        RECT 47.135 1.995 47.460 2.320 ;
        RECT 49.635 2.315 49.810 5.695 ;
        RECT 59.690 4.755 59.970 5.125 ;
        RECT 59.010 2.370 59.290 2.740 ;
        RECT 59.750 2.720 59.890 4.755 ;
        RECT 60.430 3.990 60.570 5.775 ;
        RECT 61.110 4.105 61.250 5.890 ;
        RECT 61.730 5.800 61.990 5.890 ;
        RECT 62.750 4.780 63.010 5.100 ;
        RECT 60.430 3.850 60.910 3.990 ;
        RECT 60.350 3.055 60.630 3.425 ;
        RECT 59.690 2.400 59.950 2.720 ;
        RECT 60.770 2.380 60.910 3.850 ;
        RECT 61.050 3.735 61.330 4.105 ;
        RECT 61.050 2.715 61.330 3.085 ;
        RECT 62.810 3.060 62.950 4.780 ;
        RECT 63.135 3.400 63.460 3.510 ;
        RECT 63.135 3.215 63.965 3.400 ;
        RECT 63.135 3.185 63.460 3.215 ;
        RECT 62.750 2.740 63.010 3.060 ;
        RECT 49.580 1.965 49.930 2.315 ;
        RECT 60.710 2.060 60.970 2.380 ;
        RECT 63.795 2.320 63.965 3.215 ;
        RECT 65.075 2.565 65.235 6.745 ;
        RECT 66.190 6.655 66.515 6.745 ;
        RECT 68.580 6.855 68.905 6.980 ;
        RECT 71.635 6.940 71.805 8.290 ;
        RECT 71.580 6.855 71.860 6.940 ;
        RECT 68.580 6.685 71.860 6.855 ;
        RECT 68.580 6.655 68.905 6.685 ;
        RECT 65.390 6.280 65.710 6.605 ;
        RECT 71.580 6.600 71.860 6.685 ;
        RECT 81.655 6.915 81.815 8.290 ;
        RECT 85.160 7.625 85.330 8.600 ;
        RECT 85.125 7.300 85.450 7.625 ;
        RECT 82.770 6.915 83.095 6.980 ;
        RECT 81.655 6.745 83.095 6.915 ;
        RECT 65.420 6.045 65.590 6.280 ;
        RECT 75.905 6.120 76.185 6.145 ;
        RECT 65.420 5.870 65.595 6.045 ;
        RECT 65.420 5.695 66.395 5.870 ;
        RECT 75.905 5.800 76.190 6.120 ;
        RECT 75.905 5.775 76.185 5.800 ;
        RECT 76.950 5.775 77.230 6.145 ;
        RECT 78.310 6.030 78.570 6.120 ;
        RECT 77.690 5.890 78.570 6.030 ;
        RECT 65.390 2.565 65.710 2.685 ;
        RECT 65.075 2.395 65.710 2.565 ;
        RECT 65.390 2.365 65.710 2.395 ;
        RECT 63.720 1.995 64.045 2.320 ;
        RECT 66.220 2.315 66.395 5.695 ;
        RECT 76.270 4.755 76.550 5.125 ;
        RECT 75.590 2.370 75.870 2.740 ;
        RECT 76.330 2.720 76.470 4.755 ;
        RECT 77.010 3.990 77.150 5.775 ;
        RECT 77.690 4.105 77.830 5.890 ;
        RECT 78.310 5.800 78.570 5.890 ;
        RECT 79.330 4.780 79.590 5.100 ;
        RECT 77.010 3.850 77.490 3.990 ;
        RECT 76.930 3.055 77.210 3.425 ;
        RECT 76.270 2.400 76.530 2.720 ;
        RECT 77.350 2.380 77.490 3.850 ;
        RECT 77.630 3.735 77.910 4.105 ;
        RECT 77.630 2.715 77.910 3.085 ;
        RECT 79.390 3.060 79.530 4.780 ;
        RECT 79.715 3.400 80.040 3.510 ;
        RECT 79.715 3.215 80.545 3.400 ;
        RECT 79.715 3.185 80.040 3.215 ;
        RECT 79.330 2.740 79.590 3.060 ;
        RECT 66.165 1.965 66.515 2.315 ;
        RECT 77.290 2.060 77.550 2.380 ;
        RECT 80.375 2.320 80.545 3.215 ;
        RECT 81.655 2.565 81.815 6.745 ;
        RECT 82.770 6.655 83.095 6.745 ;
        RECT 81.970 6.280 82.290 6.605 ;
        RECT 82.000 6.045 82.170 6.280 ;
        RECT 82.000 5.870 82.175 6.045 ;
        RECT 82.000 5.695 82.975 5.870 ;
        RECT 81.970 2.565 82.290 2.685 ;
        RECT 81.655 2.395 82.290 2.565 ;
        RECT 81.970 2.365 82.290 2.395 ;
        RECT 80.300 1.995 80.625 2.320 ;
        RECT 82.800 2.315 82.975 5.695 ;
        RECT 82.745 1.965 83.095 2.315 ;
      LAYER via2 ;
        RECT 4.760 7.040 5.040 7.320 ;
        RECT 21.345 7.040 21.625 7.320 ;
        RECT 9.570 5.820 9.850 6.100 ;
        RECT 10.615 5.820 10.895 6.100 ;
        RECT 9.935 4.800 10.215 5.080 ;
        RECT 10.595 3.100 10.875 3.380 ;
        RECT 9.255 2.415 9.535 2.695 ;
        RECT 11.295 3.780 11.575 4.060 ;
        RECT 11.295 2.760 11.575 3.040 ;
        RECT 37.930 7.040 38.210 7.320 ;
        RECT 26.155 5.820 26.435 6.100 ;
        RECT 27.200 5.820 27.480 6.100 ;
        RECT 26.520 4.800 26.800 5.080 ;
        RECT 27.180 3.100 27.460 3.380 ;
        RECT 25.840 2.415 26.120 2.695 ;
        RECT 27.880 3.780 28.160 4.060 ;
        RECT 27.880 2.760 28.160 3.040 ;
        RECT 54.515 7.040 54.795 7.320 ;
        RECT 42.740 5.820 43.020 6.100 ;
        RECT 43.785 5.820 44.065 6.100 ;
        RECT 43.105 4.800 43.385 5.080 ;
        RECT 43.765 3.100 44.045 3.380 ;
        RECT 42.425 2.415 42.705 2.695 ;
        RECT 44.465 3.780 44.745 4.060 ;
        RECT 44.465 2.760 44.745 3.040 ;
        RECT 71.095 7.040 71.375 7.320 ;
        RECT 59.325 5.820 59.605 6.100 ;
        RECT 60.370 5.820 60.650 6.100 ;
        RECT 59.690 4.800 59.970 5.080 ;
        RECT 60.350 3.100 60.630 3.380 ;
        RECT 59.010 2.415 59.290 2.695 ;
        RECT 61.050 3.780 61.330 4.060 ;
        RECT 61.050 2.760 61.330 3.040 ;
        RECT 75.905 5.820 76.185 6.100 ;
        RECT 76.950 5.820 77.230 6.100 ;
        RECT 76.270 4.800 76.550 5.080 ;
        RECT 76.930 3.100 77.210 3.380 ;
        RECT 75.590 2.415 75.870 2.695 ;
        RECT 77.630 3.780 77.910 4.060 ;
        RECT 77.630 2.760 77.910 3.040 ;
      LAYER met3 ;
        RECT 5.590 7.970 9.870 8.270 ;
        RECT 22.175 7.970 26.455 8.270 ;
        RECT 38.760 7.970 43.040 8.270 ;
        RECT 55.345 7.970 59.625 8.270 ;
        RECT 71.925 7.970 76.205 8.270 ;
        RECT 4.715 7.330 5.085 7.365 ;
        RECT 5.590 7.330 5.890 7.970 ;
        RECT 4.715 7.030 5.890 7.330 ;
        RECT 4.715 6.995 5.085 7.030 ;
        RECT 9.565 6.125 9.865 7.970 ;
        RECT 21.300 7.330 21.670 7.365 ;
        RECT 22.175 7.330 22.475 7.970 ;
        RECT 21.300 7.030 22.475 7.330 ;
        RECT 21.300 6.995 21.670 7.030 ;
        RECT 26.150 6.125 26.450 7.970 ;
        RECT 37.885 7.330 38.255 7.365 ;
        RECT 38.760 7.330 39.060 7.970 ;
        RECT 37.885 7.030 39.060 7.330 ;
        RECT 37.885 6.995 38.255 7.030 ;
        RECT 42.735 6.125 43.035 7.970 ;
        RECT 54.470 7.330 54.840 7.365 ;
        RECT 55.345 7.330 55.645 7.970 ;
        RECT 54.470 7.030 55.645 7.330 ;
        RECT 54.470 6.995 54.840 7.030 ;
        RECT 59.320 6.125 59.620 7.970 ;
        RECT 71.050 7.330 71.420 7.365 ;
        RECT 71.925 7.330 72.225 7.970 ;
        RECT 71.050 7.030 72.225 7.330 ;
        RECT 71.050 6.995 71.420 7.030 ;
        RECT 75.900 6.125 76.200 7.970 ;
        RECT 8.940 6.110 9.875 6.125 ;
        RECT 10.590 6.110 10.920 6.125 ;
        RECT 25.525 6.110 26.460 6.125 ;
        RECT 27.175 6.110 27.505 6.125 ;
        RECT 42.110 6.110 43.045 6.125 ;
        RECT 43.760 6.110 44.090 6.125 ;
        RECT 58.695 6.110 59.630 6.125 ;
        RECT 60.345 6.110 60.675 6.125 ;
        RECT 75.275 6.110 76.210 6.125 ;
        RECT 76.925 6.110 77.255 6.125 ;
        RECT 8.940 5.810 11.390 6.110 ;
        RECT 25.525 5.810 27.975 6.110 ;
        RECT 42.110 5.810 44.560 6.110 ;
        RECT 58.695 5.810 61.145 6.110 ;
        RECT 75.275 5.810 77.725 6.110 ;
        RECT 8.940 5.795 10.920 5.810 ;
        RECT 25.525 5.795 27.505 5.810 ;
        RECT 42.110 5.795 44.090 5.810 ;
        RECT 58.695 5.795 60.675 5.810 ;
        RECT 75.275 5.795 77.255 5.810 ;
        RECT 8.940 4.095 9.270 5.795 ;
        RECT 10.595 5.790 10.895 5.795 ;
        RECT 9.910 5.090 10.240 5.105 ;
        RECT 9.910 4.790 10.710 5.090 ;
        RECT 9.910 4.775 10.240 4.790 ;
        RECT 25.525 4.095 25.855 5.795 ;
        RECT 27.180 5.790 27.480 5.795 ;
        RECT 26.495 5.090 26.825 5.105 ;
        RECT 26.495 4.790 27.295 5.090 ;
        RECT 26.495 4.775 26.825 4.790 ;
        RECT 42.110 4.095 42.440 5.795 ;
        RECT 43.765 5.790 44.065 5.795 ;
        RECT 43.080 5.090 43.410 5.105 ;
        RECT 43.080 4.790 43.880 5.090 ;
        RECT 43.080 4.775 43.410 4.790 ;
        RECT 58.695 4.095 59.025 5.795 ;
        RECT 60.350 5.790 60.650 5.795 ;
        RECT 59.665 5.090 59.995 5.105 ;
        RECT 59.665 4.790 60.465 5.090 ;
        RECT 59.665 4.775 59.995 4.790 ;
        RECT 75.275 4.095 75.605 5.795 ;
        RECT 76.930 5.790 77.230 5.795 ;
        RECT 76.245 5.090 76.575 5.105 ;
        RECT 76.245 4.790 77.045 5.090 ;
        RECT 76.245 4.775 76.575 4.790 ;
        RECT 8.940 4.085 11.235 4.095 ;
        RECT 25.525 4.085 27.820 4.095 ;
        RECT 42.110 4.085 44.405 4.095 ;
        RECT 58.695 4.085 60.990 4.095 ;
        RECT 75.275 4.085 77.570 4.095 ;
        RECT 8.940 4.070 11.600 4.085 ;
        RECT 25.525 4.070 28.185 4.085 ;
        RECT 42.110 4.070 44.770 4.085 ;
        RECT 58.695 4.070 61.355 4.085 ;
        RECT 75.275 4.070 77.935 4.085 ;
        RECT 8.940 3.770 12.070 4.070 ;
        RECT 25.525 3.770 28.655 4.070 ;
        RECT 42.110 3.770 45.240 4.070 ;
        RECT 58.695 3.770 61.825 4.070 ;
        RECT 75.275 3.770 78.405 4.070 ;
        RECT 8.940 3.765 11.600 3.770 ;
        RECT 25.525 3.765 28.185 3.770 ;
        RECT 42.110 3.765 44.770 3.770 ;
        RECT 58.695 3.765 61.355 3.770 ;
        RECT 75.275 3.765 77.935 3.770 ;
        RECT 11.270 3.755 11.600 3.765 ;
        RECT 27.855 3.755 28.185 3.765 ;
        RECT 44.440 3.755 44.770 3.765 ;
        RECT 61.025 3.755 61.355 3.765 ;
        RECT 77.605 3.755 77.935 3.765 ;
        RECT 11.275 3.705 11.575 3.755 ;
        RECT 27.860 3.705 28.160 3.755 ;
        RECT 44.445 3.705 44.745 3.755 ;
        RECT 61.030 3.705 61.330 3.755 ;
        RECT 77.610 3.705 77.910 3.755 ;
        RECT 10.570 3.390 10.900 3.405 ;
        RECT 27.155 3.390 27.485 3.405 ;
        RECT 43.740 3.390 44.070 3.405 ;
        RECT 60.325 3.390 60.655 3.405 ;
        RECT 76.905 3.390 77.235 3.405 ;
        RECT 10.100 3.090 10.900 3.390 ;
        RECT 26.685 3.090 27.485 3.390 ;
        RECT 43.270 3.090 44.070 3.390 ;
        RECT 59.855 3.090 60.655 3.390 ;
        RECT 76.435 3.090 77.235 3.390 ;
        RECT 10.570 3.075 10.900 3.090 ;
        RECT 27.155 3.075 27.485 3.090 ;
        RECT 43.740 3.075 44.070 3.090 ;
        RECT 60.325 3.075 60.655 3.090 ;
        RECT 76.905 3.075 77.235 3.090 ;
        RECT 10.595 3.060 10.895 3.075 ;
        RECT 11.270 3.050 11.600 3.065 ;
        RECT 27.180 3.060 27.480 3.075 ;
        RECT 27.855 3.050 28.185 3.065 ;
        RECT 43.765 3.060 44.065 3.075 ;
        RECT 44.440 3.050 44.770 3.065 ;
        RECT 60.350 3.060 60.650 3.075 ;
        RECT 61.025 3.050 61.355 3.065 ;
        RECT 76.930 3.060 77.230 3.075 ;
        RECT 77.605 3.050 77.935 3.065 ;
        RECT 11.270 2.750 12.070 3.050 ;
        RECT 27.855 2.750 28.655 3.050 ;
        RECT 44.440 2.750 45.240 3.050 ;
        RECT 61.025 2.750 61.825 3.050 ;
        RECT 77.605 2.750 78.405 3.050 ;
        RECT 11.270 2.735 11.600 2.750 ;
        RECT 27.855 2.735 28.185 2.750 ;
        RECT 44.440 2.735 44.770 2.750 ;
        RECT 61.025 2.735 61.355 2.750 ;
        RECT 77.605 2.735 77.935 2.750 ;
        RECT 11.270 2.730 11.590 2.735 ;
        RECT 27.855 2.730 28.175 2.735 ;
        RECT 44.440 2.730 44.760 2.735 ;
        RECT 61.025 2.730 61.345 2.735 ;
        RECT 77.605 2.730 77.925 2.735 ;
        RECT 8.760 2.705 9.120 2.710 ;
        RECT 9.230 2.705 9.560 2.720 ;
        RECT 8.760 2.410 9.560 2.705 ;
        RECT 25.345 2.705 25.705 2.710 ;
        RECT 25.815 2.705 26.145 2.720 ;
        RECT 25.345 2.410 26.145 2.705 ;
        RECT 41.930 2.705 42.290 2.710 ;
        RECT 42.400 2.705 42.730 2.720 ;
        RECT 41.930 2.410 42.730 2.705 ;
        RECT 58.515 2.705 58.875 2.710 ;
        RECT 58.985 2.705 59.315 2.720 ;
        RECT 58.515 2.410 59.315 2.705 ;
        RECT 75.095 2.705 75.455 2.710 ;
        RECT 75.565 2.705 75.895 2.720 ;
        RECT 75.095 2.410 75.895 2.705 ;
        RECT 9.120 2.405 9.560 2.410 ;
        RECT 25.705 2.405 26.145 2.410 ;
        RECT 42.290 2.405 42.730 2.410 ;
        RECT 58.875 2.405 59.315 2.410 ;
        RECT 75.455 2.405 75.895 2.410 ;
        RECT 9.230 2.390 9.560 2.405 ;
        RECT 25.815 2.390 26.145 2.405 ;
        RECT 42.400 2.390 42.730 2.405 ;
        RECT 58.985 2.390 59.315 2.405 ;
        RECT 75.565 2.390 75.895 2.405 ;
  END
END sky130_osu_ring_oscillator_mpr2ca_8_b0r1
END LIBRARY

