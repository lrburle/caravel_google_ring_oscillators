magic
tech sky130A
magscale 1 2
timestamp 1700015195
<< obsli1 >>
rect 292000 190000 528832 491776
<< obsm1 >>
rect 289722 187416 580230 491776
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
<< obsm2 >>
rect 289728 86119 580686 491776
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 292000 484836 583520 491776
rect 292000 484436 583440 484836
rect 292000 471644 583520 484436
rect 292000 471244 583440 471644
rect 292000 458316 583520 471244
rect 292000 457916 583440 458316
rect 292000 444988 583520 457916
rect 292000 444588 583440 444988
rect 292000 431796 583520 444588
rect 292000 431396 583440 431796
rect 292000 418468 583520 431396
rect 292000 418068 583440 418468
rect 292000 405140 583520 418068
rect 292000 404740 583440 405140
rect 292000 391948 583520 404740
rect 292000 391548 583440 391948
rect 292000 378620 583520 391548
rect 292000 378220 583440 378620
rect 292000 365292 583520 378220
rect 292000 364892 583440 365292
rect 292000 352100 583520 364892
rect 292000 351700 583440 352100
rect 292000 338772 583520 351700
rect 292000 338372 583440 338772
rect 292000 325444 583520 338372
rect 292000 325044 583440 325444
rect 292000 312252 583520 325044
rect 292000 311852 583440 312252
rect 292000 298924 583520 311852
rect 292000 298524 583440 298924
rect 292000 285596 583520 298524
rect 292000 285196 583440 285596
rect 292000 272404 583520 285196
rect 292000 272004 583440 272404
rect 292000 259076 583520 272004
rect 292000 258676 583440 259076
rect 292000 245748 583520 258676
rect 292000 245348 583440 245748
rect 292000 232556 583520 245348
rect 292000 232156 583440 232556
rect 292000 219228 583520 232156
rect 292000 218828 583440 219228
rect 292000 205900 583520 218828
rect 292000 205500 583440 205900
rect 292000 192708 583520 205500
rect 292000 192308 583440 192708
rect 292000 179380 583520 192308
rect 292000 178980 583440 179380
rect 292000 166052 583520 178980
rect 292000 165652 583440 166052
rect 292000 152860 583520 165652
rect 292000 152460 583440 152860
rect 292000 139532 583520 152460
rect 292000 139132 583440 139532
rect 292000 126204 583520 139132
rect 292000 125804 583440 126204
rect 292000 113012 583520 125804
rect 292000 112612 583440 113012
rect 292000 99684 583520 112612
rect 292000 99284 583440 99684
rect 292000 86356 583520 99284
rect 292000 85956 583440 86356
rect 292000 73164 583520 85956
rect 292000 72764 583440 73164
rect 292000 59836 583520 72764
rect 292000 59436 583440 59836
rect 292000 46508 583520 59436
rect 292000 46108 583440 46508
rect 292000 33316 583520 46108
rect 292000 32916 583440 33316
rect 292000 19988 583520 32916
rect 292000 19588 583440 19988
rect 292000 6796 583520 19588
rect 292000 6564 583440 6796
<< metal4 >>
rect -3236 -2164 -2636 706100
rect -2296 -1224 -1696 705160
rect 804 -2164 1404 706100
rect 4404 -2164 5004 706100
rect 38004 -2164 38604 706100
rect 41604 -2164 42204 706100
rect 75204 -2164 75804 706100
rect 78804 -2164 79404 706100
rect 112404 -2164 113004 706100
rect 116004 -2164 116604 706100
rect 149604 -2164 150204 706100
rect 153204 -2164 153804 706100
rect 186804 -2164 187404 706100
rect 190404 -2164 191004 706100
rect 224004 -2164 224604 706100
rect 227604 -2164 228204 706100
rect 261204 -2164 261804 706100
rect 264804 -2164 265404 706100
rect 298404 372781 299004 706100
rect 302004 372781 302604 706100
rect 298404 212781 299004 368377
rect 302004 212781 302604 368377
rect 298404 -2164 299004 208377
rect 302004 -2164 302604 208377
rect 335604 -2164 336204 706100
rect 339204 -2164 339804 706100
rect 372804 -2164 373404 706100
rect 376404 -2164 377004 706100
rect 410004 -2164 410604 706100
rect 413604 -2164 414204 706100
rect 447204 -2164 447804 706100
rect 450804 -2164 451404 706100
rect 484404 -2164 485004 706100
rect 488004 -2164 488604 706100
rect 521604 421752 522204 706100
rect 525204 421752 525804 706100
rect 521604 -2164 522204 240008
rect 525204 -2164 525804 240008
rect 558804 -2164 559404 706100
rect 562404 -2164 563004 706100
rect 585620 -1224 586220 705160
rect 586560 -2164 587160 706100
<< obsm4 >>
rect 293139 372701 298324 491469
rect 299084 372701 301924 491469
rect 302684 372701 335524 491469
rect 293139 368457 335524 372701
rect 293139 212701 298324 368457
rect 299084 212701 301924 368457
rect 302684 212701 335524 368457
rect 293139 208457 335524 212701
rect 293139 6563 298324 208457
rect 299084 6563 301924 208457
rect 302684 6563 335524 208457
rect 336284 6563 339124 491469
rect 339884 6563 372724 491469
rect 373484 6563 376324 491469
rect 377084 6563 409924 491469
rect 410684 6563 413524 491469
rect 414284 6563 447124 491469
rect 447884 6563 450724 491469
rect 451484 6563 484324 491469
rect 485084 6563 487924 491469
rect 488684 421672 521524 491469
rect 522284 421672 525124 491469
rect 525884 421672 531885 491469
rect 488684 240088 531885 421672
rect 488684 6563 521524 240088
rect 522284 6563 525124 240088
rect 525884 6563 531885 240088
<< metal5 >>
rect -3236 705500 587160 706100
rect -2296 704560 586220 705160
rect -3236 675076 587160 675676
rect -3236 671476 587160 672076
rect -3236 637876 587160 638476
rect -3236 634276 587160 634876
rect -3236 600676 587160 601276
rect -3236 597076 587160 597676
rect -3236 563476 587160 564076
rect -3236 559876 587160 560476
rect -3236 526276 587160 526876
rect -3236 522676 587160 523276
rect -3236 489076 587160 489676
rect -3236 485476 587160 486076
rect -3236 451876 587160 452476
rect -3236 448276 587160 448876
rect -3236 414676 587160 415276
rect -3236 411076 587160 411676
rect -3236 377476 587160 378076
rect -3236 373876 587160 374476
rect -3236 340276 587160 340876
rect -3236 336676 587160 337276
rect -3236 303076 587160 303676
rect -3236 299476 587160 300076
rect -3236 265876 587160 266476
rect -3236 262276 587160 262876
rect -3236 228676 587160 229276
rect -3236 225076 587160 225676
rect -3236 191476 587160 192076
rect -3236 187876 587160 188476
rect -3236 154276 587160 154876
rect -3236 150676 587160 151276
rect -3236 117076 587160 117676
rect -3236 113476 587160 114076
rect -3236 79876 587160 80476
rect -3236 76276 587160 76876
rect -3236 42676 587160 43276
rect -3236 39076 587160 39676
rect -3236 5476 587160 6076
rect -3236 1876 587160 2476
rect -2296 -1224 586220 -624
rect -3236 -2164 587160 -1564
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal4 s -2296 -1224 -1696 705160 4 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -2296 -1224 586220 -624 8 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -2296 704560 586220 705160 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 585620 -1224 586220 705160 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 804 -2164 1404 706100 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 38004 -2164 38604 706100 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 75204 -2164 75804 706100 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 112404 -2164 113004 706100 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 149604 -2164 150204 706100 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 186804 -2164 187404 706100 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 224004 -2164 224604 706100 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 261204 -2164 261804 706100 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 298404 -2164 299004 208377 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 298404 212781 299004 368377 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 298404 372781 299004 706100 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 335604 -2164 336204 706100 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 372804 -2164 373404 706100 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 410004 -2164 410604 706100 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 447204 -2164 447804 706100 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 484404 -2164 485004 706100 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 521604 -2164 522204 240008 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 521604 421752 522204 706100 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s 558804 -2164 559404 706100 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 1876 587160 2476 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 39076 587160 39676 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 76276 587160 76876 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 113476 587160 114076 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 150676 587160 151276 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 187876 587160 188476 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 225076 587160 225676 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 262276 587160 262876 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 299476 587160 300076 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 336676 587160 337276 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 373876 587160 374476 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 411076 587160 411676 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 448276 587160 448876 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 485476 587160 486076 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 522676 587160 523276 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 559876 587160 560476 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 597076 587160 597676 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 634276 587160 634876 6 vccd1
port 144 nsew power bidirectional
rlabel metal5 s -3236 671476 587160 672076 6 vccd1
port 144 nsew power bidirectional
rlabel metal4 s -3236 -2164 -2636 706100 4 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 -2164 587160 -1564 8 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 705500 587160 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 586560 -2164 587160 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 4404 -2164 5004 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 41604 -2164 42204 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 78804 -2164 79404 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 116004 -2164 116604 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 153204 -2164 153804 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 190404 -2164 191004 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 227604 -2164 228204 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 264804 -2164 265404 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 302004 -2164 302604 208377 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 302004 212781 302604 368377 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 302004 372781 302604 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 339204 -2164 339804 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 376404 -2164 377004 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 413604 -2164 414204 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 450804 -2164 451404 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 488004 -2164 488604 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 525204 -2164 525804 240008 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 525204 421752 525804 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal4 s 562404 -2164 563004 706100 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 5476 587160 6076 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 42676 587160 43276 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 79876 587160 80476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 117076 587160 117676 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 154276 587160 154876 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 191476 587160 192076 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 228676 587160 229276 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 265876 587160 266476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 303076 587160 303676 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 340276 587160 340876 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 377476 587160 378076 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 414676 587160 415276 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 451876 587160 452476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 489076 587160 489676 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 526276 587160 526876 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 563476 587160 564076 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 600676 587160 601276 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 637876 587160 638476 6 vssd1
port 145 nsew ground bidirectional
rlabel metal5 s -3236 675076 587160 675676 6 vssd1
port 145 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 146 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 147 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 148 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 149 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 150 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 151 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 152 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 153 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 154 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 155 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 156 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 157 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 158 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 159 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 160 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 161 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 162 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 163 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 164 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 165 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 166 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 167 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 168 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 169 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 170 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 171 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 172 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 173 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 174 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 175 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 176 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 177 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 178 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 179 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 180 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 181 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 182 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 183 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 184 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 185 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 186 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 187 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 188 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 189 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 190 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 191 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 192 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 193 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 194 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 195 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 196 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 197 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 198 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 199 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 200 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 201 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 202 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 203 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 204 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 205 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 206 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 207 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 208 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 209 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 210 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 211 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 212 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 213 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 214 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 215 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 216 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 217 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 218 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 219 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 220 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 221 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 222 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 223 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 224 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 225 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 226 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 227 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 228 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 229 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 230 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 231 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 232 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 233 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 234 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 235 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 236 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 237 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 238 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 239 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 240 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 241 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 242 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 243 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 244 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 245 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 246 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 247 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 248 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 249 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 250 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 251 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2724116
string GDS_FILE /import/yukari1/lrburle/google_ring_oscillator/caravel/openlane/user_project_wrapper/runs/23_11_14_20_24/results/signoff/user_project_wrapper.magic.gds
string GDS_START 2371178
<< end >>

