magic
tech sky130A
magscale 1 2
timestamp 1703008989
<< obsli1 >>
rect 1104 2159 28888 7633
<< obsm1 >>
rect 934 2128 29048 7664
<< metal2 >>
rect 2962 9200 3018 10000
rect 8942 9200 8998 10000
rect 14922 9200 14978 10000
rect 20902 9200 20958 10000
rect 26882 9200 26938 10000
<< obsm2 >>
rect 938 9144 2906 9330
rect 3074 9144 8886 9330
rect 9054 9144 14866 9330
rect 15034 9144 20846 9330
rect 21014 9144 26826 9330
rect 26994 9144 29042 9330
rect 938 1119 29042 9144
<< metal3 >>
rect 29200 8712 30000 8832
rect 29200 6808 30000 6928
rect 0 4904 800 5024
rect 29200 4904 30000 5024
rect 29200 3000 30000 3120
rect 29200 1096 30000 1216
<< obsm3 >>
rect 800 8632 29120 8805
rect 800 7008 29200 8632
rect 800 6728 29120 7008
rect 800 5104 29200 6728
rect 880 4824 29120 5104
rect 800 3200 29200 4824
rect 800 2920 29120 3200
rect 800 1296 29200 2920
rect 800 1123 29120 1296
<< metal4 >>
rect 4417 2128 4737 7664
rect 7890 2128 8210 7664
rect 11363 2128 11683 7664
rect 14836 2128 15156 7664
rect 18309 2128 18629 7664
rect 21782 2128 22102 7664
rect 25255 2128 25575 7664
rect 28728 2128 29048 7664
<< labels >>
rlabel metal3 s 29200 1096 30000 1216 6 X1_Y1
port 1 nsew signal output
rlabel metal3 s 29200 3000 30000 3120 6 X2_Y1
port 2 nsew signal output
rlabel metal3 s 29200 4904 30000 5024 6 X3_Y1
port 3 nsew signal output
rlabel metal3 s 29200 6808 30000 6928 6 X4_Y1
port 4 nsew signal output
rlabel metal3 s 29200 8712 30000 8832 6 X5_Y1
port 5 nsew signal output
rlabel metal2 s 2962 9200 3018 10000 6 s1
port 6 nsew signal input
rlabel metal2 s 8942 9200 8998 10000 6 s2
port 7 nsew signal input
rlabel metal2 s 14922 9200 14978 10000 6 s3
port 8 nsew signal input
rlabel metal2 s 20902 9200 20958 10000 6 s4
port 9 nsew signal input
rlabel metal2 s 26882 9200 26938 10000 6 s5
port 10 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 start
port 11 nsew signal input
rlabel metal4 s 4417 2128 4737 7664 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 11363 2128 11683 7664 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 18309 2128 18629 7664 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 25255 2128 25575 7664 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 7890 2128 8210 7664 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 14836 2128 15156 7664 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 21782 2128 22102 7664 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 28728 2128 29048 7664 6 vssd1
port 13 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 359438
string GDS_FILE /import/yukari1/lrburle/google_ring_oscillator/caravel/openlane/b0r1_aa/runs/23_12_19_12_02/results/signoff/b0r1_aa.magic.gds
string GDS_START 293088
<< end >>

